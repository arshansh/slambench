// (C) 1992-2015 Altera Corporation. All rights reserved.                         
// Your use of Altera Corporation's design tools, logic functions and other       
// software and tools, and its AMPP partner logic functions, and any output       
// files any of the foregoing (including device programming or simulation         
// files), and any associated documentation or information are expressly subject  
// to the terms and conditions of the Altera Program License Subscription         
// Agreement, Altera MegaCore Function License Agreement, or other applicable     
// license agreement, including, without limitation, that your use is for the     
// sole purpose of programming logic devices manufactured by Altera and sold by   
// Altera or its authorized distributors.  Please refer to the applicable         
// agreement for further details.                                                 
    

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_0
	(
		input 		clock,
		input 		resetn,
		input 		start,
		input [31:0] 		input_r,
		input [31:0] 		input_global_size_0,
		input [31:0] 		input_global_size_1,
		input [31:0] 		input_e_d,
		input 		valid_in,
		output 		stall_out,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		input [31:0] 		input_acl_hw_wg_id,
		output 		valid_out,
		input 		stall_in,
		output 		lvb_bb0_cmp1622,
		output [31:0] 		lvb_bb0_sub25,
		output [31:0] 		lvb_bb0_sub29,
		output [31:0] 		lvb_bb0_mul50,
		output [63:0] 		lvb_bb0_var_,
		output [63:0] 		lvb_bb0_var__u0,
		output [31:0] 		lvb_input_global_id_0,
		output [31:0] 		lvb_input_global_id_1,
		output [31:0] 		lvb_input_acl_hw_wg_id,
		input [31:0] 		workgroup_size
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_global_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_global_id_0_staging_reg_NO_SHIFT_REG <= input_global_id_0;
				input_global_id_1_staging_reg_NO_SHIFT_REG <= input_global_id_1;
				input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub_inputs_ready;
 reg local_bb0_sub_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub_valid_out_0_NO_SHIFT_REG;
wire local_bb0_sub_stall_in_0;
 reg local_bb0_sub_valid_out_1_NO_SHIFT_REG;
wire local_bb0_sub_stall_in_1;
wire local_bb0_sub_output_regs_ready;
 reg [31:0] local_bb0_sub_NO_SHIFT_REG;
wire local_bb0_sub_causedstall;

assign local_bb0_sub_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb0_sub_output_regs_ready = (~(local_bb0_sub_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_sub_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_sub_stall_in_0)) & (~(local_bb0_sub_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_sub_stall_in_1))));
assign merge_node_stall_in_0 = (~(local_bb0_sub_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub_output_regs_ready) | ~(local_bb0_sub_inputs_ready)));
assign local_bb0_sub_causedstall = (local_bb0_sub_inputs_ready && (~(local_bb0_sub_output_regs_ready) && !(~(local_bb0_sub_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub_NO_SHIFT_REG <= 'x;
		local_bb0_sub_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_sub_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub_NO_SHIFT_REG <= 'x;
			local_bb0_sub_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_sub_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub_output_regs_ready)
			begin
				local_bb0_sub_NO_SHIFT_REG <= (32'h0 - input_r);
				local_bb0_sub_valid_out_0_NO_SHIFT_REG <= local_bb0_sub_inputs_ready;
				local_bb0_sub_valid_out_1_NO_SHIFT_REG <= local_bb0_sub_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub_stall_in_0))
				begin
					local_bb0_sub_valid_out_0_NO_SHIFT_REG <= local_bb0_sub_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_sub_stall_in_1))
				begin
					local_bb0_sub_valid_out_1_NO_SHIFT_REG <= local_bb0_sub_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub_inputs_ready)
			begin
				local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub25_inputs_ready;
 reg local_bb0_sub25_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub25_valid_out_NO_SHIFT_REG;
wire local_bb0_sub25_stall_in;
wire local_bb0_sub25_output_regs_ready;
 reg [31:0] local_bb0_sub25_NO_SHIFT_REG;
wire local_bb0_sub25_causedstall;

assign local_bb0_sub25_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign local_bb0_sub25_output_regs_ready = (~(local_bb0_sub25_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_sub25_valid_out_NO_SHIFT_REG) | ~(local_bb0_sub25_stall_in))));
assign merge_node_stall_in_2 = (~(local_bb0_sub25_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub25_output_regs_ready) | ~(local_bb0_sub25_inputs_ready)));
assign local_bb0_sub25_causedstall = (local_bb0_sub25_inputs_ready && (~(local_bb0_sub25_output_regs_ready) && !(~(local_bb0_sub25_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub25_NO_SHIFT_REG <= 'x;
		local_bb0_sub25_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub25_NO_SHIFT_REG <= 'x;
			local_bb0_sub25_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub25_output_regs_ready)
			begin
				local_bb0_sub25_NO_SHIFT_REG <= (input_global_size_0 + 32'hFFFFFFFF);
				local_bb0_sub25_valid_out_NO_SHIFT_REG <= local_bb0_sub25_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub25_stall_in))
				begin
					local_bb0_sub25_valid_out_NO_SHIFT_REG <= local_bb0_sub25_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub25_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub25_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub25_inputs_ready)
			begin
				local_bb0_sub25_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub29_inputs_ready;
 reg local_bb0_sub29_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub29_valid_out_NO_SHIFT_REG;
wire local_bb0_sub29_stall_in;
wire local_bb0_sub29_output_regs_ready;
 reg [31:0] local_bb0_sub29_NO_SHIFT_REG;
wire local_bb0_sub29_causedstall;

assign local_bb0_sub29_inputs_ready = merge_node_valid_out_3_NO_SHIFT_REG;
assign local_bb0_sub29_output_regs_ready = (~(local_bb0_sub29_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_sub29_valid_out_NO_SHIFT_REG) | ~(local_bb0_sub29_stall_in))));
assign merge_node_stall_in_3 = (~(local_bb0_sub29_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub29_output_regs_ready) | ~(local_bb0_sub29_inputs_ready)));
assign local_bb0_sub29_causedstall = (local_bb0_sub29_inputs_ready && (~(local_bb0_sub29_output_regs_ready) && !(~(local_bb0_sub29_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub29_NO_SHIFT_REG <= 'x;
		local_bb0_sub29_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub29_NO_SHIFT_REG <= 'x;
			local_bb0_sub29_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub29_output_regs_ready)
			begin
				local_bb0_sub29_NO_SHIFT_REG <= (input_global_size_1 + 32'hFFFFFFFF);
				local_bb0_sub29_valid_out_NO_SHIFT_REG <= local_bb0_sub29_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub29_stall_in))
				begin
					local_bb0_sub29_valid_out_NO_SHIFT_REG <= local_bb0_sub29_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub29_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub29_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub29_inputs_ready)
			begin
				local_bb0_sub29_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u1_inputs_ready;
 reg local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u1_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u1_stall_in;
wire local_bb0_var__u1_output_regs_ready;
 reg [31:0] local_bb0_var__u1_NO_SHIFT_REG;
wire local_bb0_var__u1_causedstall;

assign local_bb0_var__u1_inputs_ready = merge_node_valid_out_4_NO_SHIFT_REG;
assign local_bb0_var__u1_output_regs_ready = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u1_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u1_stall_in))));
assign merge_node_stall_in_4 = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u1_output_regs_ready) | ~(local_bb0_var__u1_inputs_ready)));
assign local_bb0_var__u1_causedstall = (local_bb0_var__u1_inputs_ready && (~(local_bb0_var__u1_output_regs_ready) && !(~(local_bb0_var__u1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_NO_SHIFT_REG <= 'x;
		local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_NO_SHIFT_REG <= 'x;
			local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_output_regs_ready)
			begin
				local_bb0_var__u1_NO_SHIFT_REG <= input_e_d;
				local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u1_stall_in))
				begin
					local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_inputs_ready)
			begin
				local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u0_inputs_ready;
 reg local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u0_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u0_stall_in;
wire local_bb0_var__u0_output_regs_ready;
 reg [63:0] local_bb0_var__u0_NO_SHIFT_REG;
wire local_bb0_var__u0_causedstall;

assign local_bb0_var__u0_inputs_ready = merge_node_valid_out_6_NO_SHIFT_REG;
assign local_bb0_var__u0_output_regs_ready = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u0_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u0_stall_in))));
assign merge_node_stall_in_6 = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u0_output_regs_ready) | ~(local_bb0_var__u0_inputs_ready)));
assign local_bb0_var__u0_causedstall = (local_bb0_var__u0_inputs_ready && (~(local_bb0_var__u0_output_regs_ready) && !(~(local_bb0_var__u0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_NO_SHIFT_REG <= 'x;
		local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_NO_SHIFT_REG <= 'x;
			local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_output_regs_ready)
			begin
				local_bb0_var__u0_NO_SHIFT_REG <= $signed(input_r);
				local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u0_stall_in))
				begin
					local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_inputs_ready)
			begin
				local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp1622_inputs_ready;
 reg local_bb0_cmp1622_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp1622_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp1622_stall_in;
wire local_bb0_cmp1622_output_regs_ready;
 reg local_bb0_cmp1622_NO_SHIFT_REG;
wire local_bb0_cmp1622_causedstall;

assign local_bb0_cmp1622_inputs_ready = (local_bb0_sub_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign local_bb0_cmp1622_output_regs_ready = (~(local_bb0_cmp1622_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp1622_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp1622_stall_in))));
assign local_bb0_sub_stall_in_0 = (~(local_bb0_cmp1622_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp1622_output_regs_ready) | ~(local_bb0_cmp1622_inputs_ready)));
assign merge_node_stall_in_1 = (~(local_bb0_cmp1622_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp1622_output_regs_ready) | ~(local_bb0_cmp1622_inputs_ready)));
assign local_bb0_cmp1622_causedstall = (local_bb0_cmp1622_inputs_ready && (~(local_bb0_cmp1622_output_regs_ready) && !(~(local_bb0_cmp1622_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp1622_NO_SHIFT_REG <= 'x;
		local_bb0_cmp1622_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp1622_NO_SHIFT_REG <= 'x;
			local_bb0_cmp1622_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp1622_output_regs_ready)
			begin
				local_bb0_cmp1622_NO_SHIFT_REG <= ($signed(local_bb0_sub_NO_SHIFT_REG) > $signed(input_r));
				local_bb0_cmp1622_valid_out_NO_SHIFT_REG <= local_bb0_cmp1622_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp1622_stall_in))
				begin
					local_bb0_cmp1622_valid_out_NO_SHIFT_REG <= local_bb0_cmp1622_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp1622_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp1622_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp1622_inputs_ready)
			begin
				local_bb0_cmp1622_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__inputs_ready;
 reg local_bb0_var__wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__valid_out_NO_SHIFT_REG;
wire local_bb0_var__stall_in;
wire local_bb0_var__output_regs_ready;
 reg [63:0] local_bb0_var__NO_SHIFT_REG;
wire local_bb0_var__causedstall;

assign local_bb0_var__inputs_ready = local_bb0_sub_valid_out_1_NO_SHIFT_REG;
assign local_bb0_var__output_regs_ready = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__valid_out_NO_SHIFT_REG) | ~(local_bb0_var__stall_in))));
assign local_bb0_sub_stall_in_1 = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__output_regs_ready) | ~(local_bb0_var__inputs_ready)));
assign local_bb0_var__causedstall = (local_bb0_var__inputs_ready && (~(local_bb0_var__output_regs_ready) && !(~(local_bb0_var__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__NO_SHIFT_REG <= 'x;
		local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__NO_SHIFT_REG <= 'x;
			local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__output_regs_ready)
			begin
				local_bb0_var__NO_SHIFT_REG <= $signed(local_bb0_sub_NO_SHIFT_REG);
				local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__stall_in))
				begin
					local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__inputs_ready)
			begin
				local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_2to2_bb0_var__u1_valid_out_0;
wire rstag_2to2_bb0_var__u1_stall_in_0;
wire rstag_2to2_bb0_var__u1_valid_out_1;
wire rstag_2to2_bb0_var__u1_stall_in_1;
wire rstag_2to2_bb0_var__u1_valid_out_2;
wire rstag_2to2_bb0_var__u1_stall_in_2;
wire rstag_2to2_bb0_var__u1_inputs_ready;
wire rstag_2to2_bb0_var__u1_stall_local;
 reg rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG;
wire rstag_2to2_bb0_var__u1_combined_valid;
 reg [31:0] rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_2to2_bb0_var__u1;
 reg rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG;
 reg rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG;
 reg rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG;

assign rstag_2to2_bb0_var__u1_inputs_ready = local_bb0_var__u1_valid_out_NO_SHIFT_REG;
assign rstag_2to2_bb0_var__u1 = (rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG ? rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG : local_bb0_var__u1_NO_SHIFT_REG);
assign rstag_2to2_bb0_var__u1_combined_valid = (rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG | rstag_2to2_bb0_var__u1_inputs_ready);
assign rstag_2to2_bb0_var__u1_stall_local = ((rstag_2to2_bb0_var__u1_stall_in_0 & ~(rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG)) | (rstag_2to2_bb0_var__u1_stall_in_1 & ~(rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG)) | (rstag_2to2_bb0_var__u1_stall_in_2 & ~(rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG)));
assign rstag_2to2_bb0_var__u1_valid_out_0 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG));
assign rstag_2to2_bb0_var__u1_valid_out_1 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG));
assign rstag_2to2_bb0_var__u1_valid_out_2 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG));
assign local_bb0_var__u1_stall_in = (|rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_2to2_bb0_var__u1_stall_local)
			begin
				if (~(rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG))
				begin
					rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= rstag_2to2_bb0_var__u1_inputs_ready;
				end
			end
			else
			begin
				rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG))
		begin
			rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG <= local_bb0_var__u1_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_0)) & rstag_2to2_bb0_var__u1_stall_local);
			rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_1)) & rstag_2to2_bb0_var__u1_stall_local);
			rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_2)) & rstag_2to2_bb0_var__u1_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and33_i_inputs_ready;
 reg local_bb0_and33_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and33_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and33_i_stall_in;
wire local_bb0_and33_i_output_regs_ready;
 reg [31:0] local_bb0_and33_i_NO_SHIFT_REG;
wire local_bb0_and33_i_causedstall;

assign local_bb0_and33_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_0;
assign local_bb0_and33_i_output_regs_ready = (~(local_bb0_and33_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and33_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and33_i_stall_in))));
assign rstag_2to2_bb0_var__u1_stall_in_0 = (~(local_bb0_and33_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and33_i_output_regs_ready) | ~(local_bb0_and33_i_inputs_ready)));
assign local_bb0_and33_i_causedstall = (local_bb0_and33_i_inputs_ready && (~(local_bb0_and33_i_output_regs_ready) && !(~(local_bb0_and33_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and33_i_NO_SHIFT_REG <= 'x;
		local_bb0_and33_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and33_i_NO_SHIFT_REG <= 'x;
			local_bb0_and33_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and33_i_output_regs_ready)
			begin
				local_bb0_and33_i_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1 & 32'h807FFFFF);
				local_bb0_and33_i_valid_out_NO_SHIFT_REG <= local_bb0_and33_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and33_i_stall_in))
				begin
					local_bb0_and33_i_valid_out_NO_SHIFT_REG <= local_bb0_and33_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and33_i_inputs_ready)
			begin
				local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_and2_i_valid_out;
wire local_bb0_and2_i_stall_in;
wire local_bb0_and2_i_inputs_ready;
wire local_bb0_and2_i_stall_local;
wire [31:0] local_bb0_and2_i;

assign local_bb0_and2_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_1;
assign local_bb0_and2_i = (rstag_2to2_bb0_var__u1 & 32'h7FFFFF);
assign local_bb0_and2_i_valid_out = local_bb0_and2_i_inputs_ready;
assign local_bb0_and2_i_stall_local = local_bb0_and2_i_stall_in;
assign rstag_2to2_bb0_var__u1_stall_in_1 = (|local_bb0_and2_i_stall_local);

// This section implements a registered operation.
// 
wire local_bb0_shr_i_inputs_ready;
 reg local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_shr_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_shr_i_stall_in_0;
 reg local_bb0_shr_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_shr_i_stall_in_1;
wire local_bb0_shr_i_output_regs_ready;
 reg [31:0] local_bb0_shr_i_NO_SHIFT_REG;
wire local_bb0_shr_i_causedstall;

assign local_bb0_shr_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_2;
assign local_bb0_shr_i_output_regs_ready = (~(local_bb0_shr_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_shr_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_shr_i_stall_in_0)) & (~(local_bb0_shr_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_shr_i_stall_in_1))));
assign rstag_2to2_bb0_var__u1_stall_in_2 = (~(local_bb0_shr_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_shr_i_output_regs_ready) | ~(local_bb0_shr_i_inputs_ready)));
assign local_bb0_shr_i_causedstall = (local_bb0_shr_i_inputs_ready && (~(local_bb0_shr_i_output_regs_ready) && !(~(local_bb0_shr_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_shr_i_NO_SHIFT_REG <= 'x;
		local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_shr_i_NO_SHIFT_REG <= 'x;
			local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_shr_i_output_regs_ready)
			begin
				local_bb0_shr_i_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1 >> 32'h17);
				local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= local_bb0_shr_i_inputs_ready;
				local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= local_bb0_shr_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_shr_i_stall_in_0))
				begin
					local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_shr_i_stall_in_1))
				begin
					local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_shr_i_inputs_ready)
			begin
				local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_lnot6_i_inputs_ready;
 reg local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_lnot6_i_valid_out_NO_SHIFT_REG;
wire local_bb0_lnot6_i_stall_in;
wire local_bb0_lnot6_i_output_regs_ready;
 reg local_bb0_lnot6_i_NO_SHIFT_REG;
wire local_bb0_lnot6_i_causedstall;

assign local_bb0_lnot6_i_inputs_ready = local_bb0_and2_i_valid_out;
assign local_bb0_lnot6_i_output_regs_ready = (~(local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_lnot6_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_lnot6_i_stall_in))));
assign local_bb0_and2_i_stall_in = (~(local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_lnot6_i_output_regs_ready) | ~(local_bb0_lnot6_i_inputs_ready)));
assign local_bb0_lnot6_i_causedstall = (local_bb0_lnot6_i_inputs_ready && (~(local_bb0_lnot6_i_output_regs_ready) && !(~(local_bb0_lnot6_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_lnot6_i_NO_SHIFT_REG <= 'x;
		local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_lnot6_i_NO_SHIFT_REG <= 'x;
			local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_lnot6_i_output_regs_ready)
			begin
				local_bb0_lnot6_i_NO_SHIFT_REG <= ((local_bb0_and2_i & 32'h7FFFFF) != 32'h0);
				local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= local_bb0_lnot6_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_lnot6_i_stall_in))
				begin
					local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_lnot6_i_inputs_ready)
			begin
				local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and1_i_inputs_ready;
 reg local_bb0_and1_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and1_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and1_i_stall_in;
wire local_bb0_and1_i_output_regs_ready;
 reg [31:0] local_bb0_and1_i_NO_SHIFT_REG;
wire local_bb0_and1_i_causedstall;

assign local_bb0_and1_i_inputs_ready = local_bb0_shr_i_valid_out_0_NO_SHIFT_REG;
assign local_bb0_and1_i_output_regs_ready = (~(local_bb0_and1_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and1_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and1_i_stall_in))));
assign local_bb0_shr_i_stall_in_0 = (~(local_bb0_and1_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and1_i_output_regs_ready) | ~(local_bb0_and1_i_inputs_ready)));
assign local_bb0_and1_i_causedstall = (local_bb0_and1_i_inputs_ready && (~(local_bb0_and1_i_output_regs_ready) && !(~(local_bb0_and1_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and1_i_NO_SHIFT_REG <= 'x;
		local_bb0_and1_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and1_i_NO_SHIFT_REG <= 'x;
			local_bb0_and1_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and1_i_output_regs_ready)
			begin
				local_bb0_and1_i_NO_SHIFT_REG <= ((local_bb0_shr_i_NO_SHIFT_REG & 32'h1FF) & 32'hFF);
				local_bb0_and1_i_valid_out_NO_SHIFT_REG <= local_bb0_and1_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and1_i_stall_in))
				begin
					local_bb0_and1_i_valid_out_NO_SHIFT_REG <= local_bb0_and1_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and1_i_inputs_ready)
			begin
				local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_4to4_bb0_and1_i_valid_out_0;
wire rstag_4to4_bb0_and1_i_stall_in_0;
wire rstag_4to4_bb0_and1_i_valid_out_1;
wire rstag_4to4_bb0_and1_i_stall_in_1;
wire rstag_4to4_bb0_and1_i_valid_out_2;
wire rstag_4to4_bb0_and1_i_stall_in_2;
wire rstag_4to4_bb0_and1_i_inputs_ready;
wire rstag_4to4_bb0_and1_i_stall_local;
 reg rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG;
wire rstag_4to4_bb0_and1_i_combined_valid;
 reg [31:0] rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_4to4_bb0_and1_i;
 reg rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG;
 reg rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG;
 reg rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG;

assign rstag_4to4_bb0_and1_i_inputs_ready = local_bb0_and1_i_valid_out_NO_SHIFT_REG;
assign rstag_4to4_bb0_and1_i = (rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG ? rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG : (local_bb0_and1_i_NO_SHIFT_REG & 32'hFF));
assign rstag_4to4_bb0_and1_i_combined_valid = (rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG | rstag_4to4_bb0_and1_i_inputs_ready);
assign rstag_4to4_bb0_and1_i_stall_local = ((rstag_4to4_bb0_and1_i_stall_in_0 & ~(rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG)) | (rstag_4to4_bb0_and1_i_stall_in_1 & ~(rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG)) | (rstag_4to4_bb0_and1_i_stall_in_2 & ~(rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG)));
assign rstag_4to4_bb0_and1_i_valid_out_0 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG));
assign rstag_4to4_bb0_and1_i_valid_out_1 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG));
assign rstag_4to4_bb0_and1_i_valid_out_2 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG));
assign local_bb0_and1_i_stall_in = (|rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_4to4_bb0_and1_i_stall_local)
			begin
				if (~(rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= rstag_4to4_bb0_and1_i_inputs_ready;
				end
			end
			else
			begin
				rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG <= (local_bb0_and1_i_NO_SHIFT_REG & 32'hFF);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_0)) & rstag_4to4_bb0_and1_i_stall_local);
			rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_1)) & rstag_4to4_bb0_and1_i_stall_local);
			rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_2)) & rstag_4to4_bb0_and1_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp10_i_inputs_ready;
 reg local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_cmp10_i_stall_in_0;
 reg local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_cmp10_i_stall_in_1;
wire local_bb0_cmp10_i_output_regs_ready;
 reg local_bb0_cmp10_i_NO_SHIFT_REG;
wire local_bb0_cmp10_i_causedstall;

assign local_bb0_cmp10_i_inputs_ready = rstag_4to4_bb0_and1_i_valid_out_1;
assign local_bb0_cmp10_i_output_regs_ready = (~(local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_cmp10_i_stall_in_0)) & (~(local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_cmp10_i_stall_in_1))));
assign rstag_4to4_bb0_and1_i_stall_in_1 = (~(local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp10_i_output_regs_ready) | ~(local_bb0_cmp10_i_inputs_ready)));
assign local_bb0_cmp10_i_causedstall = (local_bb0_cmp10_i_inputs_ready && (~(local_bb0_cmp10_i_output_regs_ready) && !(~(local_bb0_cmp10_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp10_i_NO_SHIFT_REG <= 'x;
		local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp10_i_NO_SHIFT_REG <= 'x;
			local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp10_i_output_regs_ready)
			begin
				local_bb0_cmp10_i_NO_SHIFT_REG <= ((rstag_4to4_bb0_and1_i & 32'hFF) == 32'h0);
				local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp10_i_inputs_ready;
				local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp10_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp10_i_stall_in_0))
				begin
					local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_cmp10_i_stall_in_1))
				begin
					local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp10_i_inputs_ready)
			begin
				local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp_i_inputs_ready;
 reg local_bb0_cmp_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp_i_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp_i_stall_in;
wire local_bb0_cmp_i_output_regs_ready;
 reg local_bb0_cmp_i_NO_SHIFT_REG;
wire local_bb0_cmp_i_causedstall;

assign local_bb0_cmp_i_inputs_ready = rstag_4to4_bb0_and1_i_valid_out_2;
assign local_bb0_cmp_i_output_regs_ready = (~(local_bb0_cmp_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp_i_stall_in))));
assign rstag_4to4_bb0_and1_i_stall_in_2 = (~(local_bb0_cmp_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp_i_output_regs_ready) | ~(local_bb0_cmp_i_inputs_ready)));
assign local_bb0_cmp_i_causedstall = (local_bb0_cmp_i_inputs_ready && (~(local_bb0_cmp_i_output_regs_ready) && !(~(local_bb0_cmp_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp_i_NO_SHIFT_REG <= 'x;
		local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp_i_NO_SHIFT_REG <= 'x;
			local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp_i_output_regs_ready)
			begin
				local_bb0_cmp_i_NO_SHIFT_REG <= ((rstag_4to4_bb0_and1_i & 32'hFF) == 32'hFF);
				local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= local_bb0_cmp_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp_i_stall_in))
				begin
					local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= local_bb0_cmp_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp_i_inputs_ready)
			begin
				local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_not_cmp10_i_valid_out;
wire local_bb0_not_cmp10_i_stall_in;
wire local_bb0_not_cmp10_i_inputs_ready;
wire local_bb0_not_cmp10_i_stall_local;
wire local_bb0_not_cmp10_i;

assign local_bb0_not_cmp10_i_inputs_ready = local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG;
assign local_bb0_not_cmp10_i = (local_bb0_cmp10_i_NO_SHIFT_REG ^ 1'b1);
assign local_bb0_not_cmp10_i_valid_out = local_bb0_not_cmp10_i_inputs_ready;
assign local_bb0_not_cmp10_i_stall_local = local_bb0_not_cmp10_i_stall_in;
assign local_bb0_cmp10_i_stall_in_1 = (|local_bb0_not_cmp10_i_stall_local);

// This section implements a staging register.
// 
wire rstag_5to5_bb0_cmp_i_valid_out_0;
wire rstag_5to5_bb0_cmp_i_stall_in_0;
wire rstag_5to5_bb0_cmp_i_valid_out_1;
wire rstag_5to5_bb0_cmp_i_stall_in_1;
wire rstag_5to5_bb0_cmp_i_valid_out_2;
wire rstag_5to5_bb0_cmp_i_stall_in_2;
wire rstag_5to5_bb0_cmp_i_valid_out_3;
wire rstag_5to5_bb0_cmp_i_stall_in_3;
wire rstag_5to5_bb0_cmp_i_inputs_ready;
wire rstag_5to5_bb0_cmp_i_stall_local;
 reg rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb0_cmp_i_combined_valid;
 reg rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG;
wire rstag_5to5_bb0_cmp_i;
 reg rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG;

assign rstag_5to5_bb0_cmp_i_inputs_ready = local_bb0_cmp_i_valid_out_NO_SHIFT_REG;
assign rstag_5to5_bb0_cmp_i = (rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG : local_bb0_cmp_i_NO_SHIFT_REG);
assign rstag_5to5_bb0_cmp_i_combined_valid = (rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG | rstag_5to5_bb0_cmp_i_inputs_ready);
assign rstag_5to5_bb0_cmp_i_stall_local = ((rstag_5to5_bb0_cmp_i_stall_in_0 & ~(rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_1 & ~(rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_2 & ~(rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_3 & ~(rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG)));
assign rstag_5to5_bb0_cmp_i_valid_out_0 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_1 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_2 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_3 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG));
assign local_bb0_cmp_i_stall_in = (|rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_5to5_bb0_cmp_i_stall_local)
			begin
				if (~(rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb0_cmp_i_inputs_ready;
				end
			end
			else
			begin
				rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG <= local_bb0_cmp_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_0)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_1)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_2)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_3)) & rstag_5to5_bb0_cmp_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_conv22_i_inputs_ready;
 reg local_bb0_conv22_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_conv22_i_valid_out_NO_SHIFT_REG;
wire local_bb0_conv22_i_stall_in;
wire local_bb0_conv22_i_output_regs_ready;
 reg [31:0] local_bb0_conv22_i_NO_SHIFT_REG;
wire local_bb0_conv22_i_causedstall;

assign local_bb0_conv22_i_inputs_ready = rstag_5to5_bb0_cmp_i_valid_out_0;
assign local_bb0_conv22_i_output_regs_ready = (~(local_bb0_conv22_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_conv22_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_conv22_i_stall_in))));
assign rstag_5to5_bb0_cmp_i_stall_in_0 = (~(local_bb0_conv22_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_conv22_i_output_regs_ready) | ~(local_bb0_conv22_i_inputs_ready)));
assign local_bb0_conv22_i_causedstall = (local_bb0_conv22_i_inputs_ready && (~(local_bb0_conv22_i_output_regs_ready) && !(~(local_bb0_conv22_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_conv22_i_NO_SHIFT_REG <= 'x;
		local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_conv22_i_NO_SHIFT_REG <= 'x;
			local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_conv22_i_output_regs_ready)
			begin
				local_bb0_conv22_i_NO_SHIFT_REG <= rstag_5to5_bb0_cmp_i;
				local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= local_bb0_conv22_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_conv22_i_stall_in))
				begin
					local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= local_bb0_conv22_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_conv22_i_inputs_ready)
			begin
				local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__7_i_inputs_ready;
 reg local_bb0__7_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__7_i_valid_out_NO_SHIFT_REG;
wire local_bb0__7_i_stall_in;
wire local_bb0__7_i_output_regs_ready;
 reg local_bb0__7_i_NO_SHIFT_REG;
wire local_bb0__7_i_causedstall;

assign local_bb0__7_i_inputs_ready = (local_bb0_not_cmp10_i_valid_out & rstag_5to5_bb0_cmp_i_valid_out_1);
assign local_bb0__7_i_output_regs_ready = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__7_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__7_i_stall_in))));
assign local_bb0_not_cmp10_i_stall_in = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__7_i_output_regs_ready) | ~(local_bb0__7_i_inputs_ready)));
assign rstag_5to5_bb0_cmp_i_stall_in_1 = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__7_i_output_regs_ready) | ~(local_bb0__7_i_inputs_ready)));
assign local_bb0__7_i_causedstall = (local_bb0__7_i_inputs_ready && (~(local_bb0__7_i_output_regs_ready) && !(~(local_bb0__7_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__7_i_NO_SHIFT_REG <= 'x;
		local_bb0__7_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__7_i_NO_SHIFT_REG <= 'x;
			local_bb0__7_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__7_i_output_regs_ready)
			begin
				local_bb0__7_i_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i | local_bb0_not_cmp10_i);
				local_bb0__7_i_valid_out_NO_SHIFT_REG <= local_bb0__7_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__7_i_stall_in))
				begin
					local_bb0__7_i_valid_out_NO_SHIFT_REG <= local_bb0__7_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__7_i_inputs_ready)
			begin
				local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_not_cmp_i_valid_out;
wire local_bb0_not_cmp_i_stall_in;
wire local_bb0_not_cmp_i_inputs_ready;
wire local_bb0_not_cmp_i_stall_local;
wire local_bb0_not_cmp_i;

assign local_bb0_not_cmp_i_inputs_ready = rstag_5to5_bb0_cmp_i_valid_out_2;
assign local_bb0_not_cmp_i = (rstag_5to5_bb0_cmp_i ^ 1'b1);
assign local_bb0_not_cmp_i_valid_out = local_bb0_not_cmp_i_inputs_ready;
assign local_bb0_not_cmp_i_stall_local = local_bb0_not_cmp_i_stall_in;
assign rstag_5to5_bb0_cmp_i_stall_in_2 = (|local_bb0_not_cmp_i_stall_local);

// This section implements a registered operation.
// 
wire local_bb0___i_inputs_ready;
 reg local_bb0___i_wii_reg_NO_SHIFT_REG;
 reg local_bb0___i_valid_out_0_NO_SHIFT_REG;
wire local_bb0___i_stall_in_0;
 reg local_bb0___i_valid_out_1_NO_SHIFT_REG;
wire local_bb0___i_stall_in_1;
wire local_bb0___i_output_regs_ready;
 reg local_bb0___i_NO_SHIFT_REG;
wire local_bb0___i_causedstall;

assign local_bb0___i_inputs_ready = (local_bb0_lnot6_i_valid_out_NO_SHIFT_REG & rstag_5to5_bb0_cmp_i_valid_out_3);
assign local_bb0___i_output_regs_ready = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0___i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0___i_stall_in_0)) & (~(local_bb0___i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0___i_stall_in_1))));
assign local_bb0_lnot6_i_stall_in = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & (~(local_bb0___i_output_regs_ready) | ~(local_bb0___i_inputs_ready)));
assign rstag_5to5_bb0_cmp_i_stall_in_3 = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & (~(local_bb0___i_output_regs_ready) | ~(local_bb0___i_inputs_ready)));
assign local_bb0___i_causedstall = (local_bb0___i_inputs_ready && (~(local_bb0___i_output_regs_ready) && !(~(local_bb0___i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0___i_NO_SHIFT_REG <= 'x;
		local_bb0___i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0___i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0___i_NO_SHIFT_REG <= 'x;
			local_bb0___i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0___i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0___i_output_regs_ready)
			begin
				local_bb0___i_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i & local_bb0_lnot6_i_NO_SHIFT_REG);
				local_bb0___i_valid_out_0_NO_SHIFT_REG <= local_bb0___i_inputs_ready;
				local_bb0___i_valid_out_1_NO_SHIFT_REG <= local_bb0___i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0___i_stall_in_0))
				begin
					local_bb0___i_valid_out_0_NO_SHIFT_REG <= local_bb0___i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0___i_stall_in_1))
				begin
					local_bb0___i_valid_out_1_NO_SHIFT_REG <= local_bb0___i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0___i_inputs_ready)
			begin
				local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_6to6_bb0__7_i_valid_out_0;
wire rstag_6to6_bb0__7_i_stall_in_0;
wire rstag_6to6_bb0__7_i_valid_out_1;
wire rstag_6to6_bb0__7_i_stall_in_1;
wire rstag_6to6_bb0__7_i_inputs_ready;
wire rstag_6to6_bb0__7_i_stall_local;
 reg rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG;
wire rstag_6to6_bb0__7_i_combined_valid;
 reg rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG;
wire rstag_6to6_bb0__7_i;
 reg rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG;
 reg rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG;

assign rstag_6to6_bb0__7_i_inputs_ready = local_bb0__7_i_valid_out_NO_SHIFT_REG;
assign rstag_6to6_bb0__7_i = (rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG ? rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG : local_bb0__7_i_NO_SHIFT_REG);
assign rstag_6to6_bb0__7_i_combined_valid = (rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG | rstag_6to6_bb0__7_i_inputs_ready);
assign rstag_6to6_bb0__7_i_stall_local = ((rstag_6to6_bb0__7_i_stall_in_0 & ~(rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG)) | (rstag_6to6_bb0__7_i_stall_in_1 & ~(rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG)));
assign rstag_6to6_bb0__7_i_valid_out_0 = (rstag_6to6_bb0__7_i_combined_valid & ~(rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG));
assign rstag_6to6_bb0__7_i_valid_out_1 = (rstag_6to6_bb0__7_i_combined_valid & ~(rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__7_i_stall_in = (|rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_6to6_bb0__7_i_stall_local)
			begin
				if (~(rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= rstag_6to6_bb0__7_i_inputs_ready;
				end
			end
			else
			begin
				rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG <= local_bb0__7_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= (rstag_6to6_bb0__7_i_combined_valid & (rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG | ~(rstag_6to6_bb0__7_i_stall_in_0)) & rstag_6to6_bb0__7_i_stall_local);
			rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= (rstag_6to6_bb0__7_i_combined_valid & (rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG | ~(rstag_6to6_bb0__7_i_stall_in_1)) & rstag_6to6_bb0__7_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__4_i_inputs_ready;
 reg local_bb0__4_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__4_i_valid_out_NO_SHIFT_REG;
wire local_bb0__4_i_stall_in;
wire local_bb0__4_i_output_regs_ready;
 reg local_bb0__4_i_NO_SHIFT_REG;
wire local_bb0__4_i_causedstall;

assign local_bb0__4_i_inputs_ready = (local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG & local_bb0_not_cmp_i_valid_out);
assign local_bb0__4_i_output_regs_ready = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__4_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__4_i_stall_in))));
assign local_bb0_cmp10_i_stall_in_0 = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__4_i_output_regs_ready) | ~(local_bb0__4_i_inputs_ready)));
assign local_bb0_not_cmp_i_stall_in = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__4_i_output_regs_ready) | ~(local_bb0__4_i_inputs_ready)));
assign local_bb0__4_i_causedstall = (local_bb0__4_i_inputs_ready && (~(local_bb0__4_i_output_regs_ready) && !(~(local_bb0__4_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__4_i_NO_SHIFT_REG <= 'x;
		local_bb0__4_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__4_i_NO_SHIFT_REG <= 'x;
			local_bb0__4_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__4_i_output_regs_ready)
			begin
				local_bb0__4_i_NO_SHIFT_REG <= (local_bb0_cmp10_i_NO_SHIFT_REG & local_bb0_not_cmp_i);
				local_bb0__4_i_valid_out_NO_SHIFT_REG <= local_bb0__4_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__4_i_stall_in))
				begin
					local_bb0__4_i_valid_out_NO_SHIFT_REG <= local_bb0__4_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__4_i_inputs_ready)
			begin
				local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_conv44_i_stall_local;
wire [31:0] local_bb0_conv44_i;

assign local_bb0_conv44_i[31:1] = 31'h0;
assign local_bb0_conv44_i[0] = local_bb0___i_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb0_cond50_i_stall_local;
wire [31:0] local_bb0_cond50_i;

assign local_bb0_cond50_i = (local_bb0___i_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements a registered operation.
// 
wire local_bb0__12_i_inputs_ready;
 reg local_bb0__12_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__12_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0__12_i_stall_in_0;
 reg local_bb0__12_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0__12_i_stall_in_1;
wire local_bb0__12_i_output_regs_ready;
 reg local_bb0__12_i_NO_SHIFT_REG;
wire local_bb0__12_i_causedstall;

assign local_bb0__12_i_inputs_ready = rstag_6to6_bb0__7_i_valid_out_0;
assign local_bb0__12_i_output_regs_ready = (~(local_bb0__12_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0__12_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0__12_i_stall_in_0)) & (~(local_bb0__12_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0__12_i_stall_in_1))));
assign rstag_6to6_bb0__7_i_stall_in_0 = (~(local_bb0__12_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__12_i_output_regs_ready) | ~(local_bb0__12_i_inputs_ready)));
assign local_bb0__12_i_causedstall = (local_bb0__12_i_inputs_ready && (~(local_bb0__12_i_output_regs_ready) && !(~(local_bb0__12_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__12_i_NO_SHIFT_REG <= 'x;
		local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__12_i_NO_SHIFT_REG <= 'x;
			local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__12_i_output_regs_ready)
			begin
				local_bb0__12_i_NO_SHIFT_REG <= (1'b0 & rstag_6to6_bb0__7_i);
				local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= local_bb0__12_i_inputs_ready;
				local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= local_bb0__12_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__12_i_stall_in_0))
				begin
					local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= local_bb0__12_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0__12_i_stall_in_1))
				begin
					local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= local_bb0__12_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__12_i_inputs_ready)
			begin
				local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__8_i_inputs_ready;
 reg local_bb0__8_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__8_i_valid_out_NO_SHIFT_REG;
wire local_bb0__8_i_stall_in;
wire local_bb0__8_i_output_regs_ready;
 reg local_bb0__8_i_NO_SHIFT_REG;
wire local_bb0__8_i_causedstall;

assign local_bb0__8_i_inputs_ready = rstag_6to6_bb0__7_i_valid_out_1;
assign local_bb0__8_i_output_regs_ready = (~(local_bb0__8_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__8_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__8_i_stall_in))));
assign rstag_6to6_bb0__7_i_stall_in_1 = (~(local_bb0__8_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__8_i_output_regs_ready) | ~(local_bb0__8_i_inputs_ready)));
assign local_bb0__8_i_causedstall = (local_bb0__8_i_inputs_ready && (~(local_bb0__8_i_output_regs_ready) && !(~(local_bb0__8_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__8_i_NO_SHIFT_REG <= 'x;
		local_bb0__8_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__8_i_NO_SHIFT_REG <= 'x;
			local_bb0__8_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__8_i_output_regs_ready)
			begin
				local_bb0__8_i_NO_SHIFT_REG <= (1'b1 & rstag_6to6_bb0__7_i);
				local_bb0__8_i_valid_out_NO_SHIFT_REG <= local_bb0__8_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__8_i_stall_in))
				begin
					local_bb0__8_i_valid_out_NO_SHIFT_REG <= local_bb0__8_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__8_i_inputs_ready)
			begin
				local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_7to7_bb0__4_i_valid_out_0;
wire rstag_7to7_bb0__4_i_stall_in_0;
wire rstag_7to7_bb0__4_i_valid_out_1;
wire rstag_7to7_bb0__4_i_stall_in_1;
wire rstag_7to7_bb0__4_i_inputs_ready;
wire rstag_7to7_bb0__4_i_stall_local;
 reg rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG;
wire rstag_7to7_bb0__4_i_combined_valid;
 reg rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG;
wire rstag_7to7_bb0__4_i;
 reg rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG;
 reg rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG;

assign rstag_7to7_bb0__4_i_inputs_ready = local_bb0__4_i_valid_out_NO_SHIFT_REG;
assign rstag_7to7_bb0__4_i = (rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG ? rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG : local_bb0__4_i_NO_SHIFT_REG);
assign rstag_7to7_bb0__4_i_combined_valid = (rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG | rstag_7to7_bb0__4_i_inputs_ready);
assign rstag_7to7_bb0__4_i_stall_local = ((rstag_7to7_bb0__4_i_stall_in_0 & ~(rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG)) | (rstag_7to7_bb0__4_i_stall_in_1 & ~(rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG)));
assign rstag_7to7_bb0__4_i_valid_out_0 = (rstag_7to7_bb0__4_i_combined_valid & ~(rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG));
assign rstag_7to7_bb0__4_i_valid_out_1 = (rstag_7to7_bb0__4_i_combined_valid & ~(rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__4_i_stall_in = (|rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_7to7_bb0__4_i_stall_local)
			begin
				if (~(rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= rstag_7to7_bb0__4_i_inputs_ready;
				end
			end
			else
			begin
				rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG <= local_bb0__4_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= (rstag_7to7_bb0__4_i_combined_valid & (rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG | ~(rstag_7to7_bb0__4_i_stall_in_0)) & rstag_7to7_bb0__4_i_stall_local);
			rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= (rstag_7to7_bb0__4_i_combined_valid & (rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG | ~(rstag_7to7_bb0__4_i_stall_in_1)) & rstag_7to7_bb0__4_i_stall_local);
		end
	end
end


// This section implements a staging register.
// 
wire rstag_7to7_bb0__8_i_valid_out_0;
wire rstag_7to7_bb0__8_i_stall_in_0;
wire rstag_7to7_bb0__8_i_valid_out_1;
wire rstag_7to7_bb0__8_i_stall_in_1;
wire rstag_7to7_bb0__8_i_inputs_ready;
wire rstag_7to7_bb0__8_i_stall_local;
 reg rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG;
wire rstag_7to7_bb0__8_i_combined_valid;
 reg rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG;
wire rstag_7to7_bb0__8_i;
 reg rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG;
 reg rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG;

assign rstag_7to7_bb0__8_i_inputs_ready = local_bb0__8_i_valid_out_NO_SHIFT_REG;
assign rstag_7to7_bb0__8_i = (rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG ? rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG : local_bb0__8_i_NO_SHIFT_REG);
assign rstag_7to7_bb0__8_i_combined_valid = (rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG | rstag_7to7_bb0__8_i_inputs_ready);
assign rstag_7to7_bb0__8_i_stall_local = ((rstag_7to7_bb0__8_i_stall_in_0 & ~(rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG)) | (rstag_7to7_bb0__8_i_stall_in_1 & ~(rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG)));
assign rstag_7to7_bb0__8_i_valid_out_0 = (rstag_7to7_bb0__8_i_combined_valid & ~(rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG));
assign rstag_7to7_bb0__8_i_valid_out_1 = (rstag_7to7_bb0__8_i_combined_valid & ~(rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__8_i_stall_in = (|rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_7to7_bb0__8_i_stall_local)
			begin
				if (~(rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= rstag_7to7_bb0__8_i_inputs_ready;
				end
			end
			else
			begin
				rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG <= local_bb0__8_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i_combined_valid & (rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG | ~(rstag_7to7_bb0__8_i_stall_in_0)) & rstag_7to7_bb0__8_i_stall_local);
			rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i_combined_valid & (rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG | ~(rstag_7to7_bb0__8_i_stall_in_1)) & rstag_7to7_bb0__8_i_stall_local);
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0__17_i_stall_local;
wire [31:0] local_bb0__17_i;

assign local_bb0__17_i = (rstag_7to7_bb0__4_i ? 32'h0 : 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb0__5_i_valid_out;
wire local_bb0__5_i_stall_in;
wire local_bb0__5_i_inputs_ready;
wire local_bb0__5_i_stall_local;
wire [31:0] local_bb0__5_i;

assign local_bb0__5_i_inputs_ready = rstag_7to7_bb0__4_i_valid_out_1;
assign local_bb0__5_i[31:1] = 31'h0;
assign local_bb0__5_i[0] = rstag_7to7_bb0__4_i;
assign local_bb0__5_i_valid_out = local_bb0__5_i_inputs_ready;
assign local_bb0__5_i_stall_local = local_bb0__5_i_stall_in;
assign rstag_7to7_bb0__4_i_stall_in_1 = (|local_bb0__5_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0__18_i_valid_out;
wire local_bb0__18_i_stall_in;
wire local_bb0__18_i_inputs_ready;
wire local_bb0__18_i_stall_local;
wire [31:0] local_bb0__18_i;

assign local_bb0__18_i_inputs_ready = (rstag_7to7_bb0__4_i_valid_out_0 & rstag_7to7_bb0__8_i_valid_out_0);
assign local_bb0__18_i = (rstag_7to7_bb0__8_i ? 32'h1 : (local_bb0__17_i & 32'h100));
assign local_bb0__18_i_valid_out = local_bb0__18_i_inputs_ready;
assign local_bb0__18_i_stall_local = local_bb0__18_i_stall_in;
assign rstag_7to7_bb0__4_i_stall_in_0 = (local_bb0__18_i_stall_local | ~(local_bb0__18_i_inputs_ready));
assign rstag_7to7_bb0__8_i_stall_in_0 = (local_bb0__18_i_stall_local | ~(local_bb0__18_i_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb0__9_i_inputs_ready;
 reg local_bb0__9_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__9_i_valid_out_NO_SHIFT_REG;
wire local_bb0__9_i_stall_in;
wire local_bb0__9_i_output_regs_ready;
 reg [31:0] local_bb0__9_i_NO_SHIFT_REG;
wire local_bb0__9_i_causedstall;

assign local_bb0__9_i_inputs_ready = (local_bb0__5_i_valid_out & rstag_7to7_bb0__8_i_valid_out_1);
assign local_bb0__9_i_output_regs_ready = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__9_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__9_i_stall_in))));
assign local_bb0__5_i_stall_in = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__9_i_output_regs_ready) | ~(local_bb0__9_i_inputs_ready)));
assign rstag_7to7_bb0__8_i_stall_in_1 = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__9_i_output_regs_ready) | ~(local_bb0__9_i_inputs_ready)));
assign local_bb0__9_i_causedstall = (local_bb0__9_i_inputs_ready && (~(local_bb0__9_i_output_regs_ready) && !(~(local_bb0__9_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__9_i_NO_SHIFT_REG <= 'x;
		local_bb0__9_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__9_i_NO_SHIFT_REG <= 'x;
			local_bb0__9_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__9_i_output_regs_ready)
			begin
				local_bb0__9_i_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i ? 32'h0 : (local_bb0__5_i & 32'h1));
				local_bb0__9_i_valid_out_NO_SHIFT_REG <= local_bb0__9_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__9_i_stall_in))
				begin
					local_bb0__9_i_valid_out_NO_SHIFT_REG <= local_bb0__9_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__9_i_inputs_ready)
			begin
				local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__19_i_inputs_ready;
 reg local_bb0__19_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__19_i_valid_out_NO_SHIFT_REG;
wire local_bb0__19_i_stall_in;
wire local_bb0__19_i_output_regs_ready;
 reg [31:0] local_bb0__19_i_NO_SHIFT_REG;
wire local_bb0__19_i_causedstall;

assign local_bb0__19_i_inputs_ready = (local_bb0__12_i_valid_out_1_NO_SHIFT_REG & local_bb0__18_i_valid_out);
assign local_bb0__19_i_output_regs_ready = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__19_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__19_i_stall_in))));
assign local_bb0__12_i_stall_in_1 = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__19_i_output_regs_ready) | ~(local_bb0__19_i_inputs_ready)));
assign local_bb0__18_i_stall_in = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__19_i_output_regs_ready) | ~(local_bb0__19_i_inputs_ready)));
assign local_bb0__19_i_causedstall = (local_bb0__19_i_inputs_ready && (~(local_bb0__19_i_output_regs_ready) && !(~(local_bb0__19_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__19_i_NO_SHIFT_REG <= 'x;
		local_bb0__19_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__19_i_NO_SHIFT_REG <= 'x;
			local_bb0__19_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__19_i_output_regs_ready)
			begin
				local_bb0__19_i_NO_SHIFT_REG <= ((local_bb0__12_i_NO_SHIFT_REG & 1'b0) ? 32'hFFFFFF00 : (local_bb0__18_i & 32'h101));
				local_bb0__19_i_valid_out_NO_SHIFT_REG <= local_bb0__19_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__19_i_stall_in))
				begin
					local_bb0__19_i_valid_out_NO_SHIFT_REG <= local_bb0__19_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__19_i_inputs_ready)
			begin
				local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0__13_i_valid_out;
wire local_bb0__13_i_stall_in;
wire local_bb0__13_i_inputs_ready;
wire local_bb0__13_i_stall_local;
wire [31:0] local_bb0__13_i;

assign local_bb0__13_i_inputs_ready = (local_bb0__12_i_valid_out_0_NO_SHIFT_REG & local_bb0__9_i_valid_out_NO_SHIFT_REG);
assign local_bb0__13_i = ((local_bb0__12_i_NO_SHIFT_REG & 1'b0) ? 32'h0 : (local_bb0__9_i_NO_SHIFT_REG & 32'h1));
assign local_bb0__13_i_valid_out = local_bb0__13_i_inputs_ready;
assign local_bb0__13_i_stall_local = local_bb0__13_i_stall_in;
assign local_bb0__12_i_stall_in_0 = (local_bb0__13_i_stall_local | ~(local_bb0__13_i_inputs_ready));
assign local_bb0__9_i_stall_in = (local_bb0__13_i_stall_local | ~(local_bb0__13_i_inputs_ready));

// This section implements a staging register.
// 
wire rstag_8to8_bb0__19_i_valid_out_0;
wire rstag_8to8_bb0__19_i_stall_in_0;
wire rstag_8to8_bb0__19_i_valid_out_1;
wire rstag_8to8_bb0__19_i_stall_in_1;
wire rstag_8to8_bb0__19_i_inputs_ready;
wire rstag_8to8_bb0__19_i_stall_local;
 reg rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG;
wire rstag_8to8_bb0__19_i_combined_valid;
 reg [31:0] rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_8to8_bb0__19_i;
 reg rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG;
 reg rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG;

assign rstag_8to8_bb0__19_i_inputs_ready = local_bb0__19_i_valid_out_NO_SHIFT_REG;
assign rstag_8to8_bb0__19_i = (rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG ? rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG : (local_bb0__19_i_NO_SHIFT_REG & 32'hFFFFFF01));
assign rstag_8to8_bb0__19_i_combined_valid = (rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG | rstag_8to8_bb0__19_i_inputs_ready);
assign rstag_8to8_bb0__19_i_stall_local = ((rstag_8to8_bb0__19_i_stall_in_0 & ~(rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG)) | (rstag_8to8_bb0__19_i_stall_in_1 & ~(rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG)));
assign rstag_8to8_bb0__19_i_valid_out_0 = (rstag_8to8_bb0__19_i_combined_valid & ~(rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG));
assign rstag_8to8_bb0__19_i_valid_out_1 = (rstag_8to8_bb0__19_i_combined_valid & ~(rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__19_i_stall_in = (|rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_8to8_bb0__19_i_stall_local)
			begin
				if (~(rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= rstag_8to8_bb0__19_i_inputs_ready;
				end
			end
			else
			begin
				rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG <= (local_bb0__19_i_NO_SHIFT_REG & 32'hFFFFFF01);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= (rstag_8to8_bb0__19_i_combined_valid & (rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG | ~(rstag_8to8_bb0__19_i_stall_in_0)) & rstag_8to8_bb0__19_i_stall_local);
			rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= (rstag_8to8_bb0__19_i_combined_valid & (rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG | ~(rstag_8to8_bb0__19_i_stall_in_1)) & rstag_8to8_bb0__19_i_stall_local);
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_fold_i_valid_out;
wire local_bb0_fold_i_stall_in;
wire local_bb0_fold_i_inputs_ready;
wire local_bb0_fold_i_stall_local;
wire [31:0] local_bb0_fold_i;

assign local_bb0_fold_i_inputs_ready = (local_bb0_shr_i_valid_out_1_NO_SHIFT_REG & rstag_8to8_bb0__19_i_valid_out_0);
assign local_bb0_fold_i = ((rstag_8to8_bb0__19_i & 32'hFFFFFF01) + (local_bb0_shr_i_NO_SHIFT_REG & 32'h1FF));
assign local_bb0_fold_i_valid_out = local_bb0_fold_i_inputs_ready;
assign local_bb0_fold_i_stall_local = local_bb0_fold_i_stall_in;
assign local_bb0_shr_i_stall_in_1 = (local_bb0_fold_i_stall_local | ~(local_bb0_fold_i_inputs_ready));
assign rstag_8to8_bb0__19_i_stall_in_0 = (local_bb0_fold_i_stall_local | ~(local_bb0_fold_i_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb0_add_i_inputs_ready;
 reg local_bb0_add_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_add_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_add_i_stall_in_0;
 reg local_bb0_add_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_add_i_stall_in_1;
wire local_bb0_add_i_output_regs_ready;
 reg [31:0] local_bb0_add_i_NO_SHIFT_REG;
wire local_bb0_add_i_causedstall;

assign local_bb0_add_i_inputs_ready = (rstag_8to8_bb0__19_i_valid_out_1 & rstag_4to4_bb0_and1_i_valid_out_0);
assign local_bb0_add_i_output_regs_ready = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_add_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_add_i_stall_in_0)) & (~(local_bb0_add_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_add_i_stall_in_1))));
assign rstag_8to8_bb0__19_i_stall_in_1 = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_add_i_output_regs_ready) | ~(local_bb0_add_i_inputs_ready)));
assign rstag_4to4_bb0_and1_i_stall_in_0 = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_add_i_output_regs_ready) | ~(local_bb0_add_i_inputs_ready)));
assign local_bb0_add_i_causedstall = (local_bb0_add_i_inputs_ready && (~(local_bb0_add_i_output_regs_ready) && !(~(local_bb0_add_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add_i_NO_SHIFT_REG <= 'x;
		local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add_i_NO_SHIFT_REG <= 'x;
			local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add_i_output_regs_ready)
			begin
				local_bb0_add_i_NO_SHIFT_REG <= ((rstag_8to8_bb0__19_i & 32'hFFFFFF01) + (rstag_4to4_bb0_and1_i & 32'hFF));
				local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= local_bb0_add_i_inputs_ready;
				local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= local_bb0_add_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_add_i_stall_in_0))
				begin
					local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= local_bb0_add_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_add_i_stall_in_1))
				begin
					local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= local_bb0_add_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add_i_inputs_ready)
			begin
				local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and32_i_inputs_ready;
 reg local_bb0_and32_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and32_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and32_i_stall_in;
wire local_bb0_and32_i_output_regs_ready;
 reg [31:0] local_bb0_and32_i_NO_SHIFT_REG;
wire local_bb0_and32_i_causedstall;

assign local_bb0_and32_i_inputs_ready = local_bb0_fold_i_valid_out;
assign local_bb0_and32_i_output_regs_ready = (~(local_bb0_and32_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and32_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and32_i_stall_in))));
assign local_bb0_fold_i_stall_in = (~(local_bb0_and32_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and32_i_output_regs_ready) | ~(local_bb0_and32_i_inputs_ready)));
assign local_bb0_and32_i_causedstall = (local_bb0_and32_i_inputs_ready && (~(local_bb0_and32_i_output_regs_ready) && !(~(local_bb0_and32_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and32_i_NO_SHIFT_REG <= 'x;
		local_bb0_and32_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and32_i_NO_SHIFT_REG <= 'x;
			local_bb0_and32_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and32_i_output_regs_ready)
			begin
				local_bb0_and32_i_NO_SHIFT_REG <= (local_bb0_fold_i << 32'h17);
				local_bb0_and32_i_valid_out_NO_SHIFT_REG <= local_bb0_and32_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and32_i_stall_in))
				begin
					local_bb0_and32_i_valid_out_NO_SHIFT_REG <= local_bb0_and32_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and32_i_inputs_ready)
			begin
				local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_cmp20_i_stall_local;
wire local_bb0_cmp20_i;

assign local_bb0_cmp20_i = ($signed(local_bb0_add_i_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb0_cmp25_i_stall_local;
wire local_bb0_cmp25_i;

assign local_bb0_cmp25_i = ($signed(local_bb0_add_i_NO_SHIFT_REG) < $signed(32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_shl_i_stall_local;
wire [31:0] local_bb0_shl_i;

assign local_bb0_shl_i = ((local_bb0_and32_i_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb0_conv_i_valid_out;
wire local_bb0_conv_i_stall_in;
wire local_bb0_conv_i_inputs_ready;
wire local_bb0_conv_i_stall_local;
wire [31:0] local_bb0_conv_i;

assign local_bb0_conv_i_inputs_ready = local_bb0_add_i_valid_out_0_NO_SHIFT_REG;
assign local_bb0_conv_i[31:1] = 31'h0;
assign local_bb0_conv_i[0] = local_bb0_cmp20_i;
assign local_bb0_conv_i_valid_out = local_bb0_conv_i_inputs_ready;
assign local_bb0_conv_i_stall_local = local_bb0_conv_i_stall_in;
assign local_bb0_add_i_stall_in_0 = (|local_bb0_conv_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0_conv26_i_valid_out;
wire local_bb0_conv26_i_stall_in;
wire local_bb0_conv26_i_inputs_ready;
wire local_bb0_conv26_i_stall_local;
wire [31:0] local_bb0_conv26_i;

assign local_bb0_conv26_i_inputs_ready = local_bb0_add_i_valid_out_1_NO_SHIFT_REG;
assign local_bb0_conv26_i[31:1] = 31'h0;
assign local_bb0_conv26_i[0] = local_bb0_cmp25_i;
assign local_bb0_conv26_i_valid_out = local_bb0_conv26_i_inputs_ready;
assign local_bb0_conv26_i_stall_local = local_bb0_conv26_i_stall_in;
assign local_bb0_add_i_stall_in_1 = (|local_bb0_conv26_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0_or34_i_stall_local;
wire [31:0] local_bb0_or34_i;

assign local_bb0_or34_i = ((local_bb0_shl_i & 32'h7F800000) | (local_bb0_and33_i_NO_SHIFT_REG & 32'h807FFFFF));

// This section implements a registered operation.
// 
wire local_bb0_or_i_inputs_ready;
 reg local_bb0_or_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_or_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_or_i_stall_in_0;
 reg local_bb0_or_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_or_i_stall_in_1;
wire local_bb0_or_i_output_regs_ready;
 reg [31:0] local_bb0_or_i_NO_SHIFT_REG;
wire local_bb0_or_i_causedstall;

assign local_bb0_or_i_inputs_ready = (local_bb0_conv_i_valid_out & local_bb0_conv22_i_valid_out_NO_SHIFT_REG);
assign local_bb0_or_i_output_regs_ready = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_or_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_or_i_stall_in_0)) & (~(local_bb0_or_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_or_i_stall_in_1))));
assign local_bb0_conv_i_stall_in = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or_i_output_regs_ready) | ~(local_bb0_or_i_inputs_ready)));
assign local_bb0_conv22_i_stall_in = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or_i_output_regs_ready) | ~(local_bb0_or_i_inputs_ready)));
assign local_bb0_or_i_causedstall = (local_bb0_or_i_inputs_ready && (~(local_bb0_or_i_output_regs_ready) && !(~(local_bb0_or_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or_i_NO_SHIFT_REG <= 'x;
		local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or_i_NO_SHIFT_REG <= 'x;
			local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or_i_output_regs_ready)
			begin
				local_bb0_or_i_NO_SHIFT_REG <= ((local_bb0_conv_i & 32'h1) | (local_bb0_conv22_i_NO_SHIFT_REG & 32'h1));
				local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= local_bb0_or_i_inputs_ready;
				local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= local_bb0_or_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_or_i_stall_in_0))
				begin
					local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= local_bb0_or_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_or_i_stall_in_1))
				begin
					local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= local_bb0_or_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or_i_inputs_ready)
			begin
				local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_or29_i_inputs_ready;
 reg local_bb0_or29_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_or29_i_valid_out_NO_SHIFT_REG;
wire local_bb0_or29_i_stall_in;
wire local_bb0_or29_i_output_regs_ready;
 reg [31:0] local_bb0_or29_i_NO_SHIFT_REG;
wire local_bb0_or29_i_causedstall;

assign local_bb0_or29_i_inputs_ready = (local_bb0_conv26_i_valid_out & local_bb0__13_i_valid_out);
assign local_bb0_or29_i_output_regs_ready = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_or29_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_or29_i_stall_in))));
assign local_bb0_conv26_i_stall_in = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or29_i_output_regs_ready) | ~(local_bb0_or29_i_inputs_ready)));
assign local_bb0__13_i_stall_in = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or29_i_output_regs_ready) | ~(local_bb0_or29_i_inputs_ready)));
assign local_bb0_or29_i_causedstall = (local_bb0_or29_i_inputs_ready && (~(local_bb0_or29_i_output_regs_ready) && !(~(local_bb0_or29_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or29_i_NO_SHIFT_REG <= 'x;
		local_bb0_or29_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or29_i_NO_SHIFT_REG <= 'x;
			local_bb0_or29_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or29_i_output_regs_ready)
			begin
				local_bb0_or29_i_NO_SHIFT_REG <= ((local_bb0_conv26_i & 32'h1) | (local_bb0__13_i & 32'h1));
				local_bb0_or29_i_valid_out_NO_SHIFT_REG <= local_bb0_or29_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_or29_i_stall_in))
				begin
					local_bb0_or29_i_valid_out_NO_SHIFT_REG <= local_bb0_or29_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or29_i_inputs_ready)
			begin
				local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_or45_i_stall_local;
wire [31:0] local_bb0_or45_i;

assign local_bb0_or45_i = ((local_bb0_or_i_NO_SHIFT_REG & 32'h1) | (local_bb0_conv44_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_or39_i_stall_local;
wire [31:0] local_bb0_or39_i;

assign local_bb0_or39_i = ((local_bb0_or29_i_NO_SHIFT_REG & 32'h1) | (local_bb0_or_i_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_tobool46_i_stall_local;
wire local_bb0_tobool46_i;

assign local_bb0_tobool46_i = ((local_bb0_or45_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_tobool40_i_stall_local;
wire local_bb0_tobool40_i;

assign local_bb0_tobool40_i = ((local_bb0_or39_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_cond47_i_stall_local;
wire [31:0] local_bb0_cond47_i;

assign local_bb0_cond47_i = (local_bb0_tobool46_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_cond_i_stall_local;
wire [31:0] local_bb0_cond_i;

assign local_bb0_cond_i = (local_bb0_tobool40_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb0_or52_i_stall_local;
wire [31:0] local_bb0_or52_i;

assign local_bb0_or52_i = ((local_bb0_cond47_i & 32'h7F800000) | (local_bb0_cond50_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb0_and51_i_stall_local;
wire [31:0] local_bb0_and51_i;

assign local_bb0_and51_i = ((local_bb0_cond_i | 32'h80000000) & local_bb0_or34_i);

// This section implements an unregistered operation.
// 
wire local_bb0_or53_i_stall_local;
wire [31:0] local_bb0_or53_i;

assign local_bb0_or53_i = ((local_bb0_or52_i & 32'h7FC00000) | local_bb0_and51_i);

// This section implements an unregistered operation.
// 
wire local_bb0_var__u2_valid_out;
wire local_bb0_var__u2_stall_in;
wire local_bb0_var__u2_inputs_ready;
wire local_bb0_var__u2_stall_local;
wire [31:0] local_bb0_var__u2;

assign local_bb0_var__u2_inputs_ready = (local_bb0_and33_i_valid_out_NO_SHIFT_REG & local_bb0_and32_i_valid_out_NO_SHIFT_REG & local_bb0___i_valid_out_1_NO_SHIFT_REG & local_bb0___i_valid_out_0_NO_SHIFT_REG & local_bb0_or_i_valid_out_1_NO_SHIFT_REG & local_bb0_or29_i_valid_out_NO_SHIFT_REG & local_bb0_or_i_valid_out_0_NO_SHIFT_REG);
assign local_bb0_var__u2 = local_bb0_or53_i;
assign local_bb0_var__u2_valid_out = local_bb0_var__u2_inputs_ready;
assign local_bb0_var__u2_stall_local = local_bb0_var__u2_stall_in;
assign local_bb0_and33_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_and32_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0___i_stall_in_1 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0___i_stall_in_0 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or_i_stall_in_1 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or29_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or_i_stall_in_0 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));

// This section implements a staging register.
// 
wire rstag_10to10_bb0_var__u2_valid_out;
wire rstag_10to10_bb0_var__u2_stall_in;
wire rstag_10to10_bb0_var__u2_inputs_ready;
wire rstag_10to10_bb0_var__u2_stall_local;
 reg rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG;
wire rstag_10to10_bb0_var__u2_combined_valid;
 reg [31:0] rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_10to10_bb0_var__u2;

assign rstag_10to10_bb0_var__u2_inputs_ready = local_bb0_var__u2_valid_out;
assign rstag_10to10_bb0_var__u2 = (rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG ? rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG : local_bb0_var__u2);
assign rstag_10to10_bb0_var__u2_combined_valid = (rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG | rstag_10to10_bb0_var__u2_inputs_ready);
assign rstag_10to10_bb0_var__u2_valid_out = rstag_10to10_bb0_var__u2_combined_valid;
assign rstag_10to10_bb0_var__u2_stall_local = rstag_10to10_bb0_var__u2_stall_in;
assign local_bb0_var__u2_stall_in = (|rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_10to10_bb0_var__u2_stall_local)
			begin
				if (~(rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG))
				begin
					rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= rstag_10to10_bb0_var__u2_inputs_ready;
				end
			end
			else
			begin
				rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG))
		begin
			rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG <= local_bb0_var__u2;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_mul50_inputs_ready;
 reg local_bb0_mul50_wii_reg_NO_SHIFT_REG;
 reg local_bb0_mul50_valid_out_NO_SHIFT_REG;
wire local_bb0_mul50_stall_in;
wire local_bb0_mul50_output_regs_ready;
wire [31:0] local_bb0_mul50;
 reg local_bb0_mul50_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb0_mul50_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb0_mul50_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb0_mul50_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb0_mul50_valid_pipe_4_NO_SHIFT_REG;
wire local_bb0_mul50_causedstall;

acl_fp_mul_ll_s5 fp_module_local_bb0_mul50 (
	.clock(clock),
	.dataa(rstag_10to10_bb0_var__u2),
	.datab(input_e_d),
	.enable(local_bb0_mul50_output_regs_ready),
	.result(local_bb0_mul50)
);


assign local_bb0_mul50_inputs_ready = (merge_node_valid_out_5_NO_SHIFT_REG & rstag_10to10_bb0_var__u2_valid_out);
assign local_bb0_mul50_output_regs_ready = (~(local_bb0_mul50_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_mul50_valid_out_NO_SHIFT_REG) | ~(local_bb0_mul50_stall_in))));
assign merge_node_stall_in_5 = (~(local_bb0_mul50_wii_reg_NO_SHIFT_REG) & (~(local_bb0_mul50_output_regs_ready) | ~(local_bb0_mul50_inputs_ready)));
assign rstag_10to10_bb0_var__u2_stall_in = (~(local_bb0_mul50_wii_reg_NO_SHIFT_REG) & (~(local_bb0_mul50_output_regs_ready) | ~(local_bb0_mul50_inputs_ready)));
assign local_bb0_mul50_causedstall = (local_bb0_mul50_inputs_ready && (~(local_bb0_mul50_output_regs_ready) && !(~(local_bb0_mul50_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul50_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul50_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul50_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul50_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul50_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul50_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul50_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul50_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul50_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul50_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul50_output_regs_ready)
			begin
				local_bb0_mul50_valid_pipe_0_NO_SHIFT_REG <= local_bb0_mul50_inputs_ready;
				local_bb0_mul50_valid_pipe_1_NO_SHIFT_REG <= local_bb0_mul50_valid_pipe_0_NO_SHIFT_REG;
				local_bb0_mul50_valid_pipe_2_NO_SHIFT_REG <= local_bb0_mul50_valid_pipe_1_NO_SHIFT_REG;
				local_bb0_mul50_valid_pipe_3_NO_SHIFT_REG <= local_bb0_mul50_valid_pipe_2_NO_SHIFT_REG;
				local_bb0_mul50_valid_pipe_4_NO_SHIFT_REG <= local_bb0_mul50_valid_pipe_3_NO_SHIFT_REG;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul50_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul50_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul50_output_regs_ready)
			begin
				local_bb0_mul50_valid_out_NO_SHIFT_REG <= local_bb0_mul50_valid_pipe_4_NO_SHIFT_REG;
			end
			else
			begin
				if (~(local_bb0_mul50_stall_in))
				begin
					local_bb0_mul50_valid_out_NO_SHIFT_REG <= local_bb0_mul50_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul50_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul50_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul50_valid_pipe_4_NO_SHIFT_REG)
			begin
				local_bb0_mul50_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg lvb_bb0_cmp1622_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_sub25_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_sub29_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_mul50_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb0_var__reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb0_var__u0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb0_var__u0_valid_out_NO_SHIFT_REG & local_bb0_var__valid_out_NO_SHIFT_REG & local_bb0_mul50_valid_out_NO_SHIFT_REG & local_bb0_sub29_valid_out_NO_SHIFT_REG & local_bb0_sub25_valid_out_NO_SHIFT_REG & local_bb0_cmp1622_valid_out_NO_SHIFT_REG & merge_node_valid_out_7_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb0_var__u0_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_var__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_mul50_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_sub29_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_sub25_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_cmp1622_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign merge_node_stall_in_7 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb0_cmp1622 = lvb_bb0_cmp1622_reg_NO_SHIFT_REG;
assign lvb_bb0_sub25 = lvb_bb0_sub25_reg_NO_SHIFT_REG;
assign lvb_bb0_sub29 = lvb_bb0_sub29_reg_NO_SHIFT_REG;
assign lvb_bb0_mul50 = lvb_bb0_mul50_reg_NO_SHIFT_REG;
assign lvb_bb0_var_ = lvb_bb0_var__reg_NO_SHIFT_REG;
assign lvb_bb0_var__u0 = lvb_bb0_var__u0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0 = lvb_input_global_id_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1 = lvb_input_global_id_1_reg_NO_SHIFT_REG;
assign lvb_input_acl_hw_wg_id = lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb0_cmp1622_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_sub25_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_sub29_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_mul50_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__u0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_reg_NO_SHIFT_REG <= 'x;
		lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb0_cmp1622_reg_NO_SHIFT_REG <= local_bb0_cmp1622_NO_SHIFT_REG;
			lvb_bb0_sub25_reg_NO_SHIFT_REG <= local_bb0_sub25_NO_SHIFT_REG;
			lvb_bb0_sub29_reg_NO_SHIFT_REG <= local_bb0_sub29_NO_SHIFT_REG;
			lvb_bb0_mul50_reg_NO_SHIFT_REG <= local_bb0_mul50;
			lvb_bb0_var__reg_NO_SHIFT_REG <= local_bb0_var__NO_SHIFT_REG;
			lvb_bb0_var__u0_reg_NO_SHIFT_REG <= local_bb0_var__u0_NO_SHIFT_REG;
			lvb_input_global_id_0_reg_NO_SHIFT_REG <= local_lvm_input_global_id_0_NO_SHIFT_REG;
			lvb_input_global_id_1_reg_NO_SHIFT_REG <= local_lvm_input_global_id_1_NO_SHIFT_REG;
			lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG <= local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_1
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_global_size_0,
		input [63:0] 		input_in,
		input 		input_wii_cmp1622,
		input [31:0] 		input_wii_sub25,
		input [31:0] 		input_wii_sub29,
		input [31:0] 		input_wii_mul50,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u3,
		input 		valid_in,
		output 		stall_out,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		input [31:0] 		input_acl_hw_wg_id,
		output 		valid_out,
		input 		stall_in,
		output [63:0] 		lvb_bb1_idxprom,
		output [31:0] 		lvb_bb1_ld_,
		output 		lvb_bb1_cmp,
		output 		lvb_bb1_var_,
		output [31:0] 		lvb_input_global_id_0,
		output [31:0] 		lvb_input_global_id_1,
		output [31:0] 		lvb_input_acl_hw_wg_id,
		input [31:0] 		workgroup_size,
		input 		start,
		input [511:0] 		avm_local_bb1_ld__readdata,
		input 		avm_local_bb1_ld__readdatavalid,
		input 		avm_local_bb1_ld__waitrequest,
		output [32:0] 		avm_local_bb1_ld__address,
		output 		avm_local_bb1_ld__read,
		output 		avm_local_bb1_ld__write,
		input 		avm_local_bb1_ld__writeack,
		output [511:0] 		avm_local_bb1_ld__writedata,
		output [63:0] 		avm_local_bb1_ld__byteenable,
		output [4:0] 		avm_local_bb1_ld__burstcount,
		output 		local_bb1_ld__active,
		input 		clock2x
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_global_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_global_id_0_staging_reg_NO_SHIFT_REG <= input_global_id_0;
				input_global_id_1_staging_reg_NO_SHIFT_REG <= input_global_id_1;
				input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb1_mul_inputs_ready;
 reg local_bb1_mul_valid_out_NO_SHIFT_REG;
wire local_bb1_mul_stall_in;
wire local_bb1_mul_output_regs_ready;
wire [31:0] local_bb1_mul;
 reg local_bb1_mul_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb1_mul_valid_pipe_1_NO_SHIFT_REG;
wire local_bb1_mul_causedstall;

acl_int_mult int_module_local_bb1_mul (
	.clock(clock),
	.dataa(input_global_size_0),
	.datab(local_lvm_input_global_id_1_NO_SHIFT_REG),
	.enable(local_bb1_mul_output_regs_ready),
	.result(local_bb1_mul)
);

defparam int_module_local_bb1_mul.INPUT1_WIDTH = 32;
defparam int_module_local_bb1_mul.INPUT2_WIDTH = 32;
defparam int_module_local_bb1_mul.OUTPUT_WIDTH = 32;
defparam int_module_local_bb1_mul.LATENCY = 3;
defparam int_module_local_bb1_mul.SIGNED = 0;

assign local_bb1_mul_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb1_mul_output_regs_ready = (&(~(local_bb1_mul_valid_out_NO_SHIFT_REG) | ~(local_bb1_mul_stall_in)));
assign merge_node_stall_in_0 = (~(local_bb1_mul_output_regs_ready) | ~(local_bb1_mul_inputs_ready));
assign local_bb1_mul_causedstall = (local_bb1_mul_inputs_ready && (~(local_bb1_mul_output_regs_ready) && !(~(local_bb1_mul_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb1_mul_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul_output_regs_ready)
		begin
			local_bb1_mul_valid_pipe_0_NO_SHIFT_REG <= local_bb1_mul_inputs_ready;
			local_bb1_mul_valid_pipe_1_NO_SHIFT_REG <= local_bb1_mul_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul_output_regs_ready)
		begin
			local_bb1_mul_valid_out_NO_SHIFT_REG <= local_bb1_mul_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb1_mul_stall_in))
			begin
				local_bb1_mul_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_input_global_id_0_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_1_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;
 reg rnode_1to4_input_global_id_0_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to4_input_global_id_0_0_consumed_1_NO_SHIFT_REG;
wire [63:0] rci_rcnode_1to168_rc2_input_global_id_1_0_reg_1;

acl_data_fifo rnode_1to4_input_global_id_0_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_lvm_input_global_id_0_NO_SHIFT_REG),
	.data_out(rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign merge_node_stall_in_1 = rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG = ((rnode_1to4_input_global_id_0_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to4_input_global_id_0_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to4_input_global_id_0_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to4_input_global_id_0_0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to4_input_global_id_0_0_valid_out_0_NO_SHIFT_REG = (rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG & ~(rnode_1to4_input_global_id_0_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to4_input_global_id_0_0_valid_out_1_NO_SHIFT_REG = (rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG & ~(rnode_1to4_input_global_id_0_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to4_input_global_id_0_0_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_1_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
assign rci_rcnode_1to168_rc2_input_global_id_1_0_reg_1[31:0] = local_lvm_input_global_id_1_NO_SHIFT_REG;
assign rci_rcnode_1to168_rc2_input_global_id_1_0_reg_1[63:32] = local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to4_input_global_id_0_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to4_input_global_id_0_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to4_input_global_id_0_0_consumed_0_NO_SHIFT_REG <= (rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG & (rnode_1to4_input_global_id_0_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to4_input_global_id_0_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG);
		rnode_1to4_input_global_id_0_0_consumed_1_NO_SHIFT_REG <= (rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG & (rnode_1to4_input_global_id_0_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to4_input_global_id_0_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 167
//  * capacity = 167
 logic rcnode_1to168_rc2_input_global_id_1_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to168_rc2_input_global_id_1_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rcnode_1to168_rc2_input_global_id_1_0_NO_SHIFT_REG;
 logic rcnode_1to168_rc2_input_global_id_1_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rcnode_1to168_rc2_input_global_id_1_0_reg_168_NO_SHIFT_REG;
 logic rcnode_1to168_rc2_input_global_id_1_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rcnode_1to168_rc2_input_global_id_1_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rcnode_1to168_rc2_input_global_id_1_0_stall_out_reg_168_IP_NO_SHIFT_REG;
 logic rcnode_1to168_rc2_input_global_id_1_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rcnode_1to168_rc2_input_global_id_1_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to168_rc2_input_global_id_1_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to168_rc2_input_global_id_1_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rcnode_1to168_rc2_input_global_id_1_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rcnode_1to168_rc2_input_global_id_1_0_stall_out_reg_168_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to168_rc2_input_global_id_1_0_reg_1),
	.data_out(rcnode_1to168_rc2_input_global_id_1_0_reg_168_NO_SHIFT_REG)
);

defparam rcnode_1to168_rc2_input_global_id_1_0_reg_168_fifo.DEPTH = 168;
defparam rcnode_1to168_rc2_input_global_id_1_0_reg_168_fifo.DATA_WIDTH = 64;
defparam rcnode_1to168_rc2_input_global_id_1_0_reg_168_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to168_rc2_input_global_id_1_0_reg_168_fifo.IMPL = "ram";

assign rcnode_1to168_rc2_input_global_id_1_0_reg_168_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign rcnode_1to168_rc2_input_global_id_1_0_stall_out_reg_168_NO_SHIFT_REG = (~(rcnode_1to168_rc2_input_global_id_1_0_reg_168_inputs_ready_NO_SHIFT_REG) | rcnode_1to168_rc2_input_global_id_1_0_stall_out_reg_168_IP_NO_SHIFT_REG);
assign merge_node_stall_in_2 = rcnode_1to168_rc2_input_global_id_1_0_stall_out_reg_168_NO_SHIFT_REG;
assign rcnode_1to168_rc2_input_global_id_1_0_NO_SHIFT_REG = rcnode_1to168_rc2_input_global_id_1_0_reg_168_NO_SHIFT_REG;
assign rcnode_1to168_rc2_input_global_id_1_0_stall_in_reg_168_NO_SHIFT_REG = rcnode_1to168_rc2_input_global_id_1_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to168_rc2_input_global_id_1_0_valid_out_NO_SHIFT_REG = rcnode_1to168_rc2_input_global_id_1_0_valid_out_reg_168_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb1_add_valid_out;
wire local_bb1_add_stall_in;
wire local_bb1_add_inputs_ready;
wire local_bb1_add_stall_local;
wire [31:0] local_bb1_add;

assign local_bb1_add_inputs_ready = (local_bb1_mul_valid_out_NO_SHIFT_REG & rnode_1to4_input_global_id_0_0_valid_out_0_NO_SHIFT_REG);
assign local_bb1_add = (local_bb1_mul + rnode_1to4_input_global_id_0_0_NO_SHIFT_REG);
assign local_bb1_add_valid_out = local_bb1_add_inputs_ready;
assign local_bb1_add_stall_local = local_bb1_add_stall_in;
assign local_bb1_mul_stall_in = (local_bb1_add_stall_local | ~(local_bb1_add_inputs_ready));
assign rnode_1to4_input_global_id_0_0_stall_in_0_NO_SHIFT_REG = (local_bb1_add_stall_local | ~(local_bb1_add_inputs_ready));

// Register node:
//  * latency = 164
//  * capacity = 164
 logic rnode_4to168_input_global_id_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to168_input_global_id_0_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to168_input_global_id_0_0_NO_SHIFT_REG;
 logic rnode_4to168_input_global_id_0_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to168_input_global_id_0_0_reg_168_NO_SHIFT_REG;
 logic rnode_4to168_input_global_id_0_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_4to168_input_global_id_0_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_4to168_input_global_id_0_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_4to168_input_global_id_0_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to168_input_global_id_0_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to168_input_global_id_0_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_4to168_input_global_id_0_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_4to168_input_global_id_0_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_1to4_input_global_id_0_1_NO_SHIFT_REG),
	.data_out(rnode_4to168_input_global_id_0_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_4to168_input_global_id_0_0_reg_168_fifo.DEPTH = 165;
defparam rnode_4to168_input_global_id_0_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_4to168_input_global_id_0_0_reg_168_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to168_input_global_id_0_0_reg_168_fifo.IMPL = "ram";

assign rnode_4to168_input_global_id_0_0_reg_168_inputs_ready_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_valid_out_1_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_stall_in_1_NO_SHIFT_REG = rnode_4to168_input_global_id_0_0_stall_out_reg_168_NO_SHIFT_REG;
assign rnode_4to168_input_global_id_0_0_NO_SHIFT_REG = rnode_4to168_input_global_id_0_0_reg_168_NO_SHIFT_REG;
assign rnode_4to168_input_global_id_0_0_stall_in_reg_168_NO_SHIFT_REG = rnode_4to168_input_global_id_0_0_stall_in_NO_SHIFT_REG;
assign rnode_4to168_input_global_id_0_0_valid_out_NO_SHIFT_REG = rnode_4to168_input_global_id_0_0_valid_out_reg_168_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb1_add_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb1_add_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb1_add_0_NO_SHIFT_REG;
 logic rnode_4to5_bb1_add_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb1_add_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb1_add_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb1_add_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb1_add_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb1_add_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb1_add_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb1_add_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb1_add_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb1_add_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb1_add),
	.data_out(rnode_4to5_bb1_add_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb1_add_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb1_add_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb1_add_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb1_add_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_4to5_bb1_add_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb1_add_valid_out;
assign local_bb1_add_stall_in = rnode_4to5_bb1_add_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb1_add_0_NO_SHIFT_REG = rnode_4to5_bb1_add_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb1_add_0_stall_in_reg_5_NO_SHIFT_REG = rnode_4to5_bb1_add_0_stall_in_NO_SHIFT_REG;
assign rnode_4to5_bb1_add_0_valid_out_NO_SHIFT_REG = rnode_4to5_bb1_add_0_valid_out_reg_5_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb1_idxprom_stall_local;
wire [63:0] local_bb1_idxprom;

assign local_bb1_idxprom[63:32] = 32'h0;
assign local_bb1_idxprom[31:0] = rnode_4to5_bb1_add_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb1_idxprom_valid_out_1;
wire local_bb1_idxprom_stall_in_1;
wire local_bb1_arrayidx_valid_out;
wire local_bb1_arrayidx_stall_in;
wire local_bb1_arrayidx_inputs_ready;
wire local_bb1_arrayidx_stall_local;
wire [63:0] local_bb1_arrayidx;
 reg local_bb1_idxprom_consumed_1_NO_SHIFT_REG;
 reg local_bb1_arrayidx_consumed_0_NO_SHIFT_REG;

assign local_bb1_arrayidx_inputs_ready = rnode_4to5_bb1_add_0_valid_out_NO_SHIFT_REG;
assign local_bb1_arrayidx = ((input_in & 64'hFFFFFFFFFFFFFC00) + ((local_bb1_idxprom & 64'hFFFFFFFF) << 6'h2));
assign local_bb1_arrayidx_stall_local = ((local_bb1_idxprom_stall_in_1 & ~(local_bb1_idxprom_consumed_1_NO_SHIFT_REG)) | (local_bb1_arrayidx_stall_in & ~(local_bb1_arrayidx_consumed_0_NO_SHIFT_REG)));
assign local_bb1_idxprom_valid_out_1 = (local_bb1_arrayidx_inputs_ready & ~(local_bb1_idxprom_consumed_1_NO_SHIFT_REG));
assign local_bb1_arrayidx_valid_out = (local_bb1_arrayidx_inputs_ready & ~(local_bb1_arrayidx_consumed_0_NO_SHIFT_REG));
assign rnode_4to5_bb1_add_0_stall_in_NO_SHIFT_REG = (|local_bb1_arrayidx_stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_idxprom_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb1_arrayidx_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb1_idxprom_consumed_1_NO_SHIFT_REG <= (local_bb1_arrayidx_inputs_ready & (local_bb1_idxprom_consumed_1_NO_SHIFT_REG | ~(local_bb1_idxprom_stall_in_1)) & local_bb1_arrayidx_stall_local);
		local_bb1_arrayidx_consumed_0_NO_SHIFT_REG <= (local_bb1_arrayidx_inputs_ready & (local_bb1_arrayidx_consumed_0_NO_SHIFT_REG | ~(local_bb1_arrayidx_stall_in)) & local_bb1_arrayidx_stall_local);
	end
end


// Register node:
//  * latency = 163
//  * capacity = 163
 logic rnode_5to168_bb1_idxprom_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to168_bb1_idxprom_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_5to168_bb1_idxprom_0_NO_SHIFT_REG;
 logic rnode_5to168_bb1_idxprom_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_5to168_bb1_idxprom_0_reg_168_NO_SHIFT_REG;
 logic rnode_5to168_bb1_idxprom_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_5to168_bb1_idxprom_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_5to168_bb1_idxprom_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_5to168_bb1_idxprom_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to168_bb1_idxprom_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to168_bb1_idxprom_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_5to168_bb1_idxprom_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_5to168_bb1_idxprom_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in((local_bb1_idxprom & 64'hFFFFFFFF)),
	.data_out(rnode_5to168_bb1_idxprom_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_5to168_bb1_idxprom_0_reg_168_fifo.DEPTH = 164;
defparam rnode_5to168_bb1_idxprom_0_reg_168_fifo.DATA_WIDTH = 64;
defparam rnode_5to168_bb1_idxprom_0_reg_168_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_5to168_bb1_idxprom_0_reg_168_fifo.IMPL = "ram";

assign rnode_5to168_bb1_idxprom_0_reg_168_inputs_ready_NO_SHIFT_REG = local_bb1_idxprom_valid_out_1;
assign local_bb1_idxprom_stall_in_1 = rnode_5to168_bb1_idxprom_0_stall_out_reg_168_NO_SHIFT_REG;
assign rnode_5to168_bb1_idxprom_0_NO_SHIFT_REG = rnode_5to168_bb1_idxprom_0_reg_168_NO_SHIFT_REG;
assign rnode_5to168_bb1_idxprom_0_stall_in_reg_168_NO_SHIFT_REG = rnode_5to168_bb1_idxprom_0_stall_in_NO_SHIFT_REG;
assign rnode_5to168_bb1_idxprom_0_valid_out_NO_SHIFT_REG = rnode_5to168_bb1_idxprom_0_valid_out_reg_168_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb1_arrayidx_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb1_arrayidx_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_5to6_bb1_arrayidx_0_NO_SHIFT_REG;
 logic rnode_5to6_bb1_arrayidx_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_5to6_bb1_arrayidx_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb1_arrayidx_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb1_arrayidx_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb1_arrayidx_0_stall_out_reg_6_NO_SHIFT_REG;
wire [159:0] rci_rcnode_168to169_rc0_input_global_id_1_0_reg_168;

acl_data_fifo rnode_5to6_bb1_arrayidx_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb1_arrayidx_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb1_arrayidx_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb1_arrayidx_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb1_arrayidx_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in((local_bb1_arrayidx & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_5to6_bb1_arrayidx_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb1_arrayidx_0_reg_6_fifo.DEPTH = 2;
defparam rnode_5to6_bb1_arrayidx_0_reg_6_fifo.DATA_WIDTH = 64;
defparam rnode_5to6_bb1_arrayidx_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_5to6_bb1_arrayidx_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_5to6_bb1_arrayidx_0_reg_6_inputs_ready_NO_SHIFT_REG = local_bb1_arrayidx_valid_out;
assign local_bb1_arrayidx_stall_in = rnode_5to6_bb1_arrayidx_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb1_arrayidx_0_NO_SHIFT_REG = rnode_5to6_bb1_arrayidx_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb1_arrayidx_0_stall_in_reg_6_NO_SHIFT_REG = rnode_5to6_bb1_arrayidx_0_stall_in_NO_SHIFT_REG;
assign rnode_5to6_bb1_arrayidx_0_valid_out_NO_SHIFT_REG = rnode_5to6_bb1_arrayidx_0_valid_out_reg_6_NO_SHIFT_REG;
assign rci_rcnode_168to169_rc0_input_global_id_1_0_reg_168[31:0] = rcnode_1to168_rc2_input_global_id_1_0_NO_SHIFT_REG[31:0];
assign rci_rcnode_168to169_rc0_input_global_id_1_0_reg_168[63:32] = rcnode_1to168_rc2_input_global_id_1_0_NO_SHIFT_REG[63:32];
assign rci_rcnode_168to169_rc0_input_global_id_1_0_reg_168[95:64] = rnode_4to168_input_global_id_0_0_NO_SHIFT_REG;
assign rci_rcnode_168to169_rc0_input_global_id_1_0_reg_168[159:96] = (rnode_5to168_bb1_idxprom_0_NO_SHIFT_REG & 64'hFFFFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_168to169_rc0_input_global_id_1_0_valid_out_NO_SHIFT_REG;
 logic rcnode_168to169_rc0_input_global_id_1_0_stall_in_NO_SHIFT_REG;
 logic [159:0] rcnode_168to169_rc0_input_global_id_1_0_NO_SHIFT_REG;
 logic rcnode_168to169_rc0_input_global_id_1_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [159:0] rcnode_168to169_rc0_input_global_id_1_0_reg_169_NO_SHIFT_REG;
 logic rcnode_168to169_rc0_input_global_id_1_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rcnode_168to169_rc0_input_global_id_1_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_IP_NO_SHIFT_REG;
 logic rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_NO_SHIFT_REG;

acl_data_fifo rcnode_168to169_rc0_input_global_id_1_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_168to169_rc0_input_global_id_1_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_168to169_rc0_input_global_id_1_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rcnode_168to169_rc0_input_global_id_1_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_168to169_rc0_input_global_id_1_0_reg_168),
	.data_out(rcnode_168to169_rc0_input_global_id_1_0_reg_169_NO_SHIFT_REG)
);

defparam rcnode_168to169_rc0_input_global_id_1_0_reg_169_fifo.DEPTH = 1;
defparam rcnode_168to169_rc0_input_global_id_1_0_reg_169_fifo.DATA_WIDTH = 160;
defparam rcnode_168to169_rc0_input_global_id_1_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_168to169_rc0_input_global_id_1_0_reg_169_fifo.IMPL = "ll_reg";

assign rcnode_168to169_rc0_input_global_id_1_0_reg_169_inputs_ready_NO_SHIFT_REG = (rnode_4to168_input_global_id_0_0_valid_out_NO_SHIFT_REG & rnode_5to168_bb1_idxprom_0_valid_out_NO_SHIFT_REG & rcnode_1to168_rc2_input_global_id_1_0_valid_out_NO_SHIFT_REG);
assign rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_NO_SHIFT_REG = (~(rcnode_168to169_rc0_input_global_id_1_0_reg_169_inputs_ready_NO_SHIFT_REG) | rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_IP_NO_SHIFT_REG);
assign rnode_4to168_input_global_id_0_0_stall_in_NO_SHIFT_REG = rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_NO_SHIFT_REG;
assign rnode_5to168_bb1_idxprom_0_stall_in_NO_SHIFT_REG = rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_NO_SHIFT_REG;
assign rcnode_1to168_rc2_input_global_id_1_0_stall_in_NO_SHIFT_REG = rcnode_168to169_rc0_input_global_id_1_0_stall_out_0_reg_169_NO_SHIFT_REG;
assign rcnode_168to169_rc0_input_global_id_1_0_NO_SHIFT_REG = rcnode_168to169_rc0_input_global_id_1_0_reg_169_NO_SHIFT_REG;
assign rcnode_168to169_rc0_input_global_id_1_0_stall_in_reg_169_NO_SHIFT_REG = rcnode_168to169_rc0_input_global_id_1_0_stall_in_NO_SHIFT_REG;
assign rcnode_168to169_rc0_input_global_id_1_0_valid_out_NO_SHIFT_REG = rcnode_168to169_rc0_input_global_id_1_0_valid_out_reg_169_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb1_ld__inputs_ready;
 reg local_bb1_ld__valid_out_NO_SHIFT_REG;
wire local_bb1_ld__stall_in;
wire local_bb1_ld__output_regs_ready;
wire local_bb1_ld__fu_stall_out;
wire local_bb1_ld__fu_valid_out;
wire [31:0] local_bb1_ld__lsu_dataout;
 reg [31:0] local_bb1_ld__NO_SHIFT_REG;
wire local_bb1_ld__causedstall;

lsu_top lsu_local_bb1_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb1_ld__fu_stall_out),
	.i_valid(local_bb1_ld__inputs_ready),
	.i_address((rnode_5to6_bb1_arrayidx_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(1'b0),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb1_ld__output_regs_ready)),
	.o_valid(local_bb1_ld__fu_valid_out),
	.o_readdata(local_bb1_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb1_ld__active),
	.avm_address(avm_local_bb1_ld__address),
	.avm_read(avm_local_bb1_ld__read),
	.avm_readdata(avm_local_bb1_ld__readdata),
	.avm_write(avm_local_bb1_ld__write),
	.avm_writeack(avm_local_bb1_ld__writeack),
	.avm_burstcount(avm_local_bb1_ld__burstcount),
	.avm_writedata(avm_local_bb1_ld__writedata),
	.avm_byteenable(avm_local_bb1_ld__byteenable),
	.avm_waitrequest(avm_local_bb1_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb1_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb1_ld_.AWIDTH = 33;
defparam lsu_local_bb1_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb1_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb1_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb1_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb1_ld_.READ = 1;
defparam lsu_local_bb1_ld_.ATOMIC = 0;
defparam lsu_local_bb1_ld_.WIDTH = 32;
defparam lsu_local_bb1_ld_.MWIDTH = 512;
defparam lsu_local_bb1_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb1_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb1_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb1_ld_.MEMORY_SIDE_MEM_LATENCY = 132;
defparam lsu_local_bb1_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb1_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb1_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb1_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb1_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb1_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb1_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb1_ld_.USECACHING = 0;
defparam lsu_local_bb1_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb1_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb1_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb1_ld_.ADDRSPACE = 1;
defparam lsu_local_bb1_ld_.STYLE = "BURST-COALESCED";

assign local_bb1_ld__inputs_ready = rnode_5to6_bb1_arrayidx_0_valid_out_NO_SHIFT_REG;
assign local_bb1_ld__output_regs_ready = (&(~(local_bb1_ld__valid_out_NO_SHIFT_REG) | ~(local_bb1_ld__stall_in)));
assign rnode_5to6_bb1_arrayidx_0_stall_in_NO_SHIFT_REG = (local_bb1_ld__fu_stall_out | ~(local_bb1_ld__inputs_ready));
assign local_bb1_ld__causedstall = (local_bb1_ld__inputs_ready && (local_bb1_ld__fu_stall_out && !(~(local_bb1_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_ld__NO_SHIFT_REG <= 'x;
		local_bb1_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_ld__output_regs_ready)
		begin
			local_bb1_ld__NO_SHIFT_REG <= local_bb1_ld__lsu_dataout;
			local_bb1_ld__valid_out_NO_SHIFT_REG <= local_bb1_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb1_ld__stall_in))
			begin
				local_bb1_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_166to166_bb1_ld__valid_out_0;
wire rstag_166to166_bb1_ld__stall_in_0;
wire rstag_166to166_bb1_ld__valid_out_1;
wire rstag_166to166_bb1_ld__stall_in_1;
wire rstag_166to166_bb1_ld__inputs_ready;
wire rstag_166to166_bb1_ld__stall_local;
 reg rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG;
wire rstag_166to166_bb1_ld__combined_valid;
 reg [31:0] rstag_166to166_bb1_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_166to166_bb1_ld_;
 reg rstag_166to166_bb1_ld__consumed_0_NO_SHIFT_REG;
 reg rstag_166to166_bb1_ld__consumed_1_NO_SHIFT_REG;

assign rstag_166to166_bb1_ld__inputs_ready = local_bb1_ld__valid_out_NO_SHIFT_REG;
assign rstag_166to166_bb1_ld_ = (rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG ? rstag_166to166_bb1_ld__staging_reg_NO_SHIFT_REG : local_bb1_ld__NO_SHIFT_REG);
assign rstag_166to166_bb1_ld__combined_valid = (rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG | rstag_166to166_bb1_ld__inputs_ready);
assign rstag_166to166_bb1_ld__stall_local = ((rstag_166to166_bb1_ld__stall_in_0 & ~(rstag_166to166_bb1_ld__consumed_0_NO_SHIFT_REG)) | (rstag_166to166_bb1_ld__stall_in_1 & ~(rstag_166to166_bb1_ld__consumed_1_NO_SHIFT_REG)));
assign rstag_166to166_bb1_ld__valid_out_0 = (rstag_166to166_bb1_ld__combined_valid & ~(rstag_166to166_bb1_ld__consumed_0_NO_SHIFT_REG));
assign rstag_166to166_bb1_ld__valid_out_1 = (rstag_166to166_bb1_ld__combined_valid & ~(rstag_166to166_bb1_ld__consumed_1_NO_SHIFT_REG));
assign local_bb1_ld__stall_in = (|rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_166to166_bb1_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_166to166_bb1_ld__stall_local)
		begin
			if (~(rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG <= rstag_166to166_bb1_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_166to166_bb1_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_166to166_bb1_ld__staging_reg_NO_SHIFT_REG <= local_bb1_ld__NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_166to166_bb1_ld__consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_166to166_bb1_ld__consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_166to166_bb1_ld__consumed_0_NO_SHIFT_REG <= (rstag_166to166_bb1_ld__combined_valid & (rstag_166to166_bb1_ld__consumed_0_NO_SHIFT_REG | ~(rstag_166to166_bb1_ld__stall_in_0)) & rstag_166to166_bb1_ld__stall_local);
		rstag_166to166_bb1_ld__consumed_1_NO_SHIFT_REG <= (rstag_166to166_bb1_ld__combined_valid & (rstag_166to166_bb1_ld__consumed_1_NO_SHIFT_REG | ~(rstag_166to166_bb1_ld__stall_in_1)) & rstag_166to166_bb1_ld__stall_local);
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_166to169_bb1_ld__0_valid_out_NO_SHIFT_REG;
 logic rnode_166to169_bb1_ld__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to169_bb1_ld__0_NO_SHIFT_REG;
 logic rnode_166to169_bb1_ld__0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to169_bb1_ld__0_reg_169_NO_SHIFT_REG;
 logic rnode_166to169_bb1_ld__0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_166to169_bb1_ld__0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_166to169_bb1_ld__0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_166to169_bb1_ld__0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to169_bb1_ld__0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to169_bb1_ld__0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_166to169_bb1_ld__0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_166to169_bb1_ld__0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rstag_166to166_bb1_ld_),
	.data_out(rnode_166to169_bb1_ld__0_reg_169_NO_SHIFT_REG)
);

defparam rnode_166to169_bb1_ld__0_reg_169_fifo.DEPTH = 4;
defparam rnode_166to169_bb1_ld__0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_166to169_bb1_ld__0_reg_169_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_166to169_bb1_ld__0_reg_169_fifo.IMPL = "ll_reg";

assign rnode_166to169_bb1_ld__0_reg_169_inputs_ready_NO_SHIFT_REG = rstag_166to166_bb1_ld__valid_out_0;
assign rstag_166to166_bb1_ld__stall_in_0 = rnode_166to169_bb1_ld__0_stall_out_reg_169_NO_SHIFT_REG;
assign rnode_166to169_bb1_ld__0_NO_SHIFT_REG = rnode_166to169_bb1_ld__0_reg_169_NO_SHIFT_REG;
assign rnode_166to169_bb1_ld__0_stall_in_reg_169_NO_SHIFT_REG = rnode_166to169_bb1_ld__0_stall_in_NO_SHIFT_REG;
assign rnode_166to169_bb1_ld__0_valid_out_NO_SHIFT_REG = rnode_166to169_bb1_ld__0_valid_out_reg_169_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb1_cmp_inputs_ready;
 reg local_bb1_cmp_valid_out_NO_SHIFT_REG;
wire local_bb1_cmp_stall_in;
wire local_bb1_cmp_output_regs_ready;
wire local_bb1_cmp;
 reg local_bb1_cmp_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb1_cmp_valid_pipe_1_NO_SHIFT_REG;
wire local_bb1_cmp_causedstall;

acl_fp_cmp fp_module_local_bb1_cmp (
	.clock(clock),
	.dataa(rstag_166to166_bb1_ld_),
	.datab(32'h0),
	.enable(local_bb1_cmp_output_regs_ready),
	.result(local_bb1_cmp)
);

defparam fp_module_local_bb1_cmp.COMPARISON_MODE = 0;

assign local_bb1_cmp_inputs_ready = rstag_166to166_bb1_ld__valid_out_1;
assign local_bb1_cmp_output_regs_ready = (&(~(local_bb1_cmp_valid_out_NO_SHIFT_REG) | ~(local_bb1_cmp_stall_in)));
assign rstag_166to166_bb1_ld__stall_in_1 = (~(local_bb1_cmp_output_regs_ready) | ~(local_bb1_cmp_inputs_ready));
assign local_bb1_cmp_causedstall = (local_bb1_cmp_inputs_ready && (~(local_bb1_cmp_output_regs_ready) && !(~(local_bb1_cmp_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_cmp_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb1_cmp_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_cmp_output_regs_ready)
		begin
			local_bb1_cmp_valid_pipe_0_NO_SHIFT_REG <= local_bb1_cmp_inputs_ready;
			local_bb1_cmp_valid_pipe_1_NO_SHIFT_REG <= local_bb1_cmp_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_cmp_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_cmp_output_regs_ready)
		begin
			local_bb1_cmp_valid_out_NO_SHIFT_REG <= local_bb1_cmp_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb1_cmp_stall_in))
			begin
				local_bb1_cmp_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_169to169_bb1_cmp_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_1_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_reg_169_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_169to169_bb1_cmp_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_169to169_bb1_cmp_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to169_bb1_cmp_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to169_bb1_cmp_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_169to169_bb1_cmp_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_169to169_bb1_cmp_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(local_bb1_cmp),
	.data_out(rnode_169to169_bb1_cmp_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_169to169_bb1_cmp_0_reg_169_fifo.DEPTH = 3;
defparam rnode_169to169_bb1_cmp_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_169to169_bb1_cmp_0_reg_169_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_169to169_bb1_cmp_0_reg_169_fifo.IMPL = "zl_reg";

assign rnode_169to169_bb1_cmp_0_reg_169_inputs_ready_NO_SHIFT_REG = local_bb1_cmp_valid_out_NO_SHIFT_REG;
assign local_bb1_cmp_stall_in = rnode_169to169_bb1_cmp_0_stall_out_reg_169_NO_SHIFT_REG;
assign rnode_169to169_bb1_cmp_0_stall_in_0_reg_169_NO_SHIFT_REG = (rnode_169to169_bb1_cmp_0_stall_in_0_NO_SHIFT_REG | rnode_169to169_bb1_cmp_0_stall_in_1_NO_SHIFT_REG);
assign rnode_169to169_bb1_cmp_0_valid_out_0_NO_SHIFT_REG = rnode_169to169_bb1_cmp_0_valid_out_0_reg_169_NO_SHIFT_REG;
assign rnode_169to169_bb1_cmp_0_valid_out_1_NO_SHIFT_REG = rnode_169to169_bb1_cmp_0_valid_out_0_reg_169_NO_SHIFT_REG;
assign rnode_169to169_bb1_cmp_0_NO_SHIFT_REG = rnode_169to169_bb1_cmp_0_reg_169_NO_SHIFT_REG;
assign rnode_169to169_bb1_cmp_1_NO_SHIFT_REG = rnode_169to169_bb1_cmp_0_reg_169_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb1_var__valid_out;
wire local_bb1_var__stall_in;
wire local_bb1_var__inputs_ready;
wire local_bb1_var__stall_local;
wire local_bb1_var_;

assign local_bb1_var__inputs_ready = rnode_169to169_bb1_cmp_0_valid_out_1_NO_SHIFT_REG;
assign local_bb1_var_ = (rnode_169to169_bb1_cmp_1_NO_SHIFT_REG | input_wii_cmp1622);
assign local_bb1_var__valid_out = local_bb1_var__inputs_ready;
assign local_bb1_var__stall_local = local_bb1_var__stall_in;
assign rnode_169to169_bb1_cmp_0_stall_in_1_NO_SHIFT_REG = (|local_bb1_var__stall_local);

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_bb1_idxprom_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb1_ld__reg_NO_SHIFT_REG;
 reg lvb_bb1_cmp_reg_NO_SHIFT_REG;
 reg lvb_bb1_var__reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb1_var__valid_out & rnode_166to169_bb1_ld__0_valid_out_NO_SHIFT_REG & rnode_169to169_bb1_cmp_0_valid_out_0_NO_SHIFT_REG & rcnode_168to169_rc0_input_global_id_1_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb1_var__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_166to169_bb1_ld__0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_169to169_bb1_cmp_0_stall_in_0_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_168to169_rc0_input_global_id_1_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb1_idxprom = lvb_bb1_idxprom_reg_NO_SHIFT_REG;
assign lvb_bb1_ld_ = lvb_bb1_ld__reg_NO_SHIFT_REG;
assign lvb_bb1_cmp = lvb_bb1_cmp_reg_NO_SHIFT_REG;
assign lvb_bb1_var_ = lvb_bb1_var__reg_NO_SHIFT_REG;
assign lvb_input_global_id_0 = lvb_input_global_id_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1 = lvb_input_global_id_1_reg_NO_SHIFT_REG;
assign lvb_input_acl_hw_wg_id = lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb1_idxprom_reg_NO_SHIFT_REG <= 'x;
		lvb_bb1_ld__reg_NO_SHIFT_REG <= 'x;
		lvb_bb1_cmp_reg_NO_SHIFT_REG <= 'x;
		lvb_bb1_var__reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_reg_NO_SHIFT_REG <= 'x;
		lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb1_idxprom_reg_NO_SHIFT_REG <= (rcnode_168to169_rc0_input_global_id_1_0_NO_SHIFT_REG[159:96] & 64'hFFFFFFFF);
			lvb_bb1_ld__reg_NO_SHIFT_REG <= rnode_166to169_bb1_ld__0_NO_SHIFT_REG;
			lvb_bb1_cmp_reg_NO_SHIFT_REG <= rnode_169to169_bb1_cmp_0_NO_SHIFT_REG;
			lvb_bb1_var__reg_NO_SHIFT_REG <= local_bb1_var_;
			lvb_input_global_id_0_reg_NO_SHIFT_REG <= rcnode_168to169_rc0_input_global_id_1_0_NO_SHIFT_REG[95:64];
			lvb_input_global_id_1_reg_NO_SHIFT_REG <= rcnode_168to169_rc0_input_global_id_1_0_NO_SHIFT_REG[31:0];
			lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG <= rcnode_168to169_rc0_input_global_id_1_0_NO_SHIFT_REG[63:32];
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_2
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_gaussian,
		input [31:0] 		input_wii_sub25,
		input [31:0] 		input_wii_sub29,
		input [31:0] 		input_wii_mul50,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u4,
		input 		valid_in_0,
		output 		stall_out_0,
		input [63:0] 		input_idxprom_0,
		input [31:0] 		input_ld__0,
		input 		input_cmp_0,
		input 		input_var__u5_0,
		input [63:0] 		input_indvars_iv29_0,
		input [31:0] 		input_t_024_0,
		input [31:0] 		input_sum_023_0,
		input [31:0] 		input_global_id_0_0,
		input [31:0] 		input_global_id_1_0,
		input [31:0] 		input_acl_hw_wg_id_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [63:0] 		input_idxprom_1,
		input [31:0] 		input_ld__1,
		input 		input_cmp_1,
		input 		input_var__u5_1,
		input [63:0] 		input_indvars_iv29_1,
		input [31:0] 		input_t_024_1,
		input [31:0] 		input_sum_023_1,
		input [31:0] 		input_global_id_0_1,
		input [31:0] 		input_global_id_1_1,
		input [31:0] 		input_acl_hw_wg_id_1,
		output 		valid_out,
		input 		stall_in,
		output [63:0] 		lvb_idxprom,
		output [31:0] 		lvb_ld_,
		output 		lvb_cmp,
		output 		lvb_var__u5,
		output [63:0] 		lvb_indvars_iv29,
		output [31:0] 		lvb_t_024,
		output [31:0] 		lvb_sum_023,
		output [31:0] 		lvb_bb2_sub25_add24,
		output [63:0] 		lvb_bb2_arrayidx43,
		output [31:0] 		lvb_input_global_id_0,
		output [31:0] 		lvb_input_global_id_1,
		output [31:0] 		lvb_input_acl_hw_wg_id,
		input [31:0] 		workgroup_size,
		input 		start
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_idxprom_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_ld__0_staging_reg_NO_SHIFT_REG;
 reg input_cmp_0_staging_reg_NO_SHIFT_REG;
 reg input_var__u5_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv29_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_024_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_023_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_idxprom_NO_SHIFT_REG;
 reg [31:0] local_lvm_ld__NO_SHIFT_REG;
 reg local_lvm_cmp_NO_SHIFT_REG;
 reg local_lvm_var__u5_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv29_NO_SHIFT_REG;
 reg [31:0] local_lvm_t_024_NO_SHIFT_REG;
 reg [31:0] local_lvm_sum_023_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_idxprom_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_ld__1_staging_reg_NO_SHIFT_REG;
 reg input_cmp_1_staging_reg_NO_SHIFT_REG;
 reg input_var__u5_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv29_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_024_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_023_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_idxprom_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_ld__0_staging_reg_NO_SHIFT_REG <= 'x;
		input_cmp_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u5_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv29_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_t_024_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_023_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_idxprom_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_ld__1_staging_reg_NO_SHIFT_REG <= 'x;
		input_cmp_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u5_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv29_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_t_024_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_023_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_idxprom_0_staging_reg_NO_SHIFT_REG <= input_idxprom_0;
				input_ld__0_staging_reg_NO_SHIFT_REG <= input_ld__0;
				input_cmp_0_staging_reg_NO_SHIFT_REG <= input_cmp_0;
				input_var__u5_0_staging_reg_NO_SHIFT_REG <= input_var__u5_0;
				input_indvars_iv29_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv29_0;
				input_t_024_0_staging_reg_NO_SHIFT_REG <= input_t_024_0;
				input_sum_023_0_staging_reg_NO_SHIFT_REG <= input_sum_023_0;
				input_global_id_0_0_staging_reg_NO_SHIFT_REG <= input_global_id_0_0;
				input_global_id_1_0_staging_reg_NO_SHIFT_REG <= input_global_id_1_0;
				input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_idxprom_1_staging_reg_NO_SHIFT_REG <= input_idxprom_1;
				input_ld__1_staging_reg_NO_SHIFT_REG <= input_ld__1;
				input_cmp_1_staging_reg_NO_SHIFT_REG <= input_cmp_1;
				input_var__u5_1_staging_reg_NO_SHIFT_REG <= input_var__u5_1;
				input_indvars_iv29_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv29_1;
				input_t_024_1_staging_reg_NO_SHIFT_REG <= input_t_024_1;
				input_sum_023_1_staging_reg_NO_SHIFT_REG <= input_sum_023_1;
				input_global_id_0_1_staging_reg_NO_SHIFT_REG <= input_global_id_0_1;
				input_global_id_1_1_staging_reg_NO_SHIFT_REG <= input_global_id_1_1;
				input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_0_staging_reg_NO_SHIFT_REG;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__0_staging_reg_NO_SHIFT_REG;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u5_NO_SHIFT_REG <= input_var__u5_0_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_0_staging_reg_NO_SHIFT_REG;
					local_lvm_t_024_NO_SHIFT_REG <= input_t_024_0_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_023_NO_SHIFT_REG <= input_sum_023_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_0;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__0;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_0;
					local_lvm_var__u5_NO_SHIFT_REG <= input_var__u5_0;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_0;
					local_lvm_t_024_NO_SHIFT_REG <= input_t_024_0;
					local_lvm_sum_023_NO_SHIFT_REG <= input_sum_023_0;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_0;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_1_staging_reg_NO_SHIFT_REG;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__1_staging_reg_NO_SHIFT_REG;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u5_NO_SHIFT_REG <= input_var__u5_1_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_1_staging_reg_NO_SHIFT_REG;
					local_lvm_t_024_NO_SHIFT_REG <= input_t_024_1_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_023_NO_SHIFT_REG <= input_sum_023_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_1;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__1;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_1;
					local_lvm_var__u5_NO_SHIFT_REG <= input_var__u5_1;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_1;
					local_lvm_t_024_NO_SHIFT_REG <= input_t_024_1;
					local_lvm_sum_023_NO_SHIFT_REG <= input_sum_023_1;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_1;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_1;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__stall_local;
wire [31:0] local_bb2_var_;

assign local_bb2_var_ = local_lvm_indvars_iv29_NO_SHIFT_REG[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u6_valid_out;
wire local_bb2_var__u6_stall_in;
wire local_bb2_var__u6_inputs_ready;
wire local_bb2_var__u6_stall_local;
wire [63:0] local_bb2_var__u6;
wire [321:0] rci_rcnode_1to3_rc3_idxprom_0_reg_1;

assign local_bb2_var__u6_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign local_bb2_var__u6 = (local_lvm_indvars_iv29_NO_SHIFT_REG + input_wii_var__u4);
assign local_bb2_var__u6_valid_out = local_bb2_var__u6_inputs_ready;
assign local_bb2_var__u6_stall_local = local_bb2_var__u6_stall_in;
assign merge_node_stall_in_2 = (|local_bb2_var__u6_stall_local);
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[63:0] = (local_lvm_idxprom_NO_SHIFT_REG & 64'hFFFFFFFF);
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[95:64] = local_lvm_ld__NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[96] = local_lvm_cmp_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[97] = local_lvm_var__u5_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[161:98] = local_lvm_indvars_iv29_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[193:162] = local_lvm_t_024_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[225:194] = local_lvm_sum_023_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[257:226] = local_lvm_input_global_id_0_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[289:258] = local_lvm_input_global_id_1_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc3_idxprom_0_reg_1[321:290] = local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rcnode_1to3_rc3_idxprom_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to3_rc3_idxprom_0_stall_in_NO_SHIFT_REG;
 logic [321:0] rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG;
 logic rcnode_1to3_rc3_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [321:0] rcnode_1to3_rc3_idxprom_0_reg_3_NO_SHIFT_REG;
 logic rcnode_1to3_rc3_idxprom_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rcnode_1to3_rc3_idxprom_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rcnode_1to3_rc3_idxprom_0_stall_out_reg_3_IP_NO_SHIFT_REG;
 logic rcnode_1to3_rc3_idxprom_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rcnode_1to3_rc3_idxprom_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to3_rc3_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to3_rc3_idxprom_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rcnode_1to3_rc3_idxprom_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rcnode_1to3_rc3_idxprom_0_stall_out_reg_3_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to3_rc3_idxprom_0_reg_1),
	.data_out(rcnode_1to3_rc3_idxprom_0_reg_3_NO_SHIFT_REG)
);

defparam rcnode_1to3_rc3_idxprom_0_reg_3_fifo.DEPTH = 3;
defparam rcnode_1to3_rc3_idxprom_0_reg_3_fifo.DATA_WIDTH = 322;
defparam rcnode_1to3_rc3_idxprom_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to3_rc3_idxprom_0_reg_3_fifo.IMPL = "ll_reg";

assign rcnode_1to3_rc3_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_3_NO_SHIFT_REG;
assign rcnode_1to3_rc3_idxprom_0_stall_out_reg_3_NO_SHIFT_REG = (~(rcnode_1to3_rc3_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG) | rcnode_1to3_rc3_idxprom_0_stall_out_reg_3_IP_NO_SHIFT_REG);
assign merge_node_stall_in_3 = rcnode_1to3_rc3_idxprom_0_stall_out_reg_3_NO_SHIFT_REG;
assign rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG = rcnode_1to3_rc3_idxprom_0_reg_3_NO_SHIFT_REG;
assign rcnode_1to3_rc3_idxprom_0_stall_in_reg_3_NO_SHIFT_REG = rcnode_1to3_rc3_idxprom_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to3_rc3_idxprom_0_valid_out_NO_SHIFT_REG = rcnode_1to3_rc3_idxprom_0_valid_out_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_add24_valid_out;
wire local_bb2_add24_stall_in;
wire local_bb2_add24_inputs_ready;
wire local_bb2_add24_stall_local;
wire [31:0] local_bb2_add24;

assign local_bb2_add24_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign local_bb2_add24 = (local_bb2_var_ + local_lvm_input_global_id_0_NO_SHIFT_REG);
assign local_bb2_add24_valid_out = local_bb2_add24_inputs_ready;
assign local_bb2_add24_stall_local = local_bb2_add24_stall_in;
assign merge_node_stall_in_0 = (local_bb2_add24_stall_local | ~(local_bb2_add24_inputs_ready));
assign merge_node_stall_in_1 = (local_bb2_add24_stall_local | ~(local_bb2_add24_inputs_ready));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb2_var__u6_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u6_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb2_var__u6_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u6_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb2_var__u6_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u6_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u6_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u6_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb2_var__u6_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb2_var__u6_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb2_var__u6_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb2_var__u6_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb2_var__u6_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb2_var__u6),
	.data_out(rnode_1to2_bb2_var__u6_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb2_var__u6_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb2_var__u6_0_reg_2_fifo.DATA_WIDTH = 64;
defparam rnode_1to2_bb2_var__u6_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb2_var__u6_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb2_var__u6_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb2_var__u6_valid_out;
assign local_bb2_var__u6_stall_in = rnode_1to2_bb2_var__u6_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u6_0_NO_SHIFT_REG = rnode_1to2_bb2_var__u6_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u6_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb2_var__u6_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u6_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb2_var__u6_0_valid_out_reg_2_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb2_add24_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add24_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_add24_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add24_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add24_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_add24_1_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add24_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_add24_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add24_0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add24_0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add24_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb2_add24_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb2_add24_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb2_add24_0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb2_add24_0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb2_add24_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb2_add24),
	.data_out(rnode_1to2_bb2_add24_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb2_add24_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb2_add24_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb2_add24_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb2_add24_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb2_add24_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb2_add24_valid_out;
assign local_bb2_add24_stall_in = rnode_1to2_bb2_add24_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_add24_0_stall_in_0_reg_2_NO_SHIFT_REG = (rnode_1to2_bb2_add24_0_stall_in_0_NO_SHIFT_REG | rnode_1to2_bb2_add24_0_stall_in_1_NO_SHIFT_REG);
assign rnode_1to2_bb2_add24_0_valid_out_0_NO_SHIFT_REG = rnode_1to2_bb2_add24_0_valid_out_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_add24_0_valid_out_1_NO_SHIFT_REG = rnode_1to2_bb2_add24_0_valid_out_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_add24_0_NO_SHIFT_REG = rnode_1to2_bb2_add24_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_add24_1_NO_SHIFT_REG = rnode_1to2_bb2_add24_0_reg_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx43_valid_out;
wire local_bb2_arrayidx43_stall_in;
wire local_bb2_arrayidx43_inputs_ready;
wire local_bb2_arrayidx43_stall_local;
wire [63:0] local_bb2_arrayidx43;

assign local_bb2_arrayidx43_inputs_ready = rnode_1to2_bb2_var__u6_0_valid_out_NO_SHIFT_REG;
assign local_bb2_arrayidx43 = ((input_gaussian & 64'hFFFFFFFFFFFFFC00) + (rnode_1to2_bb2_var__u6_0_NO_SHIFT_REG << 6'h2));
assign local_bb2_arrayidx43_valid_out = local_bb2_arrayidx43_inputs_ready;
assign local_bb2_arrayidx43_stall_local = local_bb2_arrayidx43_stall_in;
assign rnode_1to2_bb2_var__u6_0_stall_in_NO_SHIFT_REG = (|local_bb2_arrayidx43_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp1_i_valid_out;
wire local_bb2_cmp1_i_stall_in;
wire local_bb2_cmp1_i_inputs_ready;
wire local_bb2_cmp1_i_stall_local;
wire local_bb2_cmp1_i;

assign local_bb2_cmp1_i_inputs_ready = rnode_1to2_bb2_add24_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_cmp1_i = (rnode_1to2_bb2_add24_0_NO_SHIFT_REG > input_wii_sub25);
assign local_bb2_cmp1_i_valid_out = local_bb2_cmp1_i_inputs_ready;
assign local_bb2_cmp1_i_stall_local = local_bb2_cmp1_i_stall_in;
assign rnode_1to2_bb2_add24_0_stall_in_0_NO_SHIFT_REG = (|local_bb2_cmp1_i_stall_local);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb2_arrayidx43_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx43_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb2_arrayidx43_0_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx43_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb2_arrayidx43_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx43_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx43_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx43_0_stall_out_reg_3_NO_SHIFT_REG;
wire [32:0] rci_rcnode_2to3_rc0_bb2_cmp1_i_0_reg_2;

acl_data_fifo rnode_2to3_bb2_arrayidx43_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb2_arrayidx43_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb2_arrayidx43_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb2_arrayidx43_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb2_arrayidx43_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in((local_bb2_arrayidx43 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_2to3_bb2_arrayidx43_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb2_arrayidx43_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb2_arrayidx43_0_reg_3_fifo.DATA_WIDTH = 64;
defparam rnode_2to3_bb2_arrayidx43_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb2_arrayidx43_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_2to3_bb2_arrayidx43_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb2_arrayidx43_valid_out;
assign local_bb2_arrayidx43_stall_in = rnode_2to3_bb2_arrayidx43_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx43_0_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx43_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx43_0_stall_in_reg_3_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx43_0_stall_in_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx43_0_valid_out_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx43_0_valid_out_reg_3_NO_SHIFT_REG;
assign rci_rcnode_2to3_rc0_bb2_cmp1_i_0_reg_2[0] = local_bb2_cmp1_i;
assign rci_rcnode_2to3_rc0_bb2_cmp1_i_0_reg_2[32:1] = rnode_1to2_bb2_add24_1_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_2to3_rc0_bb2_cmp1_i_0_valid_out_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb2_cmp1_i_0_stall_in_NO_SHIFT_REG;
 logic [32:0] rcnode_2to3_rc0_bb2_cmp1_i_0_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [32:0] rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb2_cmp1_i_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb2_cmp1_i_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb2_cmp1_i_0_stall_out_0_reg_3_IP_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb2_cmp1_i_0_stall_out_0_reg_3_NO_SHIFT_REG;

acl_data_fifo rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_2to3_rc0_bb2_cmp1_i_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rcnode_2to3_rc0_bb2_cmp1_i_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rcnode_2to3_rc0_bb2_cmp1_i_0_stall_out_0_reg_3_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_2to3_rc0_bb2_cmp1_i_0_reg_2),
	.data_out(rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_NO_SHIFT_REG)
);

defparam rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_fifo.DEPTH = 1;
defparam rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_fifo.DATA_WIDTH = 33;
defparam rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_fifo.IMPL = "ll_reg";

assign rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_inputs_ready_NO_SHIFT_REG = (local_bb2_cmp1_i_valid_out & rnode_1to2_bb2_add24_0_valid_out_1_NO_SHIFT_REG);
assign rcnode_2to3_rc0_bb2_cmp1_i_0_stall_out_0_reg_3_NO_SHIFT_REG = (~(rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_inputs_ready_NO_SHIFT_REG) | rcnode_2to3_rc0_bb2_cmp1_i_0_stall_out_0_reg_3_IP_NO_SHIFT_REG);
assign local_bb2_cmp1_i_stall_in = rcnode_2to3_rc0_bb2_cmp1_i_0_stall_out_0_reg_3_NO_SHIFT_REG;
assign rnode_1to2_bb2_add24_0_stall_in_1_NO_SHIFT_REG = rcnode_2to3_rc0_bb2_cmp1_i_0_stall_out_0_reg_3_NO_SHIFT_REG;
assign rcnode_2to3_rc0_bb2_cmp1_i_0_NO_SHIFT_REG = rcnode_2to3_rc0_bb2_cmp1_i_0_reg_3_NO_SHIFT_REG;
assign rcnode_2to3_rc0_bb2_cmp1_i_0_stall_in_reg_3_NO_SHIFT_REG = rcnode_2to3_rc0_bb2_cmp1_i_0_stall_in_NO_SHIFT_REG;
assign rcnode_2to3_rc0_bb2_cmp1_i_0_valid_out_NO_SHIFT_REG = rcnode_2to3_rc0_bb2_cmp1_i_0_valid_out_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_sub25_add24_valid_out;
wire local_bb2_sub25_add24_stall_in;
wire local_bb2_sub25_add24_inputs_ready;
wire local_bb2_sub25_add24_stall_local;
wire [31:0] local_bb2_sub25_add24;

assign local_bb2_sub25_add24_inputs_ready = rcnode_2to3_rc0_bb2_cmp1_i_0_valid_out_NO_SHIFT_REG;
assign local_bb2_sub25_add24 = (rcnode_2to3_rc0_bb2_cmp1_i_0_NO_SHIFT_REG[0] ? input_wii_sub25 : rcnode_2to3_rc0_bb2_cmp1_i_0_NO_SHIFT_REG[32:1]);
assign local_bb2_sub25_add24_valid_out = local_bb2_sub25_add24_inputs_ready;
assign local_bb2_sub25_add24_stall_local = local_bb2_sub25_add24_stall_in;
assign rcnode_2to3_rc0_bb2_cmp1_i_0_stall_in_NO_SHIFT_REG = (|local_bb2_sub25_add24_stall_local);

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_idxprom_reg_NO_SHIFT_REG;
 reg [31:0] lvb_ld__reg_NO_SHIFT_REG;
 reg lvb_cmp_reg_NO_SHIFT_REG;
 reg lvb_var__u5_reg_NO_SHIFT_REG;
 reg [63:0] lvb_indvars_iv29_reg_NO_SHIFT_REG;
 reg [31:0] lvb_t_024_reg_NO_SHIFT_REG;
 reg [31:0] lvb_sum_023_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb2_sub25_add24_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb2_arrayidx43_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb2_sub25_add24_valid_out & rnode_2to3_bb2_arrayidx43_0_valid_out_NO_SHIFT_REG & rcnode_1to3_rc3_idxprom_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb2_sub25_add24_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_2to3_bb2_arrayidx43_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_1to3_rc3_idxprom_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_idxprom = lvb_idxprom_reg_NO_SHIFT_REG;
assign lvb_ld_ = lvb_ld__reg_NO_SHIFT_REG;
assign lvb_cmp = lvb_cmp_reg_NO_SHIFT_REG;
assign lvb_var__u5 = lvb_var__u5_reg_NO_SHIFT_REG;
assign lvb_indvars_iv29 = lvb_indvars_iv29_reg_NO_SHIFT_REG;
assign lvb_t_024 = lvb_t_024_reg_NO_SHIFT_REG;
assign lvb_sum_023 = lvb_sum_023_reg_NO_SHIFT_REG;
assign lvb_bb2_sub25_add24 = lvb_bb2_sub25_add24_reg_NO_SHIFT_REG;
assign lvb_bb2_arrayidx43 = lvb_bb2_arrayidx43_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0 = lvb_input_global_id_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1 = lvb_input_global_id_1_reg_NO_SHIFT_REG;
assign lvb_input_acl_hw_wg_id = lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_idxprom_reg_NO_SHIFT_REG <= 'x;
		lvb_ld__reg_NO_SHIFT_REG <= 'x;
		lvb_cmp_reg_NO_SHIFT_REG <= 'x;
		lvb_var__u5_reg_NO_SHIFT_REG <= 'x;
		lvb_indvars_iv29_reg_NO_SHIFT_REG <= 'x;
		lvb_t_024_reg_NO_SHIFT_REG <= 'x;
		lvb_sum_023_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_sub25_add24_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_arrayidx43_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_reg_NO_SHIFT_REG <= 'x;
		lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_idxprom_reg_NO_SHIFT_REG <= (rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[63:0] & 64'hFFFFFFFF);
			lvb_ld__reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[95:64];
			lvb_cmp_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[96];
			lvb_var__u5_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[97];
			lvb_indvars_iv29_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[161:98];
			lvb_t_024_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[193:162];
			lvb_sum_023_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[225:194];
			lvb_bb2_sub25_add24_reg_NO_SHIFT_REG <= local_bb2_sub25_add24;
			lvb_bb2_arrayidx43_reg_NO_SHIFT_REG <= (rnode_2to3_bb2_arrayidx43_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
			lvb_input_global_id_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[257:226];
			lvb_input_global_id_1_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[289:258];
			lvb_input_acl_hw_wg_id_reg_NO_SHIFT_REG <= rcnode_1to3_rc3_idxprom_0_NO_SHIFT_REG[321:290];
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_3
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_gaussian,
		input [31:0] 		input_r,
		input [31:0] 		input_global_size_0,
		input [63:0] 		input_in,
		input [31:0] 		input_wii_sub25,
		input [31:0] 		input_wii_sub29,
		input [31:0] 		input_wii_mul50,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u7,
		input 		valid_in_0,
		output 		stall_out_0,
		input [63:0] 		input_idxprom_0,
		input [31:0] 		input_ld__0,
		input 		input_cmp_0,
		input 		input_var__u8_0,
		input [63:0] 		input_indvars_iv29_0,
		input [31:0] 		input_sub25_add24_0,
		input [63:0] 		input_arrayidx43_0,
		input [63:0] 		input_indvars_iv_0,
		input [31:0] 		input_t_119_0,
		input [31:0] 		input_sum_118_0,
		input [31:0] 		input_global_id_0_0,
		input [31:0] 		input_global_id_1_0,
		input [31:0] 		input_acl_hw_wg_id_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [63:0] 		input_idxprom_1,
		input [31:0] 		input_ld__1,
		input 		input_cmp_1,
		input 		input_var__u8_1,
		input [63:0] 		input_indvars_iv29_1,
		input [31:0] 		input_sub25_add24_1,
		input [63:0] 		input_arrayidx43_1,
		input [63:0] 		input_indvars_iv_1,
		input [31:0] 		input_t_119_1,
		input [31:0] 		input_sum_118_1,
		input [31:0] 		input_global_id_0_1,
		input [31:0] 		input_global_id_1_1,
		input [31:0] 		input_acl_hw_wg_id_1,
		output 		valid_out_0,
		input 		stall_in_0,
		output [63:0] 		lvb_idxprom_0,
		output [31:0] 		lvb_ld__0,
		output 		lvb_cmp_0,
		output 		lvb_var__u8_0,
		output [63:0] 		lvb_indvars_iv29_0,
		output [31:0] 		lvb_sub25_add24_0,
		output [63:0] 		lvb_arrayidx43_0,
		output [63:0] 		lvb_bb3_indvars_iv_next_0,
		output [31:0] 		lvb_bb3_c0_exe1_0,
		output [31:0] 		lvb_bb3_c0_exe2_0,
		output [31:0] 		lvb_input_global_id_0_0,
		output [31:0] 		lvb_input_global_id_1_0,
		output [31:0] 		lvb_input_acl_hw_wg_id_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [63:0] 		lvb_idxprom_1,
		output [31:0] 		lvb_ld__1,
		output 		lvb_cmp_1,
		output 		lvb_var__u8_1,
		output [63:0] 		lvb_indvars_iv29_1,
		output [31:0] 		lvb_sub25_add24_1,
		output [63:0] 		lvb_arrayidx43_1,
		output [63:0] 		lvb_bb3_indvars_iv_next_1,
		output [31:0] 		lvb_bb3_c0_exe1_1,
		output [31:0] 		lvb_bb3_c0_exe2_1,
		output [31:0] 		lvb_input_global_id_0_1,
		output [31:0] 		lvb_input_global_id_1_1,
		output [31:0] 		lvb_input_acl_hw_wg_id_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input [511:0] 		avm_local_bb3_ld__readdata,
		input 		avm_local_bb3_ld__readdatavalid,
		input 		avm_local_bb3_ld__waitrequest,
		output [32:0] 		avm_local_bb3_ld__address,
		output 		avm_local_bb3_ld__read,
		output 		avm_local_bb3_ld__write,
		input 		avm_local_bb3_ld__writeack,
		output [511:0] 		avm_local_bb3_ld__writedata,
		output [63:0] 		avm_local_bb3_ld__byteenable,
		output [4:0] 		avm_local_bb3_ld__burstcount,
		output 		local_bb3_ld__active,
		input 		clock2x,
		input [511:0] 		avm_local_bb3_ld__u12_readdata,
		input 		avm_local_bb3_ld__u12_readdatavalid,
		input 		avm_local_bb3_ld__u12_waitrequest,
		output [32:0] 		avm_local_bb3_ld__u12_address,
		output 		avm_local_bb3_ld__u12_read,
		output 		avm_local_bb3_ld__u12_write,
		input 		avm_local_bb3_ld__u12_writeack,
		output [511:0] 		avm_local_bb3_ld__u12_writedata,
		output [63:0] 		avm_local_bb3_ld__u12_byteenable,
		output [4:0] 		avm_local_bb3_ld__u12_burstcount,
		output 		local_bb3_ld__u12_active,
		input [511:0] 		avm_local_bb3_ld__u13_readdata,
		input 		avm_local_bb3_ld__u13_readdatavalid,
		input 		avm_local_bb3_ld__u13_waitrequest,
		output [32:0] 		avm_local_bb3_ld__u13_address,
		output 		avm_local_bb3_ld__u13_read,
		output 		avm_local_bb3_ld__u13_write,
		input 		avm_local_bb3_ld__u13_writeack,
		output [511:0] 		avm_local_bb3_ld__u13_writedata,
		output [63:0] 		avm_local_bb3_ld__u13_byteenable,
		output [4:0] 		avm_local_bb3_ld__u13_burstcount,
		output 		local_bb3_ld__u13_active
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_node_stall_in_8;
 reg merge_node_valid_out_8_NO_SHIFT_REG;
wire merge_node_stall_in_9;
 reg merge_node_valid_out_9_NO_SHIFT_REG;
wire merge_node_stall_in_10;
 reg merge_node_valid_out_10_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_idxprom_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_ld__0_staging_reg_NO_SHIFT_REG;
 reg input_cmp_0_staging_reg_NO_SHIFT_REG;
 reg input_var__u8_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv29_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sub25_add24_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_arrayidx43_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_119_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_118_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_idxprom_NO_SHIFT_REG;
 reg [31:0] local_lvm_ld__NO_SHIFT_REG;
 reg local_lvm_cmp_NO_SHIFT_REG;
 reg local_lvm_var__u8_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv29_NO_SHIFT_REG;
 reg [31:0] local_lvm_sub25_add24_NO_SHIFT_REG;
 reg [63:0] local_lvm_arrayidx43_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv_NO_SHIFT_REG;
 reg [31:0] local_lvm_t_119_NO_SHIFT_REG;
 reg [31:0] local_lvm_sum_118_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_idxprom_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_ld__1_staging_reg_NO_SHIFT_REG;
 reg input_cmp_1_staging_reg_NO_SHIFT_REG;
 reg input_var__u8_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv29_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sub25_add24_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_arrayidx43_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_119_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_118_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG) | (merge_node_stall_in_8 & merge_node_valid_out_8_NO_SHIFT_REG) | (merge_node_stall_in_9 & merge_node_valid_out_9_NO_SHIFT_REG) | (merge_node_stall_in_10 & merge_node_valid_out_10_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_idxprom_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_ld__0_staging_reg_NO_SHIFT_REG <= 'x;
		input_cmp_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u8_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv29_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_sub25_add24_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_arrayidx43_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_t_119_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_118_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_idxprom_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_ld__1_staging_reg_NO_SHIFT_REG <= 'x;
		input_cmp_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u8_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv29_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_sub25_add24_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_arrayidx43_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_t_119_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_118_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_idxprom_0_staging_reg_NO_SHIFT_REG <= input_idxprom_0;
				input_ld__0_staging_reg_NO_SHIFT_REG <= input_ld__0;
				input_cmp_0_staging_reg_NO_SHIFT_REG <= input_cmp_0;
				input_var__u8_0_staging_reg_NO_SHIFT_REG <= input_var__u8_0;
				input_indvars_iv29_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv29_0;
				input_sub25_add24_0_staging_reg_NO_SHIFT_REG <= input_sub25_add24_0;
				input_arrayidx43_0_staging_reg_NO_SHIFT_REG <= input_arrayidx43_0;
				input_indvars_iv_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv_0;
				input_t_119_0_staging_reg_NO_SHIFT_REG <= input_t_119_0;
				input_sum_118_0_staging_reg_NO_SHIFT_REG <= input_sum_118_0;
				input_global_id_0_0_staging_reg_NO_SHIFT_REG <= input_global_id_0_0;
				input_global_id_1_0_staging_reg_NO_SHIFT_REG <= input_global_id_1_0;
				input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_idxprom_1_staging_reg_NO_SHIFT_REG <= input_idxprom_1;
				input_ld__1_staging_reg_NO_SHIFT_REG <= input_ld__1;
				input_cmp_1_staging_reg_NO_SHIFT_REG <= input_cmp_1;
				input_var__u8_1_staging_reg_NO_SHIFT_REG <= input_var__u8_1;
				input_indvars_iv29_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv29_1;
				input_sub25_add24_1_staging_reg_NO_SHIFT_REG <= input_sub25_add24_1;
				input_arrayidx43_1_staging_reg_NO_SHIFT_REG <= input_arrayidx43_1;
				input_indvars_iv_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv_1;
				input_t_119_1_staging_reg_NO_SHIFT_REG <= input_t_119_1;
				input_sum_118_1_staging_reg_NO_SHIFT_REG <= input_sum_118_1;
				input_global_id_0_1_staging_reg_NO_SHIFT_REG <= input_global_id_0_1;
				input_global_id_1_1_staging_reg_NO_SHIFT_REG <= input_global_id_1_1;
				input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_0_staging_reg_NO_SHIFT_REG;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__0_staging_reg_NO_SHIFT_REG;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u8_NO_SHIFT_REG <= input_var__u8_0_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_0_staging_reg_NO_SHIFT_REG;
					local_lvm_sub25_add24_NO_SHIFT_REG <= input_sub25_add24_0_staging_reg_NO_SHIFT_REG;
					local_lvm_arrayidx43_NO_SHIFT_REG <= input_arrayidx43_0_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_0_staging_reg_NO_SHIFT_REG;
					local_lvm_t_119_NO_SHIFT_REG <= input_t_119_0_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_118_NO_SHIFT_REG <= input_sum_118_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_0;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__0;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_0;
					local_lvm_var__u8_NO_SHIFT_REG <= input_var__u8_0;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_0;
					local_lvm_sub25_add24_NO_SHIFT_REG <= input_sub25_add24_0;
					local_lvm_arrayidx43_NO_SHIFT_REG <= input_arrayidx43_0;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_0;
					local_lvm_t_119_NO_SHIFT_REG <= input_t_119_0;
					local_lvm_sum_118_NO_SHIFT_REG <= input_sum_118_0;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_0;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_1_staging_reg_NO_SHIFT_REG;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__1_staging_reg_NO_SHIFT_REG;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u8_NO_SHIFT_REG <= input_var__u8_1_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_1_staging_reg_NO_SHIFT_REG;
					local_lvm_sub25_add24_NO_SHIFT_REG <= input_sub25_add24_1_staging_reg_NO_SHIFT_REG;
					local_lvm_arrayidx43_NO_SHIFT_REG <= input_arrayidx43_1_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_1_staging_reg_NO_SHIFT_REG;
					local_lvm_t_119_NO_SHIFT_REG <= input_t_119_1_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_118_NO_SHIFT_REG <= input_sum_118_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_1;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__1;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_1;
					local_lvm_var__u8_NO_SHIFT_REG <= input_var__u8_1;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_1;
					local_lvm_sub25_add24_NO_SHIFT_REG <= input_sub25_add24_1;
					local_lvm_arrayidx43_NO_SHIFT_REG <= input_arrayidx43_1;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_1;
					local_lvm_t_119_NO_SHIFT_REG <= input_t_119_1;
					local_lvm_sum_118_NO_SHIFT_REG <= input_sum_118_1;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_1;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_1;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_9_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_10_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_8_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_9_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_10_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_8))
			begin
				merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_9))
			begin
				merge_node_valid_out_9_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_10))
			begin
				merge_node_valid_out_10_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_var__stall_local;
wire [31:0] local_bb3_var_;

assign local_bb3_var_ = local_lvm_indvars_iv_NO_SHIFT_REG[31:0];

// Register node:
//  * latency = 167
//  * capacity = 167
 logic rnode_1to168_var__u7_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to168_var__u7_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to168_var__u7_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to168_var__u7_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_1to168_var__u7_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_1to168_var__u7_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_1to168_var__u7_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to168_var__u7_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to168_var__u7_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_1to168_var__u7_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_1to168_var__u7_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to168_var__u7_0_reg_168_fifo.DEPTH = 168;
defparam rnode_1to168_var__u7_0_reg_168_fifo.DATA_WIDTH = 0;
defparam rnode_1to168_var__u7_0_reg_168_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to168_var__u7_0_reg_168_fifo.IMPL = "ram";

assign rnode_1to168_var__u7_0_reg_168_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign merge_node_stall_in_2 = rnode_1to168_var__u7_0_stall_out_reg_168_NO_SHIFT_REG;
assign rnode_1to168_var__u7_0_stall_in_reg_168_NO_SHIFT_REG = rnode_1to168_var__u7_0_stall_in_NO_SHIFT_REG;
assign rnode_1to168_var__u7_0_valid_out_NO_SHIFT_REG = rnode_1to168_var__u7_0_valid_out_reg_168_NO_SHIFT_REG;

// Register node:
//  * latency = 167
//  * capacity = 167
 logic rnode_1to168_indvars_iv_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to168_indvars_iv_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_1to168_indvars_iv_0_NO_SHIFT_REG;
 logic rnode_1to168_indvars_iv_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to168_indvars_iv_0_reg_168_NO_SHIFT_REG;
 logic rnode_1to168_indvars_iv_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_1to168_indvars_iv_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_1to168_indvars_iv_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_1to168_indvars_iv_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to168_indvars_iv_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to168_indvars_iv_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_1to168_indvars_iv_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_1to168_indvars_iv_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(local_lvm_indvars_iv_NO_SHIFT_REG),
	.data_out(rnode_1to168_indvars_iv_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_1to168_indvars_iv_0_reg_168_fifo.DEPTH = 168;
defparam rnode_1to168_indvars_iv_0_reg_168_fifo.DATA_WIDTH = 64;
defparam rnode_1to168_indvars_iv_0_reg_168_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to168_indvars_iv_0_reg_168_fifo.IMPL = "ram";

assign rnode_1to168_indvars_iv_0_reg_168_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_3_NO_SHIFT_REG;
assign merge_node_stall_in_3 = rnode_1to168_indvars_iv_0_stall_out_reg_168_NO_SHIFT_REG;
assign rnode_1to168_indvars_iv_0_NO_SHIFT_REG = rnode_1to168_indvars_iv_0_reg_168_NO_SHIFT_REG;
assign rnode_1to168_indvars_iv_0_stall_in_reg_168_NO_SHIFT_REG = rnode_1to168_indvars_iv_0_stall_in_NO_SHIFT_REG;
assign rnode_1to168_indvars_iv_0_valid_out_NO_SHIFT_REG = rnode_1to168_indvars_iv_0_valid_out_reg_168_NO_SHIFT_REG;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_1to8_var__u8_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_1_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_reg_8_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_valid_out_0_reg_8_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_stall_in_0_reg_8_NO_SHIFT_REG;
 logic rnode_1to8_var__u8_0_stall_out_reg_8_NO_SHIFT_REG;
 reg rnode_1to8_var__u8_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to8_var__u8_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_1to8_var__u8_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to8_var__u8_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to8_var__u8_0_stall_in_0_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_1to8_var__u8_0_valid_out_0_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_1to8_var__u8_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_lvm_var__u8_NO_SHIFT_REG),
	.data_out(rnode_1to8_var__u8_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_1to8_var__u8_0_reg_8_fifo.DEPTH = 8;
defparam rnode_1to8_var__u8_0_reg_8_fifo.DATA_WIDTH = 1;
defparam rnode_1to8_var__u8_0_reg_8_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to8_var__u8_0_reg_8_fifo.IMPL = "ll_reg";

assign rnode_1to8_var__u8_0_reg_8_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_4_NO_SHIFT_REG;
assign merge_node_stall_in_4 = rnode_1to8_var__u8_0_stall_out_reg_8_NO_SHIFT_REG;
assign rnode_1to8_var__u8_0_stall_in_0_reg_8_NO_SHIFT_REG = ((rnode_1to8_var__u8_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to8_var__u8_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to8_var__u8_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to8_var__u8_0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to8_var__u8_0_valid_out_0_NO_SHIFT_REG = (rnode_1to8_var__u8_0_valid_out_0_reg_8_NO_SHIFT_REG & ~(rnode_1to8_var__u8_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to8_var__u8_0_valid_out_1_NO_SHIFT_REG = (rnode_1to8_var__u8_0_valid_out_0_reg_8_NO_SHIFT_REG & ~(rnode_1to8_var__u8_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to8_var__u8_0_NO_SHIFT_REG = rnode_1to8_var__u8_0_reg_8_NO_SHIFT_REG;
assign rnode_1to8_var__u8_1_NO_SHIFT_REG = rnode_1to8_var__u8_0_reg_8_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to8_var__u8_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to8_var__u8_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to8_var__u8_0_consumed_0_NO_SHIFT_REG <= (rnode_1to8_var__u8_0_valid_out_0_reg_8_NO_SHIFT_REG & (rnode_1to8_var__u8_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to8_var__u8_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to8_var__u8_0_stall_in_0_reg_8_NO_SHIFT_REG);
		rnode_1to8_var__u8_0_consumed_1_NO_SHIFT_REG <= (rnode_1to8_var__u8_0_valid_out_0_reg_8_NO_SHIFT_REG & (rnode_1to8_var__u8_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to8_var__u8_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to8_var__u8_0_stall_in_0_reg_8_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_1to6_sub25_add24_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to6_sub25_add24_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to6_sub25_add24_0_NO_SHIFT_REG;
 logic rnode_1to6_sub25_add24_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to6_sub25_add24_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to6_sub25_add24_1_NO_SHIFT_REG;
 logic rnode_1to6_sub25_add24_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to6_sub25_add24_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_sub25_add24_0_valid_out_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_sub25_add24_0_stall_in_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_sub25_add24_0_stall_out_reg_6_NO_SHIFT_REG;
 reg rnode_1to6_sub25_add24_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to6_sub25_add24_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_1to6_sub25_add24_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to6_sub25_add24_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to6_sub25_add24_0_stall_in_0_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_1to6_sub25_add24_0_valid_out_0_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_1to6_sub25_add24_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_lvm_sub25_add24_NO_SHIFT_REG),
	.data_out(rnode_1to6_sub25_add24_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_1to6_sub25_add24_0_reg_6_fifo.DEPTH = 6;
defparam rnode_1to6_sub25_add24_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_1to6_sub25_add24_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to6_sub25_add24_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_1to6_sub25_add24_0_reg_6_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign merge_node_stall_in_5 = rnode_1to6_sub25_add24_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_1to6_sub25_add24_0_stall_in_0_reg_6_NO_SHIFT_REG = ((rnode_1to6_sub25_add24_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to6_sub25_add24_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to6_sub25_add24_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to6_sub25_add24_0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to6_sub25_add24_0_valid_out_0_NO_SHIFT_REG = (rnode_1to6_sub25_add24_0_valid_out_0_reg_6_NO_SHIFT_REG & ~(rnode_1to6_sub25_add24_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to6_sub25_add24_0_valid_out_1_NO_SHIFT_REG = (rnode_1to6_sub25_add24_0_valid_out_0_reg_6_NO_SHIFT_REG & ~(rnode_1to6_sub25_add24_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to6_sub25_add24_0_NO_SHIFT_REG = rnode_1to6_sub25_add24_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_sub25_add24_1_NO_SHIFT_REG = rnode_1to6_sub25_add24_0_reg_6_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to6_sub25_add24_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to6_sub25_add24_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to6_sub25_add24_0_consumed_0_NO_SHIFT_REG <= (rnode_1to6_sub25_add24_0_valid_out_0_reg_6_NO_SHIFT_REG & (rnode_1to6_sub25_add24_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to6_sub25_add24_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to6_sub25_add24_0_stall_in_0_reg_6_NO_SHIFT_REG);
		rnode_1to6_sub25_add24_0_consumed_1_NO_SHIFT_REG <= (rnode_1to6_sub25_add24_0_valid_out_0_reg_6_NO_SHIFT_REG & (rnode_1to6_sub25_add24_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to6_sub25_add24_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to6_sub25_add24_0_stall_in_0_reg_6_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 169
//  * capacity = 169
 logic rnode_1to170_arrayidx43_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to170_arrayidx43_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_1to170_arrayidx43_0_NO_SHIFT_REG;
 logic rnode_1to170_arrayidx43_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to170_arrayidx43_0_reg_170_NO_SHIFT_REG;
 logic rnode_1to170_arrayidx43_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_1to170_arrayidx43_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_1to170_arrayidx43_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_1to170_arrayidx43_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to170_arrayidx43_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to170_arrayidx43_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_1to170_arrayidx43_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_1to170_arrayidx43_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in((local_lvm_arrayidx43_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_1to170_arrayidx43_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_1to170_arrayidx43_0_reg_170_fifo.DEPTH = 170;
defparam rnode_1to170_arrayidx43_0_reg_170_fifo.DATA_WIDTH = 64;
defparam rnode_1to170_arrayidx43_0_reg_170_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to170_arrayidx43_0_reg_170_fifo.IMPL = "ram";

assign rnode_1to170_arrayidx43_0_reg_170_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_6_NO_SHIFT_REG;
assign merge_node_stall_in_6 = rnode_1to170_arrayidx43_0_stall_out_reg_170_NO_SHIFT_REG;
assign rnode_1to170_arrayidx43_0_NO_SHIFT_REG = rnode_1to170_arrayidx43_0_reg_170_NO_SHIFT_REG;
assign rnode_1to170_arrayidx43_0_stall_in_reg_170_NO_SHIFT_REG = rnode_1to170_arrayidx43_0_stall_in_NO_SHIFT_REG;
assign rnode_1to170_arrayidx43_0_valid_out_NO_SHIFT_REG = rnode_1to170_arrayidx43_0_valid_out_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 329
//  * capacity = 329
 logic rnode_1to330_ld__0_valid_out_NO_SHIFT_REG;
 logic rnode_1to330_ld__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to330_ld__0_NO_SHIFT_REG;
 logic rnode_1to330_ld__0_reg_330_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to330_ld__0_reg_330_NO_SHIFT_REG;
 logic rnode_1to330_ld__0_valid_out_reg_330_NO_SHIFT_REG;
 logic rnode_1to330_ld__0_stall_in_reg_330_NO_SHIFT_REG;
 logic rnode_1to330_ld__0_stall_out_reg_330_NO_SHIFT_REG;
wire [63:0] rci_rcnode_1to330_rc8_t_119_0_reg_1;

acl_data_fifo rnode_1to330_ld__0_reg_330_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to330_ld__0_reg_330_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to330_ld__0_stall_in_reg_330_NO_SHIFT_REG),
	.valid_out(rnode_1to330_ld__0_valid_out_reg_330_NO_SHIFT_REG),
	.stall_out(rnode_1to330_ld__0_stall_out_reg_330_NO_SHIFT_REG),
	.data_in(local_lvm_ld__NO_SHIFT_REG),
	.data_out(rnode_1to330_ld__0_reg_330_NO_SHIFT_REG)
);

defparam rnode_1to330_ld__0_reg_330_fifo.DEPTH = 330;
defparam rnode_1to330_ld__0_reg_330_fifo.DATA_WIDTH = 32;
defparam rnode_1to330_ld__0_reg_330_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to330_ld__0_reg_330_fifo.IMPL = "ram";

assign rnode_1to330_ld__0_reg_330_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_7_NO_SHIFT_REG;
assign merge_node_stall_in_7 = rnode_1to330_ld__0_stall_out_reg_330_NO_SHIFT_REG;
assign rnode_1to330_ld__0_NO_SHIFT_REG = rnode_1to330_ld__0_reg_330_NO_SHIFT_REG;
assign rnode_1to330_ld__0_stall_in_reg_330_NO_SHIFT_REG = rnode_1to330_ld__0_stall_in_NO_SHIFT_REG;
assign rnode_1to330_ld__0_valid_out_NO_SHIFT_REG = rnode_1to330_ld__0_valid_out_reg_330_NO_SHIFT_REG;
assign rci_rcnode_1to330_rc8_t_119_0_reg_1[31:0] = local_lvm_t_119_NO_SHIFT_REG;
assign rci_rcnode_1to330_rc8_t_119_0_reg_1[63:32] = local_lvm_sum_118_NO_SHIFT_REG;

// Register node:
//  * latency = 329
//  * capacity = 329
 logic rcnode_1to330_rc8_t_119_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to330_rc8_t_119_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rcnode_1to330_rc8_t_119_0_NO_SHIFT_REG;
 logic rcnode_1to330_rc8_t_119_0_reg_330_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rcnode_1to330_rc8_t_119_0_reg_330_NO_SHIFT_REG;
 logic rcnode_1to330_rc8_t_119_0_valid_out_reg_330_NO_SHIFT_REG;
 logic rcnode_1to330_rc8_t_119_0_stall_in_reg_330_NO_SHIFT_REG;
 logic rcnode_1to330_rc8_t_119_0_stall_out_reg_330_IP_NO_SHIFT_REG;
 logic rcnode_1to330_rc8_t_119_0_stall_out_reg_330_NO_SHIFT_REG;
wire [160:0] rci_rcnode_1to398_rc9_idxprom_0_reg_1;

acl_data_fifo rcnode_1to330_rc8_t_119_0_reg_330_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to330_rc8_t_119_0_reg_330_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to330_rc8_t_119_0_stall_in_reg_330_NO_SHIFT_REG),
	.valid_out(rcnode_1to330_rc8_t_119_0_valid_out_reg_330_NO_SHIFT_REG),
	.stall_out(rcnode_1to330_rc8_t_119_0_stall_out_reg_330_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to330_rc8_t_119_0_reg_1),
	.data_out(rcnode_1to330_rc8_t_119_0_reg_330_NO_SHIFT_REG)
);

defparam rcnode_1to330_rc8_t_119_0_reg_330_fifo.DEPTH = 330;
defparam rcnode_1to330_rc8_t_119_0_reg_330_fifo.DATA_WIDTH = 64;
defparam rcnode_1to330_rc8_t_119_0_reg_330_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to330_rc8_t_119_0_reg_330_fifo.IMPL = "ram";

assign rcnode_1to330_rc8_t_119_0_reg_330_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_8_NO_SHIFT_REG;
assign rcnode_1to330_rc8_t_119_0_stall_out_reg_330_NO_SHIFT_REG = (~(rcnode_1to330_rc8_t_119_0_reg_330_inputs_ready_NO_SHIFT_REG) | rcnode_1to330_rc8_t_119_0_stall_out_reg_330_IP_NO_SHIFT_REG);
assign merge_node_stall_in_8 = rcnode_1to330_rc8_t_119_0_stall_out_reg_330_NO_SHIFT_REG;
assign rcnode_1to330_rc8_t_119_0_NO_SHIFT_REG = rcnode_1to330_rc8_t_119_0_reg_330_NO_SHIFT_REG;
assign rcnode_1to330_rc8_t_119_0_stall_in_reg_330_NO_SHIFT_REG = rcnode_1to330_rc8_t_119_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to330_rc8_t_119_0_valid_out_NO_SHIFT_REG = rcnode_1to330_rc8_t_119_0_valid_out_reg_330_NO_SHIFT_REG;
assign rci_rcnode_1to398_rc9_idxprom_0_reg_1[63:0] = (local_lvm_idxprom_NO_SHIFT_REG & 64'hFFFFFFFF);
assign rci_rcnode_1to398_rc9_idxprom_0_reg_1[64] = local_lvm_cmp_NO_SHIFT_REG;
assign rci_rcnode_1to398_rc9_idxprom_0_reg_1[128:65] = local_lvm_indvars_iv29_NO_SHIFT_REG;
assign rci_rcnode_1to398_rc9_idxprom_0_reg_1[160:129] = local_lvm_input_global_id_0_NO_SHIFT_REG;

// Register node:
//  * latency = 397
//  * capacity = 397
 logic rcnode_1to398_rc9_idxprom_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to398_rc9_idxprom_0_stall_in_NO_SHIFT_REG;
 logic [160:0] rcnode_1to398_rc9_idxprom_0_NO_SHIFT_REG;
 logic rcnode_1to398_rc9_idxprom_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [160:0] rcnode_1to398_rc9_idxprom_0_reg_398_NO_SHIFT_REG;
 logic rcnode_1to398_rc9_idxprom_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rcnode_1to398_rc9_idxprom_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rcnode_1to398_rc9_idxprom_0_stall_out_reg_398_IP_NO_SHIFT_REG;
 logic rcnode_1to398_rc9_idxprom_0_stall_out_reg_398_NO_SHIFT_REG;
wire [63:0] rci_rcnode_1to398_rc10_input_global_id_1_0_reg_1;

acl_data_fifo rcnode_1to398_rc9_idxprom_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to398_rc9_idxprom_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to398_rc9_idxprom_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rcnode_1to398_rc9_idxprom_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rcnode_1to398_rc9_idxprom_0_stall_out_reg_398_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to398_rc9_idxprom_0_reg_1),
	.data_out(rcnode_1to398_rc9_idxprom_0_reg_398_NO_SHIFT_REG)
);

defparam rcnode_1to398_rc9_idxprom_0_reg_398_fifo.DEPTH = 398;
defparam rcnode_1to398_rc9_idxprom_0_reg_398_fifo.DATA_WIDTH = 161;
defparam rcnode_1to398_rc9_idxprom_0_reg_398_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to398_rc9_idxprom_0_reg_398_fifo.IMPL = "ram";

assign rcnode_1to398_rc9_idxprom_0_reg_398_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_9_NO_SHIFT_REG;
assign rcnode_1to398_rc9_idxprom_0_stall_out_reg_398_NO_SHIFT_REG = (~(rcnode_1to398_rc9_idxprom_0_reg_398_inputs_ready_NO_SHIFT_REG) | rcnode_1to398_rc9_idxprom_0_stall_out_reg_398_IP_NO_SHIFT_REG);
assign merge_node_stall_in_9 = rcnode_1to398_rc9_idxprom_0_stall_out_reg_398_NO_SHIFT_REG;
assign rcnode_1to398_rc9_idxprom_0_NO_SHIFT_REG = rcnode_1to398_rc9_idxprom_0_reg_398_NO_SHIFT_REG;
assign rcnode_1to398_rc9_idxprom_0_stall_in_reg_398_NO_SHIFT_REG = rcnode_1to398_rc9_idxprom_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to398_rc9_idxprom_0_valid_out_NO_SHIFT_REG = rcnode_1to398_rc9_idxprom_0_valid_out_reg_398_NO_SHIFT_REG;
assign rci_rcnode_1to398_rc10_input_global_id_1_0_reg_1[31:0] = local_lvm_input_global_id_1_NO_SHIFT_REG;
assign rci_rcnode_1to398_rc10_input_global_id_1_0_reg_1[63:32] = local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;

// Register node:
//  * latency = 397
//  * capacity = 397
 logic rcnode_1to398_rc10_input_global_id_1_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to398_rc10_input_global_id_1_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rcnode_1to398_rc10_input_global_id_1_0_NO_SHIFT_REG;
 logic rcnode_1to398_rc10_input_global_id_1_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rcnode_1to398_rc10_input_global_id_1_0_reg_398_NO_SHIFT_REG;
 logic rcnode_1to398_rc10_input_global_id_1_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rcnode_1to398_rc10_input_global_id_1_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rcnode_1to398_rc10_input_global_id_1_0_stall_out_reg_398_IP_NO_SHIFT_REG;
 logic rcnode_1to398_rc10_input_global_id_1_0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rcnode_1to398_rc10_input_global_id_1_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to398_rc10_input_global_id_1_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to398_rc10_input_global_id_1_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rcnode_1to398_rc10_input_global_id_1_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rcnode_1to398_rc10_input_global_id_1_0_stall_out_reg_398_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to398_rc10_input_global_id_1_0_reg_1),
	.data_out(rcnode_1to398_rc10_input_global_id_1_0_reg_398_NO_SHIFT_REG)
);

defparam rcnode_1to398_rc10_input_global_id_1_0_reg_398_fifo.DEPTH = 398;
defparam rcnode_1to398_rc10_input_global_id_1_0_reg_398_fifo.DATA_WIDTH = 64;
defparam rcnode_1to398_rc10_input_global_id_1_0_reg_398_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to398_rc10_input_global_id_1_0_reg_398_fifo.IMPL = "ram";

assign rcnode_1to398_rc10_input_global_id_1_0_reg_398_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_10_NO_SHIFT_REG;
assign rcnode_1to398_rc10_input_global_id_1_0_stall_out_reg_398_NO_SHIFT_REG = (~(rcnode_1to398_rc10_input_global_id_1_0_reg_398_inputs_ready_NO_SHIFT_REG) | rcnode_1to398_rc10_input_global_id_1_0_stall_out_reg_398_IP_NO_SHIFT_REG);
assign merge_node_stall_in_10 = rcnode_1to398_rc10_input_global_id_1_0_stall_out_reg_398_NO_SHIFT_REG;
assign rcnode_1to398_rc10_input_global_id_1_0_NO_SHIFT_REG = rcnode_1to398_rc10_input_global_id_1_0_reg_398_NO_SHIFT_REG;
assign rcnode_1to398_rc10_input_global_id_1_0_stall_in_reg_398_NO_SHIFT_REG = rcnode_1to398_rc10_input_global_id_1_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to398_rc10_input_global_id_1_0_valid_out_NO_SHIFT_REG = rcnode_1to398_rc10_input_global_id_1_0_valid_out_reg_398_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_add28_valid_out;
wire local_bb3_add28_stall_in;
wire local_bb3_add28_inputs_ready;
wire local_bb3_add28_stall_local;
wire [31:0] local_bb3_add28;

assign local_bb3_add28_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign local_bb3_add28 = (local_bb3_var_ + local_lvm_input_global_id_1_NO_SHIFT_REG);
assign local_bb3_add28_valid_out = local_bb3_add28_inputs_ready;
assign local_bb3_add28_stall_local = local_bb3_add28_stall_in;
assign merge_node_stall_in_0 = (local_bb3_add28_stall_local | ~(local_bb3_add28_inputs_ready));
assign merge_node_stall_in_1 = (local_bb3_add28_stall_local | ~(local_bb3_add28_inputs_ready));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_var__u7_0_valid_out_NO_SHIFT_REG;
 logic rnode_168to169_var__u7_0_stall_in_NO_SHIFT_REG;
 logic rnode_168to169_var__u7_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_168to169_var__u7_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_var__u7_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_var__u7_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_var__u7_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_var__u7_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_var__u7_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_var__u7_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_var__u7_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_168to169_var__u7_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_var__u7_0_reg_169_fifo.DATA_WIDTH = 0;
defparam rnode_168to169_var__u7_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_var__u7_0_reg_169_fifo.IMPL = "ll_reg";

assign rnode_168to169_var__u7_0_reg_169_inputs_ready_NO_SHIFT_REG = rnode_1to168_var__u7_0_valid_out_NO_SHIFT_REG;
assign rnode_1to168_var__u7_0_stall_in_NO_SHIFT_REG = rnode_168to169_var__u7_0_stall_out_reg_169_NO_SHIFT_REG;
assign rnode_168to169_var__u7_0_stall_in_reg_169_NO_SHIFT_REG = rnode_168to169_var__u7_0_stall_in_NO_SHIFT_REG;
assign rnode_168to169_var__u7_0_valid_out_NO_SHIFT_REG = rnode_168to169_var__u7_0_valid_out_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_indvars_iv_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_indvars_iv_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_168to169_indvars_iv_0_NO_SHIFT_REG;
 logic rnode_168to169_indvars_iv_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_indvars_iv_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_168to169_indvars_iv_1_NO_SHIFT_REG;
 logic rnode_168to169_indvars_iv_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_168to169_indvars_iv_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_indvars_iv_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_indvars_iv_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_indvars_iv_0_stall_out_reg_169_NO_SHIFT_REG;
 reg rnode_168to169_indvars_iv_0_consumed_0_NO_SHIFT_REG;
 reg rnode_168to169_indvars_iv_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_indvars_iv_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_indvars_iv_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_indvars_iv_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_indvars_iv_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_indvars_iv_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_1to168_indvars_iv_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_indvars_iv_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_indvars_iv_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_indvars_iv_0_reg_169_fifo.DATA_WIDTH = 64;
defparam rnode_168to169_indvars_iv_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_indvars_iv_0_reg_169_fifo.IMPL = "ll_reg";

assign rnode_168to169_indvars_iv_0_reg_169_inputs_ready_NO_SHIFT_REG = rnode_1to168_indvars_iv_0_valid_out_NO_SHIFT_REG;
assign rnode_1to168_indvars_iv_0_stall_in_NO_SHIFT_REG = rnode_168to169_indvars_iv_0_stall_out_reg_169_NO_SHIFT_REG;
assign rnode_168to169_indvars_iv_0_stall_in_0_reg_169_NO_SHIFT_REG = ((rnode_168to169_indvars_iv_0_stall_in_0_NO_SHIFT_REG & ~(rnode_168to169_indvars_iv_0_consumed_0_NO_SHIFT_REG)) | (rnode_168to169_indvars_iv_0_stall_in_1_NO_SHIFT_REG & ~(rnode_168to169_indvars_iv_0_consumed_1_NO_SHIFT_REG)));
assign rnode_168to169_indvars_iv_0_valid_out_0_NO_SHIFT_REG = (rnode_168to169_indvars_iv_0_valid_out_0_reg_169_NO_SHIFT_REG & ~(rnode_168to169_indvars_iv_0_consumed_0_NO_SHIFT_REG));
assign rnode_168to169_indvars_iv_0_valid_out_1_NO_SHIFT_REG = (rnode_168to169_indvars_iv_0_valid_out_0_reg_169_NO_SHIFT_REG & ~(rnode_168to169_indvars_iv_0_consumed_1_NO_SHIFT_REG));
assign rnode_168to169_indvars_iv_0_NO_SHIFT_REG = rnode_168to169_indvars_iv_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_indvars_iv_1_NO_SHIFT_REG = rnode_168to169_indvars_iv_0_reg_169_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_168to169_indvars_iv_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_168to169_indvars_iv_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_168to169_indvars_iv_0_consumed_0_NO_SHIFT_REG <= (rnode_168to169_indvars_iv_0_valid_out_0_reg_169_NO_SHIFT_REG & (rnode_168to169_indvars_iv_0_consumed_0_NO_SHIFT_REG | ~(rnode_168to169_indvars_iv_0_stall_in_0_NO_SHIFT_REG)) & rnode_168to169_indvars_iv_0_stall_in_0_reg_169_NO_SHIFT_REG);
		rnode_168to169_indvars_iv_0_consumed_1_NO_SHIFT_REG <= (rnode_168to169_indvars_iv_0_valid_out_0_reg_169_NO_SHIFT_REG & (rnode_168to169_indvars_iv_0_consumed_1_NO_SHIFT_REG | ~(rnode_168to169_indvars_iv_0_stall_in_1_NO_SHIFT_REG)) & rnode_168to169_indvars_iv_0_stall_in_0_reg_169_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_8to170_var__u8_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to170_var__u8_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to170_var__u8_0_NO_SHIFT_REG;
 logic rnode_8to170_var__u8_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to170_var__u8_0_reg_170_NO_SHIFT_REG;
 logic rnode_8to170_var__u8_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_8to170_var__u8_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_8to170_var__u8_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_8to170_var__u8_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to170_var__u8_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to170_var__u8_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_8to170_var__u8_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_8to170_var__u8_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_1to8_var__u8_1_NO_SHIFT_REG),
	.data_out(rnode_8to170_var__u8_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_8to170_var__u8_0_reg_170_fifo.DEPTH = 163;
defparam rnode_8to170_var__u8_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_8to170_var__u8_0_reg_170_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_8to170_var__u8_0_reg_170_fifo.IMPL = "ram";

assign rnode_8to170_var__u8_0_reg_170_inputs_ready_NO_SHIFT_REG = rnode_1to8_var__u8_0_valid_out_1_NO_SHIFT_REG;
assign rnode_1to8_var__u8_0_stall_in_1_NO_SHIFT_REG = rnode_8to170_var__u8_0_stall_out_reg_170_NO_SHIFT_REG;
assign rnode_8to170_var__u8_0_NO_SHIFT_REG = rnode_8to170_var__u8_0_reg_170_NO_SHIFT_REG;
assign rnode_8to170_var__u8_0_stall_in_reg_170_NO_SHIFT_REG = rnode_8to170_var__u8_0_stall_in_NO_SHIFT_REG;
assign rnode_8to170_var__u8_0_valid_out_NO_SHIFT_REG = rnode_8to170_var__u8_0_valid_out_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 392
//  * capacity = 392
 logic rnode_6to398_sub25_add24_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to398_sub25_add24_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_6to398_sub25_add24_0_NO_SHIFT_REG;
 logic rnode_6to398_sub25_add24_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_6to398_sub25_add24_0_reg_398_NO_SHIFT_REG;
 logic rnode_6to398_sub25_add24_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rnode_6to398_sub25_add24_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rnode_6to398_sub25_add24_0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_6to398_sub25_add24_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to398_sub25_add24_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to398_sub25_add24_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_6to398_sub25_add24_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_6to398_sub25_add24_0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(rnode_1to6_sub25_add24_1_NO_SHIFT_REG),
	.data_out(rnode_6to398_sub25_add24_0_reg_398_NO_SHIFT_REG)
);

defparam rnode_6to398_sub25_add24_0_reg_398_fifo.DEPTH = 393;
defparam rnode_6to398_sub25_add24_0_reg_398_fifo.DATA_WIDTH = 32;
defparam rnode_6to398_sub25_add24_0_reg_398_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_6to398_sub25_add24_0_reg_398_fifo.IMPL = "ram";

assign rnode_6to398_sub25_add24_0_reg_398_inputs_ready_NO_SHIFT_REG = rnode_1to6_sub25_add24_0_valid_out_1_NO_SHIFT_REG;
assign rnode_1to6_sub25_add24_0_stall_in_1_NO_SHIFT_REG = rnode_6to398_sub25_add24_0_stall_out_reg_398_NO_SHIFT_REG;
assign rnode_6to398_sub25_add24_0_NO_SHIFT_REG = rnode_6to398_sub25_add24_0_reg_398_NO_SHIFT_REG;
assign rnode_6to398_sub25_add24_0_stall_in_reg_398_NO_SHIFT_REG = rnode_6to398_sub25_add24_0_stall_in_NO_SHIFT_REG;
assign rnode_6to398_sub25_add24_0_valid_out_NO_SHIFT_REG = rnode_6to398_sub25_add24_0_valid_out_reg_398_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_arrayidx43_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_arrayidx43_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_170to171_arrayidx43_0_NO_SHIFT_REG;
 logic rnode_170to171_arrayidx43_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_arrayidx43_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_170to171_arrayidx43_1_NO_SHIFT_REG;
 logic rnode_170to171_arrayidx43_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_170to171_arrayidx43_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_arrayidx43_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_arrayidx43_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_arrayidx43_0_stall_out_reg_171_NO_SHIFT_REG;
 reg rnode_170to171_arrayidx43_0_consumed_0_NO_SHIFT_REG;
 reg rnode_170to171_arrayidx43_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_arrayidx43_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_arrayidx43_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_arrayidx43_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_arrayidx43_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_arrayidx43_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in((rnode_1to170_arrayidx43_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_170to171_arrayidx43_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_arrayidx43_0_reg_171_fifo.DEPTH = 2;
defparam rnode_170to171_arrayidx43_0_reg_171_fifo.DATA_WIDTH = 64;
defparam rnode_170to171_arrayidx43_0_reg_171_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_170to171_arrayidx43_0_reg_171_fifo.IMPL = "ll_reg";

assign rnode_170to171_arrayidx43_0_reg_171_inputs_ready_NO_SHIFT_REG = rnode_1to170_arrayidx43_0_valid_out_NO_SHIFT_REG;
assign rnode_1to170_arrayidx43_0_stall_in_NO_SHIFT_REG = rnode_170to171_arrayidx43_0_stall_out_reg_171_NO_SHIFT_REG;
assign rnode_170to171_arrayidx43_0_stall_in_0_reg_171_NO_SHIFT_REG = ((rnode_170to171_arrayidx43_0_stall_in_0_NO_SHIFT_REG & ~(rnode_170to171_arrayidx43_0_consumed_0_NO_SHIFT_REG)) | (rnode_170to171_arrayidx43_0_stall_in_1_NO_SHIFT_REG & ~(rnode_170to171_arrayidx43_0_consumed_1_NO_SHIFT_REG)));
assign rnode_170to171_arrayidx43_0_valid_out_0_NO_SHIFT_REG = (rnode_170to171_arrayidx43_0_valid_out_0_reg_171_NO_SHIFT_REG & ~(rnode_170to171_arrayidx43_0_consumed_0_NO_SHIFT_REG));
assign rnode_170to171_arrayidx43_0_valid_out_1_NO_SHIFT_REG = (rnode_170to171_arrayidx43_0_valid_out_0_reg_171_NO_SHIFT_REG & ~(rnode_170to171_arrayidx43_0_consumed_1_NO_SHIFT_REG));
assign rnode_170to171_arrayidx43_0_NO_SHIFT_REG = rnode_170to171_arrayidx43_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_arrayidx43_1_NO_SHIFT_REG = rnode_170to171_arrayidx43_0_reg_171_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_170to171_arrayidx43_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_170to171_arrayidx43_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_170to171_arrayidx43_0_consumed_0_NO_SHIFT_REG <= (rnode_170to171_arrayidx43_0_valid_out_0_reg_171_NO_SHIFT_REG & (rnode_170to171_arrayidx43_0_consumed_0_NO_SHIFT_REG | ~(rnode_170to171_arrayidx43_0_stall_in_0_NO_SHIFT_REG)) & rnode_170to171_arrayidx43_0_stall_in_0_reg_171_NO_SHIFT_REG);
		rnode_170to171_arrayidx43_0_consumed_1_NO_SHIFT_REG <= (rnode_170to171_arrayidx43_0_valid_out_0_reg_171_NO_SHIFT_REG & (rnode_170to171_arrayidx43_0_consumed_1_NO_SHIFT_REG | ~(rnode_170to171_arrayidx43_0_stall_in_1_NO_SHIFT_REG)) & rnode_170to171_arrayidx43_0_stall_in_0_reg_171_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_330to331_ld__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_330to331_ld__0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_330to331_ld__0_NO_SHIFT_REG;
 logic rnode_330to331_ld__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_330to331_ld__0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_330to331_ld__1_NO_SHIFT_REG;
 logic rnode_330to331_ld__0_reg_331_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_330to331_ld__0_reg_331_NO_SHIFT_REG;
 logic rnode_330to331_ld__0_valid_out_0_reg_331_NO_SHIFT_REG;
 logic rnode_330to331_ld__0_stall_in_0_reg_331_NO_SHIFT_REG;
 logic rnode_330to331_ld__0_stall_out_reg_331_NO_SHIFT_REG;
 reg rnode_330to331_ld__0_consumed_0_NO_SHIFT_REG;
 reg rnode_330to331_ld__0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_330to331_ld__0_reg_331_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_330to331_ld__0_reg_331_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_330to331_ld__0_stall_in_0_reg_331_NO_SHIFT_REG),
	.valid_out(rnode_330to331_ld__0_valid_out_0_reg_331_NO_SHIFT_REG),
	.stall_out(rnode_330to331_ld__0_stall_out_reg_331_NO_SHIFT_REG),
	.data_in(rnode_1to330_ld__0_NO_SHIFT_REG),
	.data_out(rnode_330to331_ld__0_reg_331_NO_SHIFT_REG)
);

defparam rnode_330to331_ld__0_reg_331_fifo.DEPTH = 1;
defparam rnode_330to331_ld__0_reg_331_fifo.DATA_WIDTH = 32;
defparam rnode_330to331_ld__0_reg_331_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_330to331_ld__0_reg_331_fifo.IMPL = "ll_reg";

assign rnode_330to331_ld__0_reg_331_inputs_ready_NO_SHIFT_REG = rnode_1to330_ld__0_valid_out_NO_SHIFT_REG;
assign rnode_1to330_ld__0_stall_in_NO_SHIFT_REG = rnode_330to331_ld__0_stall_out_reg_331_NO_SHIFT_REG;
assign rnode_330to331_ld__0_stall_in_0_reg_331_NO_SHIFT_REG = ((rnode_330to331_ld__0_stall_in_0_NO_SHIFT_REG & ~(rnode_330to331_ld__0_consumed_0_NO_SHIFT_REG)) | (rnode_330to331_ld__0_stall_in_1_NO_SHIFT_REG & ~(rnode_330to331_ld__0_consumed_1_NO_SHIFT_REG)));
assign rnode_330to331_ld__0_valid_out_0_NO_SHIFT_REG = (rnode_330to331_ld__0_valid_out_0_reg_331_NO_SHIFT_REG & ~(rnode_330to331_ld__0_consumed_0_NO_SHIFT_REG));
assign rnode_330to331_ld__0_valid_out_1_NO_SHIFT_REG = (rnode_330to331_ld__0_valid_out_0_reg_331_NO_SHIFT_REG & ~(rnode_330to331_ld__0_consumed_1_NO_SHIFT_REG));
assign rnode_330to331_ld__0_NO_SHIFT_REG = rnode_330to331_ld__0_reg_331_NO_SHIFT_REG;
assign rnode_330to331_ld__1_NO_SHIFT_REG = rnode_330to331_ld__0_reg_331_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_330to331_ld__0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_330to331_ld__0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_330to331_ld__0_consumed_0_NO_SHIFT_REG <= (rnode_330to331_ld__0_valid_out_0_reg_331_NO_SHIFT_REG & (rnode_330to331_ld__0_consumed_0_NO_SHIFT_REG | ~(rnode_330to331_ld__0_stall_in_0_NO_SHIFT_REG)) & rnode_330to331_ld__0_stall_in_0_reg_331_NO_SHIFT_REG);
		rnode_330to331_ld__0_consumed_1_NO_SHIFT_REG <= (rnode_330to331_ld__0_valid_out_0_reg_331_NO_SHIFT_REG & (rnode_330to331_ld__0_consumed_1_NO_SHIFT_REG | ~(rnode_330to331_ld__0_stall_in_1_NO_SHIFT_REG)) & rnode_330to331_ld__0_stall_in_0_reg_331_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_add28_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add28_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_add28_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add28_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add28_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_add28_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add28_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_add28_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add28_0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add28_0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add28_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_add28_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_add28_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_add28_0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_add28_0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_add28_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_add28),
	.data_out(rnode_1to2_bb3_add28_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_add28_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_add28_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb3_add28_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_add28_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb3_add28_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb3_add28_valid_out;
assign local_bb3_add28_stall_in = rnode_1to2_bb3_add28_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_add28_0_stall_in_0_reg_2_NO_SHIFT_REG = (rnode_1to2_bb3_add28_0_stall_in_0_NO_SHIFT_REG | rnode_1to2_bb3_add28_0_stall_in_1_NO_SHIFT_REG);
assign rnode_1to2_bb3_add28_0_valid_out_0_NO_SHIFT_REG = rnode_1to2_bb3_add28_0_valid_out_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_add28_0_valid_out_1_NO_SHIFT_REG = rnode_1to2_bb3_add28_0_valid_out_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_add28_0_NO_SHIFT_REG = rnode_1to2_bb3_add28_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_add28_1_NO_SHIFT_REG = rnode_1to2_bb3_add28_0_reg_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u9_valid_out;
wire local_bb3_var__u9_stall_in;
wire local_bb3_var__u9_inputs_ready;
wire local_bb3_var__u9_stall_local;
wire [63:0] local_bb3_var__u9;

assign local_bb3_var__u9_inputs_ready = (rnode_168to169_var__u7_0_valid_out_NO_SHIFT_REG & rnode_168to169_indvars_iv_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3_var__u9 = (rnode_168to169_indvars_iv_0_NO_SHIFT_REG + input_wii_var__u7);
assign local_bb3_var__u9_valid_out = local_bb3_var__u9_inputs_ready;
assign local_bb3_var__u9_stall_local = local_bb3_var__u9_stall_in;
assign rnode_168to169_var__u7_0_stall_in_NO_SHIFT_REG = (local_bb3_var__u9_stall_local | ~(local_bb3_var__u9_inputs_ready));
assign rnode_168to169_indvars_iv_0_stall_in_0_NO_SHIFT_REG = (local_bb3_var__u9_stall_local | ~(local_bb3_var__u9_inputs_ready));

// Register node:
//  * latency = 227
//  * capacity = 227
 logic rnode_169to396_indvars_iv_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to396_indvars_iv_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_169to396_indvars_iv_0_NO_SHIFT_REG;
 logic rnode_169to396_indvars_iv_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_169to396_indvars_iv_0_reg_396_NO_SHIFT_REG;
 logic rnode_169to396_indvars_iv_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_169to396_indvars_iv_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_169to396_indvars_iv_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_169to396_indvars_iv_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to396_indvars_iv_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to396_indvars_iv_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_169to396_indvars_iv_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_169to396_indvars_iv_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(rnode_168to169_indvars_iv_1_NO_SHIFT_REG),
	.data_out(rnode_169to396_indvars_iv_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_169to396_indvars_iv_0_reg_396_fifo.DEPTH = 228;
defparam rnode_169to396_indvars_iv_0_reg_396_fifo.DATA_WIDTH = 64;
defparam rnode_169to396_indvars_iv_0_reg_396_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_169to396_indvars_iv_0_reg_396_fifo.IMPL = "ram";

assign rnode_169to396_indvars_iv_0_reg_396_inputs_ready_NO_SHIFT_REG = rnode_168to169_indvars_iv_0_valid_out_1_NO_SHIFT_REG;
assign rnode_168to169_indvars_iv_0_stall_in_1_NO_SHIFT_REG = rnode_169to396_indvars_iv_0_stall_out_reg_396_NO_SHIFT_REG;
assign rnode_169to396_indvars_iv_0_NO_SHIFT_REG = rnode_169to396_indvars_iv_0_reg_396_NO_SHIFT_REG;
assign rnode_169to396_indvars_iv_0_stall_in_reg_396_NO_SHIFT_REG = rnode_169to396_indvars_iv_0_stall_in_NO_SHIFT_REG;
assign rnode_169to396_indvars_iv_0_valid_out_NO_SHIFT_REG = rnode_169to396_indvars_iv_0_valid_out_reg_396_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_var__u8_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_1_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_var__u8_0_stall_out_reg_171_NO_SHIFT_REG;
 reg rnode_170to171_var__u8_0_consumed_0_NO_SHIFT_REG;
 reg rnode_170to171_var__u8_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_var__u8_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_var__u8_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_var__u8_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_var__u8_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_var__u8_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(rnode_8to170_var__u8_0_NO_SHIFT_REG),
	.data_out(rnode_170to171_var__u8_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_var__u8_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_var__u8_0_reg_171_fifo.DATA_WIDTH = 1;
defparam rnode_170to171_var__u8_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_var__u8_0_reg_171_fifo.IMPL = "ll_reg";

assign rnode_170to171_var__u8_0_reg_171_inputs_ready_NO_SHIFT_REG = rnode_8to170_var__u8_0_valid_out_NO_SHIFT_REG;
assign rnode_8to170_var__u8_0_stall_in_NO_SHIFT_REG = rnode_170to171_var__u8_0_stall_out_reg_171_NO_SHIFT_REG;
assign rnode_170to171_var__u8_0_stall_in_0_reg_171_NO_SHIFT_REG = ((rnode_170to171_var__u8_0_stall_in_0_NO_SHIFT_REG & ~(rnode_170to171_var__u8_0_consumed_0_NO_SHIFT_REG)) | (rnode_170to171_var__u8_0_stall_in_1_NO_SHIFT_REG & ~(rnode_170to171_var__u8_0_consumed_1_NO_SHIFT_REG)));
assign rnode_170to171_var__u8_0_valid_out_0_NO_SHIFT_REG = (rnode_170to171_var__u8_0_valid_out_0_reg_171_NO_SHIFT_REG & ~(rnode_170to171_var__u8_0_consumed_0_NO_SHIFT_REG));
assign rnode_170to171_var__u8_0_valid_out_1_NO_SHIFT_REG = (rnode_170to171_var__u8_0_valid_out_0_reg_171_NO_SHIFT_REG & ~(rnode_170to171_var__u8_0_consumed_1_NO_SHIFT_REG));
assign rnode_170to171_var__u8_0_NO_SHIFT_REG = rnode_170to171_var__u8_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_var__u8_1_NO_SHIFT_REG = rnode_170to171_var__u8_0_reg_171_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_170to171_var__u8_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_170to171_var__u8_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_170to171_var__u8_0_consumed_0_NO_SHIFT_REG <= (rnode_170to171_var__u8_0_valid_out_0_reg_171_NO_SHIFT_REG & (rnode_170to171_var__u8_0_consumed_0_NO_SHIFT_REG | ~(rnode_170to171_var__u8_0_stall_in_0_NO_SHIFT_REG)) & rnode_170to171_var__u8_0_stall_in_0_reg_171_NO_SHIFT_REG);
		rnode_170to171_var__u8_0_consumed_1_NO_SHIFT_REG <= (rnode_170to171_var__u8_0_valid_out_0_reg_171_NO_SHIFT_REG & (rnode_170to171_var__u8_0_consumed_1_NO_SHIFT_REG | ~(rnode_170to171_var__u8_0_stall_in_1_NO_SHIFT_REG)) & rnode_170to171_var__u8_0_stall_in_0_reg_171_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 67
//  * capacity = 67
 logic rnode_331to398_ld__0_valid_out_NO_SHIFT_REG;
 logic rnode_331to398_ld__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_331to398_ld__0_NO_SHIFT_REG;
 logic rnode_331to398_ld__0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_331to398_ld__0_reg_398_NO_SHIFT_REG;
 logic rnode_331to398_ld__0_valid_out_reg_398_NO_SHIFT_REG;
 logic rnode_331to398_ld__0_stall_in_reg_398_NO_SHIFT_REG;
 logic rnode_331to398_ld__0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_331to398_ld__0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_331to398_ld__0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_331to398_ld__0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_331to398_ld__0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_331to398_ld__0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(rnode_330to331_ld__1_NO_SHIFT_REG),
	.data_out(rnode_331to398_ld__0_reg_398_NO_SHIFT_REG)
);

defparam rnode_331to398_ld__0_reg_398_fifo.DEPTH = 68;
defparam rnode_331to398_ld__0_reg_398_fifo.DATA_WIDTH = 32;
defparam rnode_331to398_ld__0_reg_398_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_331to398_ld__0_reg_398_fifo.IMPL = "ram";

assign rnode_331to398_ld__0_reg_398_inputs_ready_NO_SHIFT_REG = rnode_330to331_ld__0_valid_out_1_NO_SHIFT_REG;
assign rnode_330to331_ld__0_stall_in_1_NO_SHIFT_REG = rnode_331to398_ld__0_stall_out_reg_398_NO_SHIFT_REG;
assign rnode_331to398_ld__0_NO_SHIFT_REG = rnode_331to398_ld__0_reg_398_NO_SHIFT_REG;
assign rnode_331to398_ld__0_stall_in_reg_398_NO_SHIFT_REG = rnode_331to398_ld__0_stall_in_NO_SHIFT_REG;
assign rnode_331to398_ld__0_valid_out_NO_SHIFT_REG = rnode_331to398_ld__0_valid_out_reg_398_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp1_i9_valid_out;
wire local_bb3_cmp1_i9_stall_in;
wire local_bb3_cmp1_i9_inputs_ready;
wire local_bb3_cmp1_i9_stall_local;
wire local_bb3_cmp1_i9;

assign local_bb3_cmp1_i9_inputs_ready = rnode_1to2_bb3_add28_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_cmp1_i9 = (rnode_1to2_bb3_add28_0_NO_SHIFT_REG > input_wii_sub29);
assign local_bb3_cmp1_i9_valid_out = local_bb3_cmp1_i9_inputs_ready;
assign local_bb3_cmp1_i9_stall_local = local_bb3_cmp1_i9_stall_in;
assign rnode_1to2_bb3_add28_0_stall_in_0_NO_SHIFT_REG = (|local_bb3_cmp1_i9_stall_local);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb3_var__u9_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb3_var__u9_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_169to170_bb3_var__u9_0_NO_SHIFT_REG;
 logic rnode_169to170_bb3_var__u9_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_169to170_bb3_var__u9_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb3_var__u9_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb3_var__u9_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb3_var__u9_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb3_var__u9_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb3_var__u9_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb3_var__u9_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb3_var__u9_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb3_var__u9_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb3_var__u9),
	.data_out(rnode_169to170_bb3_var__u9_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb3_var__u9_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb3_var__u9_0_reg_170_fifo.DATA_WIDTH = 64;
defparam rnode_169to170_bb3_var__u9_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb3_var__u9_0_reg_170_fifo.IMPL = "ll_reg";

assign rnode_169to170_bb3_var__u9_0_reg_170_inputs_ready_NO_SHIFT_REG = local_bb3_var__u9_valid_out;
assign local_bb3_var__u9_stall_in = rnode_169to170_bb3_var__u9_0_stall_out_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb3_var__u9_0_NO_SHIFT_REG = rnode_169to170_bb3_var__u9_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb3_var__u9_0_stall_in_reg_170_NO_SHIFT_REG = rnode_169to170_bb3_var__u9_0_stall_in_NO_SHIFT_REG;
assign rnode_169to170_bb3_var__u9_0_valid_out_NO_SHIFT_REG = rnode_169to170_bb3_var__u9_0_valid_out_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_indvars_iv_0_valid_out_NO_SHIFT_REG;
 logic rnode_396to397_indvars_iv_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_396to397_indvars_iv_0_NO_SHIFT_REG;
 logic rnode_396to397_indvars_iv_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_396to397_indvars_iv_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_indvars_iv_0_valid_out_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_indvars_iv_0_stall_in_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_indvars_iv_0_stall_out_reg_397_NO_SHIFT_REG;
wire [64:0] rci_rcnode_171to398_rc1_arrayidx43_0_reg_171;

acl_data_fifo rnode_396to397_indvars_iv_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_indvars_iv_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_indvars_iv_0_stall_in_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_indvars_iv_0_valid_out_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_indvars_iv_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(rnode_169to396_indvars_iv_0_NO_SHIFT_REG),
	.data_out(rnode_396to397_indvars_iv_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_indvars_iv_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_indvars_iv_0_reg_397_fifo.DATA_WIDTH = 64;
defparam rnode_396to397_indvars_iv_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_indvars_iv_0_reg_397_fifo.IMPL = "ll_reg";

assign rnode_396to397_indvars_iv_0_reg_397_inputs_ready_NO_SHIFT_REG = rnode_169to396_indvars_iv_0_valid_out_NO_SHIFT_REG;
assign rnode_169to396_indvars_iv_0_stall_in_NO_SHIFT_REG = rnode_396to397_indvars_iv_0_stall_out_reg_397_NO_SHIFT_REG;
assign rnode_396to397_indvars_iv_0_NO_SHIFT_REG = rnode_396to397_indvars_iv_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_indvars_iv_0_stall_in_reg_397_NO_SHIFT_REG = rnode_396to397_indvars_iv_0_stall_in_NO_SHIFT_REG;
assign rnode_396to397_indvars_iv_0_valid_out_NO_SHIFT_REG = rnode_396to397_indvars_iv_0_valid_out_reg_397_NO_SHIFT_REG;
assign rci_rcnode_171to398_rc1_arrayidx43_0_reg_171[63:0] = (rnode_170to171_arrayidx43_1_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign rci_rcnode_171to398_rc1_arrayidx43_0_reg_171[64] = rnode_170to171_var__u8_1_NO_SHIFT_REG;

// Register node:
//  * latency = 227
//  * capacity = 227
 logic rcnode_171to398_rc1_arrayidx43_0_valid_out_NO_SHIFT_REG;
 logic rcnode_171to398_rc1_arrayidx43_0_stall_in_NO_SHIFT_REG;
 logic [64:0] rcnode_171to398_rc1_arrayidx43_0_NO_SHIFT_REG;
 logic rcnode_171to398_rc1_arrayidx43_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [64:0] rcnode_171to398_rc1_arrayidx43_0_reg_398_NO_SHIFT_REG;
 logic rcnode_171to398_rc1_arrayidx43_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rcnode_171to398_rc1_arrayidx43_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rcnode_171to398_rc1_arrayidx43_0_stall_out_0_reg_398_IP_NO_SHIFT_REG;
 logic rcnode_171to398_rc1_arrayidx43_0_stall_out_0_reg_398_NO_SHIFT_REG;
wire [32:0] rci_rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_2;

acl_data_fifo rcnode_171to398_rc1_arrayidx43_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_171to398_rc1_arrayidx43_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_171to398_rc1_arrayidx43_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rcnode_171to398_rc1_arrayidx43_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rcnode_171to398_rc1_arrayidx43_0_stall_out_0_reg_398_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_171to398_rc1_arrayidx43_0_reg_171),
	.data_out(rcnode_171to398_rc1_arrayidx43_0_reg_398_NO_SHIFT_REG)
);

defparam rcnode_171to398_rc1_arrayidx43_0_reg_398_fifo.DEPTH = 228;
defparam rcnode_171to398_rc1_arrayidx43_0_reg_398_fifo.DATA_WIDTH = 65;
defparam rcnode_171to398_rc1_arrayidx43_0_reg_398_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_171to398_rc1_arrayidx43_0_reg_398_fifo.IMPL = "ram";

assign rcnode_171to398_rc1_arrayidx43_0_reg_398_inputs_ready_NO_SHIFT_REG = (rnode_170to171_arrayidx43_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_var__u8_0_valid_out_1_NO_SHIFT_REG);
assign rcnode_171to398_rc1_arrayidx43_0_stall_out_0_reg_398_NO_SHIFT_REG = (~(rcnode_171to398_rc1_arrayidx43_0_reg_398_inputs_ready_NO_SHIFT_REG) | rcnode_171to398_rc1_arrayidx43_0_stall_out_0_reg_398_IP_NO_SHIFT_REG);
assign rnode_170to171_arrayidx43_0_stall_in_1_NO_SHIFT_REG = rcnode_171to398_rc1_arrayidx43_0_stall_out_0_reg_398_NO_SHIFT_REG;
assign rnode_170to171_var__u8_0_stall_in_1_NO_SHIFT_REG = rcnode_171to398_rc1_arrayidx43_0_stall_out_0_reg_398_NO_SHIFT_REG;
assign rcnode_171to398_rc1_arrayidx43_0_NO_SHIFT_REG = rcnode_171to398_rc1_arrayidx43_0_reg_398_NO_SHIFT_REG;
assign rcnode_171to398_rc1_arrayidx43_0_stall_in_reg_398_NO_SHIFT_REG = rcnode_171to398_rc1_arrayidx43_0_stall_in_NO_SHIFT_REG;
assign rcnode_171to398_rc1_arrayidx43_0_valid_out_NO_SHIFT_REG = rcnode_171to398_rc1_arrayidx43_0_valid_out_reg_398_NO_SHIFT_REG;
assign rci_rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_2[0] = local_bb3_cmp1_i9;
assign rci_rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_2[32:1] = rnode_1to2_bb3_add28_1_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_2to3_rc0_bb3_cmp1_i9_0_valid_out_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_in_NO_SHIFT_REG;
 logic [32:0] rcnode_2to3_rc0_bb3_cmp1_i9_0_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [32:0] rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb3_cmp1_i9_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_out_0_reg_3_IP_NO_SHIFT_REG;
 logic rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_out_0_reg_3_NO_SHIFT_REG;

acl_data_fifo rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rcnode_2to3_rc0_bb3_cmp1_i9_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_out_0_reg_3_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_2),
	.data_out(rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_NO_SHIFT_REG)
);

defparam rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_fifo.DEPTH = 1;
defparam rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_fifo.DATA_WIDTH = 33;
defparam rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_fifo.IMPL = "ll_reg";

assign rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_inputs_ready_NO_SHIFT_REG = (local_bb3_cmp1_i9_valid_out & rnode_1to2_bb3_add28_0_valid_out_1_NO_SHIFT_REG);
assign rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_out_0_reg_3_NO_SHIFT_REG = (~(rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_inputs_ready_NO_SHIFT_REG) | rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_out_0_reg_3_IP_NO_SHIFT_REG);
assign local_bb3_cmp1_i9_stall_in = rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_out_0_reg_3_NO_SHIFT_REG;
assign rnode_1to2_bb3_add28_0_stall_in_1_NO_SHIFT_REG = rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_out_0_reg_3_NO_SHIFT_REG;
assign rcnode_2to3_rc0_bb3_cmp1_i9_0_NO_SHIFT_REG = rcnode_2to3_rc0_bb3_cmp1_i9_0_reg_3_NO_SHIFT_REG;
assign rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_in_reg_3_NO_SHIFT_REG = rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_in_NO_SHIFT_REG;
assign rcnode_2to3_rc0_bb3_cmp1_i9_0_valid_out_NO_SHIFT_REG = rcnode_2to3_rc0_bb3_cmp1_i9_0_valid_out_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_arrayidx46_valid_out;
wire local_bb3_arrayidx46_stall_in;
wire local_bb3_arrayidx46_inputs_ready;
wire local_bb3_arrayidx46_stall_local;
wire [63:0] local_bb3_arrayidx46;

assign local_bb3_arrayidx46_inputs_ready = rnode_169to170_bb3_var__u9_0_valid_out_NO_SHIFT_REG;
assign local_bb3_arrayidx46 = ((input_gaussian & 64'hFFFFFFFFFFFFFC00) + (rnode_169to170_bb3_var__u9_0_NO_SHIFT_REG << 6'h2));
assign local_bb3_arrayidx46_valid_out = local_bb3_arrayidx46_inputs_ready;
assign local_bb3_arrayidx46_stall_local = local_bb3_arrayidx46_stall_in;
assign rnode_169to170_bb3_var__u9_0_stall_in_NO_SHIFT_REG = (|local_bb3_arrayidx46_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb3_indvars_iv_next_stall_local;
wire [63:0] local_bb3_indvars_iv_next;
wire [353:0] rci_rcnode_398to399_rc0_idxprom_0_reg_398;

assign local_bb3_indvars_iv_next = (rnode_396to397_indvars_iv_0_NO_SHIFT_REG + 64'h1);
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[63:0] = (rcnode_1to398_rc9_idxprom_0_NO_SHIFT_REG[63:0] & 64'hFFFFFFFF);
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[64] = rcnode_1to398_rc9_idxprom_0_NO_SHIFT_REG[64];
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[128:65] = rcnode_1to398_rc9_idxprom_0_NO_SHIFT_REG[128:65];
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[160:129] = rcnode_1to398_rc9_idxprom_0_NO_SHIFT_REG[160:129];
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[192:161] = rcnode_1to398_rc10_input_global_id_1_0_NO_SHIFT_REG[31:0];
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[224:193] = rcnode_1to398_rc10_input_global_id_1_0_NO_SHIFT_REG[63:32];
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[256:225] = rnode_6to398_sub25_add24_0_NO_SHIFT_REG;
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[320:257] = (rcnode_171to398_rc1_arrayidx43_0_NO_SHIFT_REG[63:0] & 64'hFFFFFFFFFFFFFFFC);
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[352:321] = rnode_331to398_ld__0_NO_SHIFT_REG;
assign rci_rcnode_398to399_rc0_idxprom_0_reg_398[353] = rcnode_171to398_rc1_arrayidx43_0_NO_SHIFT_REG[64];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_398to399_rc0_idxprom_0_valid_out_0_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_stall_in_0_NO_SHIFT_REG;
 logic [353:0] rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_valid_out_1_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_stall_in_1_NO_SHIFT_REG;
 logic [353:0] rcnode_398to399_rc0_idxprom_1_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [353:0] rcnode_398to399_rc0_idxprom_0_reg_399_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_valid_out_0_reg_399_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_stall_in_0_reg_399_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_IP_NO_SHIFT_REG;
 logic rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_NO_SHIFT_REG;

acl_data_fifo rcnode_398to399_rc0_idxprom_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_398to399_rc0_idxprom_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_398to399_rc0_idxprom_0_stall_in_0_reg_399_NO_SHIFT_REG),
	.valid_out(rcnode_398to399_rc0_idxprom_0_valid_out_0_reg_399_NO_SHIFT_REG),
	.stall_out(rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_398to399_rc0_idxprom_0_reg_398),
	.data_out(rcnode_398to399_rc0_idxprom_0_reg_399_NO_SHIFT_REG)
);

defparam rcnode_398to399_rc0_idxprom_0_reg_399_fifo.DEPTH = 1;
defparam rcnode_398to399_rc0_idxprom_0_reg_399_fifo.DATA_WIDTH = 354;
defparam rcnode_398to399_rc0_idxprom_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_398to399_rc0_idxprom_0_reg_399_fifo.IMPL = "ll_reg";

assign rcnode_398to399_rc0_idxprom_0_reg_399_inputs_ready_NO_SHIFT_REG = (rnode_6to398_sub25_add24_0_valid_out_NO_SHIFT_REG & rnode_331to398_ld__0_valid_out_NO_SHIFT_REG & rcnode_1to398_rc9_idxprom_0_valid_out_NO_SHIFT_REG & rcnode_1to398_rc10_input_global_id_1_0_valid_out_NO_SHIFT_REG & rcnode_171to398_rc1_arrayidx43_0_valid_out_NO_SHIFT_REG);
assign rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_NO_SHIFT_REG = (~(rcnode_398to399_rc0_idxprom_0_reg_399_inputs_ready_NO_SHIFT_REG) | rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_IP_NO_SHIFT_REG);
assign rnode_6to398_sub25_add24_0_stall_in_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_NO_SHIFT_REG;
assign rnode_331to398_ld__0_stall_in_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_NO_SHIFT_REG;
assign rcnode_1to398_rc9_idxprom_0_stall_in_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_NO_SHIFT_REG;
assign rcnode_1to398_rc10_input_global_id_1_0_stall_in_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_NO_SHIFT_REG;
assign rcnode_171to398_rc1_arrayidx43_0_stall_in_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_stall_out_0_reg_399_NO_SHIFT_REG;
assign rcnode_398to399_rc0_idxprom_0_stall_in_0_reg_399_NO_SHIFT_REG = (rcnode_398to399_rc0_idxprom_0_stall_in_0_NO_SHIFT_REG | rcnode_398to399_rc0_idxprom_0_stall_in_1_NO_SHIFT_REG);
assign rcnode_398to399_rc0_idxprom_0_valid_out_0_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_valid_out_0_reg_399_NO_SHIFT_REG;
assign rcnode_398to399_rc0_idxprom_0_valid_out_1_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_valid_out_0_reg_399_NO_SHIFT_REG;
assign rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_reg_399_NO_SHIFT_REG;
assign rcnode_398to399_rc0_idxprom_1_NO_SHIFT_REG = rcnode_398to399_rc0_idxprom_0_reg_399_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_sub29_add28_valid_out;
wire local_bb3_sub29_add28_stall_in;
wire local_bb3_sub29_add28_inputs_ready;
wire local_bb3_sub29_add28_stall_local;
wire [31:0] local_bb3_sub29_add28;

assign local_bb3_sub29_add28_inputs_ready = rcnode_2to3_rc0_bb3_cmp1_i9_0_valid_out_NO_SHIFT_REG;
assign local_bb3_sub29_add28 = (rcnode_2to3_rc0_bb3_cmp1_i9_0_NO_SHIFT_REG[0] ? input_wii_sub29 : rcnode_2to3_rc0_bb3_cmp1_i9_0_NO_SHIFT_REG[32:1]);
assign local_bb3_sub29_add28_valid_out = local_bb3_sub29_add28_inputs_ready;
assign local_bb3_sub29_add28_stall_local = local_bb3_sub29_add28_stall_in;
assign rcnode_2to3_rc0_bb3_cmp1_i9_0_stall_in_NO_SHIFT_REG = (|local_bb3_sub29_add28_stall_local);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb3_arrayidx46_0_valid_out_NO_SHIFT_REG;
 logic rnode_170to171_bb3_arrayidx46_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_170to171_bb3_arrayidx46_0_NO_SHIFT_REG;
 logic rnode_170to171_bb3_arrayidx46_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_170to171_bb3_arrayidx46_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb3_arrayidx46_0_valid_out_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb3_arrayidx46_0_stall_in_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb3_arrayidx46_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb3_arrayidx46_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb3_arrayidx46_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb3_arrayidx46_0_stall_in_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb3_arrayidx46_0_valid_out_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb3_arrayidx46_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in((local_bb3_arrayidx46 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_170to171_bb3_arrayidx46_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb3_arrayidx46_0_reg_171_fifo.DEPTH = 2;
defparam rnode_170to171_bb3_arrayidx46_0_reg_171_fifo.DATA_WIDTH = 64;
defparam rnode_170to171_bb3_arrayidx46_0_reg_171_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_170to171_bb3_arrayidx46_0_reg_171_fifo.IMPL = "ll_reg";

assign rnode_170to171_bb3_arrayidx46_0_reg_171_inputs_ready_NO_SHIFT_REG = local_bb3_arrayidx46_valid_out;
assign local_bb3_arrayidx46_stall_in = rnode_170to171_bb3_arrayidx46_0_stall_out_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb3_arrayidx46_0_NO_SHIFT_REG = rnode_170to171_bb3_arrayidx46_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb3_arrayidx46_0_stall_in_reg_171_NO_SHIFT_REG = rnode_170to171_bb3_arrayidx46_0_stall_in_NO_SHIFT_REG;
assign rnode_170to171_bb3_arrayidx46_0_valid_out_NO_SHIFT_REG = rnode_170to171_bb3_arrayidx46_0_valid_out_reg_171_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_indvars_iv_next_valid_out_1;
wire local_bb3_indvars_iv_next_stall_in_1;
wire local_bb3_var__u10_valid_out;
wire local_bb3_var__u10_stall_in;
wire local_bb3_var__u10_inputs_ready;
wire local_bb3_var__u10_stall_local;
wire [31:0] local_bb3_var__u10;
 reg local_bb3_indvars_iv_next_consumed_1_NO_SHIFT_REG;
 reg local_bb3_var__u10_consumed_0_NO_SHIFT_REG;

assign local_bb3_var__u10_inputs_ready = rnode_396to397_indvars_iv_0_valid_out_NO_SHIFT_REG;
assign local_bb3_var__u10 = local_bb3_indvars_iv_next[31:0];
assign local_bb3_var__u10_stall_local = ((local_bb3_indvars_iv_next_stall_in_1 & ~(local_bb3_indvars_iv_next_consumed_1_NO_SHIFT_REG)) | (local_bb3_var__u10_stall_in & ~(local_bb3_var__u10_consumed_0_NO_SHIFT_REG)));
assign local_bb3_indvars_iv_next_valid_out_1 = (local_bb3_var__u10_inputs_ready & ~(local_bb3_indvars_iv_next_consumed_1_NO_SHIFT_REG));
assign local_bb3_var__u10_valid_out = (local_bb3_var__u10_inputs_ready & ~(local_bb3_var__u10_consumed_0_NO_SHIFT_REG));
assign rnode_396to397_indvars_iv_0_stall_in_NO_SHIFT_REG = (|local_bb3_var__u10_stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_indvars_iv_next_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_var__u10_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb3_indvars_iv_next_consumed_1_NO_SHIFT_REG <= (local_bb3_var__u10_inputs_ready & (local_bb3_indvars_iv_next_consumed_1_NO_SHIFT_REG | ~(local_bb3_indvars_iv_next_stall_in_1)) & local_bb3_var__u10_stall_local);
		local_bb3_var__u10_consumed_0_NO_SHIFT_REG <= (local_bb3_var__u10_inputs_ready & (local_bb3_var__u10_consumed_0_NO_SHIFT_REG | ~(local_bb3_var__u10_stall_in)) & local_bb3_var__u10_stall_local);
	end
end


// This section implements a registered operation.
// 
wire local_bb3_mul32_inputs_ready;
 reg local_bb3_mul32_valid_out_NO_SHIFT_REG;
wire local_bb3_mul32_stall_in;
wire local_bb3_mul32_output_regs_ready;
wire [31:0] local_bb3_mul32;
 reg local_bb3_mul32_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_mul32_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_mul32_causedstall;

acl_int_mult int_module_local_bb3_mul32 (
	.clock(clock),
	.dataa(local_bb3_sub29_add28),
	.datab(input_global_size_0),
	.enable(local_bb3_mul32_output_regs_ready),
	.result(local_bb3_mul32)
);

defparam int_module_local_bb3_mul32.INPUT1_WIDTH = 32;
defparam int_module_local_bb3_mul32.INPUT2_WIDTH = 32;
defparam int_module_local_bb3_mul32.OUTPUT_WIDTH = 32;
defparam int_module_local_bb3_mul32.LATENCY = 3;
defparam int_module_local_bb3_mul32.SIGNED = 0;

assign local_bb3_mul32_inputs_ready = local_bb3_sub29_add28_valid_out;
assign local_bb3_mul32_output_regs_ready = (&(~(local_bb3_mul32_valid_out_NO_SHIFT_REG) | ~(local_bb3_mul32_stall_in)));
assign local_bb3_sub29_add28_stall_in = (~(local_bb3_mul32_output_regs_ready) | ~(local_bb3_mul32_inputs_ready));
assign local_bb3_mul32_causedstall = (local_bb3_mul32_inputs_ready && (~(local_bb3_mul32_output_regs_ready) && !(~(local_bb3_mul32_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul32_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul32_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul32_output_regs_ready)
		begin
			local_bb3_mul32_valid_pipe_0_NO_SHIFT_REG <= local_bb3_mul32_inputs_ready;
			local_bb3_mul32_valid_pipe_1_NO_SHIFT_REG <= local_bb3_mul32_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul32_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul32_output_regs_ready)
		begin
			local_bb3_mul32_valid_out_NO_SHIFT_REG <= local_bb3_mul32_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb3_mul32_stall_in))
			begin
				local_bb3_mul32_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_397to399_bb3_indvars_iv_next_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to399_bb3_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_397to399_bb3_indvars_iv_next_0_NO_SHIFT_REG;
 logic rnode_397to399_bb3_indvars_iv_next_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_397to399_bb3_indvars_iv_next_0_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb3_indvars_iv_next_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb3_indvars_iv_next_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb3_indvars_iv_next_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_397to399_bb3_indvars_iv_next_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to399_bb3_indvars_iv_next_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to399_bb3_indvars_iv_next_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_397to399_bb3_indvars_iv_next_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_397to399_bb3_indvars_iv_next_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in(local_bb3_indvars_iv_next),
	.data_out(rnode_397to399_bb3_indvars_iv_next_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_397to399_bb3_indvars_iv_next_0_reg_399_fifo.DEPTH = 3;
defparam rnode_397to399_bb3_indvars_iv_next_0_reg_399_fifo.DATA_WIDTH = 64;
defparam rnode_397to399_bb3_indvars_iv_next_0_reg_399_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_397to399_bb3_indvars_iv_next_0_reg_399_fifo.IMPL = "ll_reg";

assign rnode_397to399_bb3_indvars_iv_next_0_reg_399_inputs_ready_NO_SHIFT_REG = local_bb3_indvars_iv_next_valid_out_1;
assign local_bb3_indvars_iv_next_stall_in_1 = rnode_397to399_bb3_indvars_iv_next_0_stall_out_reg_399_NO_SHIFT_REG;
assign rnode_397to399_bb3_indvars_iv_next_0_NO_SHIFT_REG = rnode_397to399_bb3_indvars_iv_next_0_reg_399_NO_SHIFT_REG;
assign rnode_397to399_bb3_indvars_iv_next_0_stall_in_reg_399_NO_SHIFT_REG = rnode_397to399_bb3_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
assign rnode_397to399_bb3_indvars_iv_next_0_valid_out_NO_SHIFT_REG = rnode_397to399_bb3_indvars_iv_next_0_valid_out_reg_399_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_397to398_bb3_var__u10_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to398_bb3_var__u10_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb3_var__u10_0_NO_SHIFT_REG;
 logic rnode_397to398_bb3_var__u10_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb3_var__u10_0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb3_var__u10_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb3_var__u10_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb3_var__u10_0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_397to398_bb3_var__u10_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to398_bb3_var__u10_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to398_bb3_var__u10_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_397to398_bb3_var__u10_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_397to398_bb3_var__u10_0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(local_bb3_var__u10),
	.data_out(rnode_397to398_bb3_var__u10_0_reg_398_NO_SHIFT_REG)
);

defparam rnode_397to398_bb3_var__u10_0_reg_398_fifo.DEPTH = 1;
defparam rnode_397to398_bb3_var__u10_0_reg_398_fifo.DATA_WIDTH = 32;
defparam rnode_397to398_bb3_var__u10_0_reg_398_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to398_bb3_var__u10_0_reg_398_fifo.IMPL = "ll_reg";

assign rnode_397to398_bb3_var__u10_0_reg_398_inputs_ready_NO_SHIFT_REG = local_bb3_var__u10_valid_out;
assign local_bb3_var__u10_stall_in = rnode_397to398_bb3_var__u10_0_stall_out_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb3_var__u10_0_NO_SHIFT_REG = rnode_397to398_bb3_var__u10_0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb3_var__u10_0_stall_in_reg_398_NO_SHIFT_REG = rnode_397to398_bb3_var__u10_0_stall_in_NO_SHIFT_REG;
assign rnode_397to398_bb3_var__u10_0_valid_out_NO_SHIFT_REG = rnode_397to398_bb3_var__u10_0_valid_out_reg_398_NO_SHIFT_REG;

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_6to6_bb3_mul32_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to6_bb3_mul32_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_6to6_bb3_mul32_0_NO_SHIFT_REG;
 logic rnode_6to6_bb3_mul32_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_6to6_bb3_mul32_0_reg_6_NO_SHIFT_REG;
 logic rnode_6to6_bb3_mul32_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_6to6_bb3_mul32_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_6to6_bb3_mul32_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_6to6_bb3_mul32_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to6_bb3_mul32_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to6_bb3_mul32_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_6to6_bb3_mul32_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_6to6_bb3_mul32_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_mul32),
	.data_out(rnode_6to6_bb3_mul32_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_6to6_bb3_mul32_0_reg_6_fifo.DEPTH = 3;
defparam rnode_6to6_bb3_mul32_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_6to6_bb3_mul32_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_6to6_bb3_mul32_0_reg_6_fifo.IMPL = "zl_reg";

assign rnode_6to6_bb3_mul32_0_reg_6_inputs_ready_NO_SHIFT_REG = local_bb3_mul32_valid_out_NO_SHIFT_REG;
assign local_bb3_mul32_stall_in = rnode_6to6_bb3_mul32_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_6to6_bb3_mul32_0_NO_SHIFT_REG = rnode_6to6_bb3_mul32_0_reg_6_NO_SHIFT_REG;
assign rnode_6to6_bb3_mul32_0_stall_in_reg_6_NO_SHIFT_REG = rnode_6to6_bb3_mul32_0_stall_in_NO_SHIFT_REG;
assign rnode_6to6_bb3_mul32_0_valid_out_NO_SHIFT_REG = rnode_6to6_bb3_mul32_0_valid_out_reg_6_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp20_valid_out;
wire local_bb3_cmp20_stall_in;
wire local_bb3_cmp20_inputs_ready;
wire local_bb3_cmp20_stall_local;
wire local_bb3_cmp20;

assign local_bb3_cmp20_inputs_ready = rnode_397to398_bb3_var__u10_0_valid_out_NO_SHIFT_REG;
assign local_bb3_cmp20 = ($signed(rnode_397to398_bb3_var__u10_0_NO_SHIFT_REG) > $signed(input_r));
assign local_bb3_cmp20_valid_out = local_bb3_cmp20_inputs_ready;
assign local_bb3_cmp20_stall_local = local_bb3_cmp20_stall_in;
assign rnode_397to398_bb3_var__u10_0_stall_in_NO_SHIFT_REG = (|local_bb3_cmp20_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb3_add33_valid_out;
wire local_bb3_add33_stall_in;
wire local_bb3_add33_inputs_ready;
wire local_bb3_add33_stall_local;
wire [31:0] local_bb3_add33;

assign local_bb3_add33_inputs_ready = (rnode_1to6_sub25_add24_0_valid_out_0_NO_SHIFT_REG & rnode_6to6_bb3_mul32_0_valid_out_NO_SHIFT_REG);
assign local_bb3_add33 = (rnode_6to6_bb3_mul32_0_NO_SHIFT_REG + rnode_1to6_sub25_add24_0_NO_SHIFT_REG);
assign local_bb3_add33_valid_out = local_bb3_add33_inputs_ready;
assign local_bb3_add33_stall_local = local_bb3_add33_stall_in;
assign rnode_1to6_sub25_add24_0_stall_in_0_NO_SHIFT_REG = (local_bb3_add33_stall_local | ~(local_bb3_add33_inputs_ready));
assign rnode_6to6_bb3_mul32_0_stall_in_NO_SHIFT_REG = (local_bb3_add33_stall_local | ~(local_bb3_add33_inputs_ready));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_398to399_bb3_cmp20_0_valid_out_NO_SHIFT_REG;
 logic rnode_398to399_bb3_cmp20_0_stall_in_NO_SHIFT_REG;
 logic rnode_398to399_bb3_cmp20_0_NO_SHIFT_REG;
 logic rnode_398to399_bb3_cmp20_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic rnode_398to399_bb3_cmp20_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb3_cmp20_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb3_cmp20_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb3_cmp20_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_398to399_bb3_cmp20_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to399_bb3_cmp20_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to399_bb3_cmp20_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_398to399_bb3_cmp20_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_398to399_bb3_cmp20_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in(local_bb3_cmp20),
	.data_out(rnode_398to399_bb3_cmp20_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_398to399_bb3_cmp20_0_reg_399_fifo.DEPTH = 1;
defparam rnode_398to399_bb3_cmp20_0_reg_399_fifo.DATA_WIDTH = 1;
defparam rnode_398to399_bb3_cmp20_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to399_bb3_cmp20_0_reg_399_fifo.IMPL = "ll_reg";

assign rnode_398to399_bb3_cmp20_0_reg_399_inputs_ready_NO_SHIFT_REG = local_bb3_cmp20_valid_out;
assign local_bb3_cmp20_stall_in = rnode_398to399_bb3_cmp20_0_stall_out_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb3_cmp20_0_NO_SHIFT_REG = rnode_398to399_bb3_cmp20_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb3_cmp20_0_stall_in_reg_399_NO_SHIFT_REG = rnode_398to399_bb3_cmp20_0_stall_in_NO_SHIFT_REG;
assign rnode_398to399_bb3_cmp20_0_valid_out_NO_SHIFT_REG = rnode_398to399_bb3_cmp20_0_valid_out_reg_399_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb3_add33_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb3_add33_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb3_add33_0_NO_SHIFT_REG;
 logic rnode_6to7_bb3_add33_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb3_add33_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb3_add33_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb3_add33_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb3_add33_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb3_add33_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb3_add33_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb3_add33_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb3_add33_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb3_add33_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb3_add33),
	.data_out(rnode_6to7_bb3_add33_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb3_add33_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb3_add33_0_reg_7_fifo.DATA_WIDTH = 32;
defparam rnode_6to7_bb3_add33_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb3_add33_0_reg_7_fifo.IMPL = "ll_reg";

assign rnode_6to7_bb3_add33_0_reg_7_inputs_ready_NO_SHIFT_REG = local_bb3_add33_valid_out;
assign local_bb3_add33_stall_in = rnode_6to7_bb3_add33_0_stall_out_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb3_add33_0_NO_SHIFT_REG = rnode_6to7_bb3_add33_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb3_add33_0_stall_in_reg_7_NO_SHIFT_REG = rnode_6to7_bb3_add33_0_stall_in_NO_SHIFT_REG;
assign rnode_6to7_bb3_add33_0_valid_out_NO_SHIFT_REG = rnode_6to7_bb3_add33_0_valid_out_reg_7_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u11_valid_out;
wire local_bb3_var__u11_stall_in;
wire local_bb3_var__u11_inputs_ready;
wire local_bb3_var__u11_stall_local;
wire local_bb3_var__u11;

assign local_bb3_var__u11_inputs_ready = (rnode_398to399_bb3_cmp20_0_valid_out_NO_SHIFT_REG & rcnode_398to399_rc0_idxprom_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_var__u11 = (rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[353] | rnode_398to399_bb3_cmp20_0_NO_SHIFT_REG);
assign local_bb3_var__u11_valid_out = local_bb3_var__u11_inputs_ready;
assign local_bb3_var__u11_stall_local = local_bb3_var__u11_stall_in;
assign rnode_398to399_bb3_cmp20_0_stall_in_NO_SHIFT_REG = (local_bb3_var__u11_stall_local | ~(local_bb3_var__u11_inputs_ready));
assign rcnode_398to399_rc0_idxprom_0_stall_in_1_NO_SHIFT_REG = (local_bb3_var__u11_stall_local | ~(local_bb3_var__u11_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb3_idxprom34_stall_local;
wire [63:0] local_bb3_idxprom34;

assign local_bb3_idxprom34[63:32] = 32'h0;
assign local_bb3_idxprom34[31:0] = rnode_6to7_bb3_add33_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_arrayidx35_valid_out;
wire local_bb3_arrayidx35_stall_in;
wire local_bb3_arrayidx35_inputs_ready;
wire local_bb3_arrayidx35_stall_local;
wire [63:0] local_bb3_arrayidx35;

assign local_bb3_arrayidx35_inputs_ready = rnode_6to7_bb3_add33_0_valid_out_NO_SHIFT_REG;
assign local_bb3_arrayidx35 = ((input_in & 64'hFFFFFFFFFFFFFC00) + ((local_bb3_idxprom34 & 64'hFFFFFFFF) << 6'h2));
assign local_bb3_arrayidx35_valid_out = local_bb3_arrayidx35_inputs_ready;
assign local_bb3_arrayidx35_stall_local = local_bb3_arrayidx35_stall_in;
assign rnode_6to7_bb3_add33_0_stall_in_NO_SHIFT_REG = (|local_bb3_arrayidx35_stall_local);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb3_arrayidx35_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb3_arrayidx35_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_7to8_bb3_arrayidx35_0_NO_SHIFT_REG;
 logic rnode_7to8_bb3_arrayidx35_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_7to8_bb3_arrayidx35_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb3_arrayidx35_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb3_arrayidx35_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb3_arrayidx35_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb3_arrayidx35_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb3_arrayidx35_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb3_arrayidx35_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb3_arrayidx35_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb3_arrayidx35_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in((local_bb3_arrayidx35 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_7to8_bb3_arrayidx35_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb3_arrayidx35_0_reg_8_fifo.DEPTH = 2;
defparam rnode_7to8_bb3_arrayidx35_0_reg_8_fifo.DATA_WIDTH = 64;
defparam rnode_7to8_bb3_arrayidx35_0_reg_8_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_7to8_bb3_arrayidx35_0_reg_8_fifo.IMPL = "ll_reg";

assign rnode_7to8_bb3_arrayidx35_0_reg_8_inputs_ready_NO_SHIFT_REG = local_bb3_arrayidx35_valid_out;
assign local_bb3_arrayidx35_stall_in = rnode_7to8_bb3_arrayidx35_0_stall_out_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb3_arrayidx35_0_NO_SHIFT_REG = rnode_7to8_bb3_arrayidx35_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb3_arrayidx35_0_stall_in_reg_8_NO_SHIFT_REG = rnode_7to8_bb3_arrayidx35_0_stall_in_NO_SHIFT_REG;
assign rnode_7to8_bb3_arrayidx35_0_valid_out_NO_SHIFT_REG = rnode_7to8_bb3_arrayidx35_0_valid_out_reg_8_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb3_ld__inputs_ready;
 reg local_bb3_ld__valid_out_NO_SHIFT_REG;
wire local_bb3_ld__stall_in;
wire local_bb3_ld__output_regs_ready;
wire local_bb3_ld__fu_stall_out;
wire local_bb3_ld__fu_valid_out;
wire [31:0] local_bb3_ld__lsu_dataout;
 reg [31:0] local_bb3_ld__NO_SHIFT_REG;
wire local_bb3_ld__causedstall;

lsu_top lsu_local_bb3_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb3_ld__fu_stall_out),
	.i_valid(local_bb3_ld__inputs_ready),
	.i_address((rnode_7to8_bb3_arrayidx35_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rnode_1to8_var__u8_0_NO_SHIFT_REG),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb3_ld__output_regs_ready)),
	.o_valid(local_bb3_ld__fu_valid_out),
	.o_readdata(local_bb3_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb3_ld__active),
	.avm_address(avm_local_bb3_ld__address),
	.avm_read(avm_local_bb3_ld__read),
	.avm_readdata(avm_local_bb3_ld__readdata),
	.avm_write(avm_local_bb3_ld__write),
	.avm_writeack(avm_local_bb3_ld__writeack),
	.avm_burstcount(avm_local_bb3_ld__burstcount),
	.avm_writedata(avm_local_bb3_ld__writedata),
	.avm_byteenable(avm_local_bb3_ld__byteenable),
	.avm_waitrequest(avm_local_bb3_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb3_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb3_ld_.AWIDTH = 33;
defparam lsu_local_bb3_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb3_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb3_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb3_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb3_ld_.READ = 1;
defparam lsu_local_bb3_ld_.ATOMIC = 0;
defparam lsu_local_bb3_ld_.WIDTH = 32;
defparam lsu_local_bb3_ld_.MWIDTH = 512;
defparam lsu_local_bb3_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb3_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb3_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb3_ld_.MEMORY_SIDE_MEM_LATENCY = 132;
defparam lsu_local_bb3_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb3_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb3_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb3_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb3_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb3_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb3_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb3_ld_.USECACHING = 1;
defparam lsu_local_bb3_ld_.CACHESIZE = 1024;
defparam lsu_local_bb3_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb3_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb3_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb3_ld_.ADDRSPACE = 1;
defparam lsu_local_bb3_ld_.STYLE = "BURST-COALESCED";

assign local_bb3_ld__inputs_ready = (rnode_7to8_bb3_arrayidx35_0_valid_out_NO_SHIFT_REG & rnode_1to8_var__u8_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3_ld__output_regs_ready = (&(~(local_bb3_ld__valid_out_NO_SHIFT_REG) | ~(local_bb3_ld__stall_in)));
assign rnode_7to8_bb3_arrayidx35_0_stall_in_NO_SHIFT_REG = (local_bb3_ld__fu_stall_out | ~(local_bb3_ld__inputs_ready));
assign rnode_1to8_var__u8_0_stall_in_0_NO_SHIFT_REG = (local_bb3_ld__fu_stall_out | ~(local_bb3_ld__inputs_ready));
assign local_bb3_ld__causedstall = (local_bb3_ld__inputs_ready && (local_bb3_ld__fu_stall_out && !(~(local_bb3_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_ld__NO_SHIFT_REG <= 'x;
		local_bb3_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_ld__output_regs_ready)
		begin
			local_bb3_ld__NO_SHIFT_REG <= local_bb3_ld__lsu_dataout;
			local_bb3_ld__valid_out_NO_SHIFT_REG <= local_bb3_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_ld__stall_in))
			begin
				local_bb3_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_168to168_bb3_ld__valid_out_0;
wire rstag_168to168_bb3_ld__stall_in_0;
wire rstag_168to168_bb3_ld__valid_out_1;
wire rstag_168to168_bb3_ld__stall_in_1;
wire rstag_168to168_bb3_ld__inputs_ready;
wire rstag_168to168_bb3_ld__stall_local;
 reg rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG;
wire rstag_168to168_bb3_ld__combined_valid;
 reg [31:0] rstag_168to168_bb3_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_168to168_bb3_ld_;
 reg rstag_168to168_bb3_ld__consumed_0_NO_SHIFT_REG;
 reg rstag_168to168_bb3_ld__consumed_1_NO_SHIFT_REG;

assign rstag_168to168_bb3_ld__inputs_ready = local_bb3_ld__valid_out_NO_SHIFT_REG;
assign rstag_168to168_bb3_ld_ = (rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG ? rstag_168to168_bb3_ld__staging_reg_NO_SHIFT_REG : local_bb3_ld__NO_SHIFT_REG);
assign rstag_168to168_bb3_ld__combined_valid = (rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG | rstag_168to168_bb3_ld__inputs_ready);
assign rstag_168to168_bb3_ld__stall_local = ((rstag_168to168_bb3_ld__stall_in_0 & ~(rstag_168to168_bb3_ld__consumed_0_NO_SHIFT_REG)) | (rstag_168to168_bb3_ld__stall_in_1 & ~(rstag_168to168_bb3_ld__consumed_1_NO_SHIFT_REG)));
assign rstag_168to168_bb3_ld__valid_out_0 = (rstag_168to168_bb3_ld__combined_valid & ~(rstag_168to168_bb3_ld__consumed_0_NO_SHIFT_REG));
assign rstag_168to168_bb3_ld__valid_out_1 = (rstag_168to168_bb3_ld__combined_valid & ~(rstag_168to168_bb3_ld__consumed_1_NO_SHIFT_REG));
assign local_bb3_ld__stall_in = (|rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_168to168_bb3_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_168to168_bb3_ld__stall_local)
		begin
			if (~(rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG <= rstag_168to168_bb3_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_168to168_bb3_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_168to168_bb3_ld__staging_reg_NO_SHIFT_REG <= local_bb3_ld__NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_168to168_bb3_ld__consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_168to168_bb3_ld__consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_168to168_bb3_ld__consumed_0_NO_SHIFT_REG <= (rstag_168to168_bb3_ld__combined_valid & (rstag_168to168_bb3_ld__consumed_0_NO_SHIFT_REG | ~(rstag_168to168_bb3_ld__stall_in_0)) & rstag_168to168_bb3_ld__stall_local);
		rstag_168to168_bb3_ld__consumed_1_NO_SHIFT_REG <= (rstag_168to168_bb3_ld__combined_valid & (rstag_168to168_bb3_ld__consumed_1_NO_SHIFT_REG | ~(rstag_168to168_bb3_ld__stall_in_1)) & rstag_168to168_bb3_ld__stall_local);
	end
end


// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_168to330_bb3_ld__0_valid_out_NO_SHIFT_REG;
 logic rnode_168to330_bb3_ld__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_168to330_bb3_ld__0_NO_SHIFT_REG;
 logic rnode_168to330_bb3_ld__0_reg_330_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to330_bb3_ld__0_reg_330_NO_SHIFT_REG;
 logic rnode_168to330_bb3_ld__0_valid_out_reg_330_NO_SHIFT_REG;
 logic rnode_168to330_bb3_ld__0_stall_in_reg_330_NO_SHIFT_REG;
 logic rnode_168to330_bb3_ld__0_stall_out_reg_330_NO_SHIFT_REG;

acl_data_fifo rnode_168to330_bb3_ld__0_reg_330_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to330_bb3_ld__0_reg_330_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to330_bb3_ld__0_stall_in_reg_330_NO_SHIFT_REG),
	.valid_out(rnode_168to330_bb3_ld__0_valid_out_reg_330_NO_SHIFT_REG),
	.stall_out(rnode_168to330_bb3_ld__0_stall_out_reg_330_NO_SHIFT_REG),
	.data_in(rstag_168to168_bb3_ld_),
	.data_out(rnode_168to330_bb3_ld__0_reg_330_NO_SHIFT_REG)
);

defparam rnode_168to330_bb3_ld__0_reg_330_fifo.DEPTH = 163;
defparam rnode_168to330_bb3_ld__0_reg_330_fifo.DATA_WIDTH = 32;
defparam rnode_168to330_bb3_ld__0_reg_330_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_168to330_bb3_ld__0_reg_330_fifo.IMPL = "ram";

assign rnode_168to330_bb3_ld__0_reg_330_inputs_ready_NO_SHIFT_REG = rstag_168to168_bb3_ld__valid_out_0;
assign rstag_168to168_bb3_ld__stall_in_0 = rnode_168to330_bb3_ld__0_stall_out_reg_330_NO_SHIFT_REG;
assign rnode_168to330_bb3_ld__0_NO_SHIFT_REG = rnode_168to330_bb3_ld__0_reg_330_NO_SHIFT_REG;
assign rnode_168to330_bb3_ld__0_stall_in_reg_330_NO_SHIFT_REG = rnode_168to330_bb3_ld__0_stall_in_NO_SHIFT_REG;
assign rnode_168to330_bb3_ld__0_valid_out_NO_SHIFT_REG = rnode_168to330_bb3_ld__0_valid_out_reg_330_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb3_cmp36_inputs_ready;
 reg local_bb3_cmp36_valid_out_NO_SHIFT_REG;
wire local_bb3_cmp36_stall_in;
wire local_bb3_cmp36_output_regs_ready;
wire local_bb3_cmp36;
 reg local_bb3_cmp36_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_cmp36_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_cmp36_causedstall;

acl_fp_cmp fp_module_local_bb3_cmp36 (
	.clock(clock),
	.dataa(rstag_168to168_bb3_ld_),
	.datab(32'h0),
	.enable(local_bb3_cmp36_output_regs_ready),
	.result(local_bb3_cmp36)
);

defparam fp_module_local_bb3_cmp36.COMPARISON_MODE = 3;

assign local_bb3_cmp36_inputs_ready = rstag_168to168_bb3_ld__valid_out_1;
assign local_bb3_cmp36_output_regs_ready = (&(~(local_bb3_cmp36_valid_out_NO_SHIFT_REG) | ~(local_bb3_cmp36_stall_in)));
assign rstag_168to168_bb3_ld__stall_in_1 = (~(local_bb3_cmp36_output_regs_ready) | ~(local_bb3_cmp36_inputs_ready));
assign local_bb3_cmp36_causedstall = (local_bb3_cmp36_inputs_ready && (~(local_bb3_cmp36_output_regs_ready) && !(~(local_bb3_cmp36_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_cmp36_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_cmp36_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_cmp36_output_regs_ready)
		begin
			local_bb3_cmp36_valid_pipe_0_NO_SHIFT_REG <= local_bb3_cmp36_inputs_ready;
			local_bb3_cmp36_valid_pipe_1_NO_SHIFT_REG <= local_bb3_cmp36_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_cmp36_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_cmp36_output_regs_ready)
		begin
			local_bb3_cmp36_valid_out_NO_SHIFT_REG <= local_bb3_cmp36_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb3_cmp36_stall_in))
			begin
				local_bb3_cmp36_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_171to171_bb3_cmp36_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_1_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_reg_171_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_171to171_bb3_cmp36_0_stall_out_reg_171_NO_SHIFT_REG;
 reg rnode_171to171_bb3_cmp36_0_consumed_0_NO_SHIFT_REG;
 reg rnode_171to171_bb3_cmp36_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_171to171_bb3_cmp36_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to171_bb3_cmp36_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to171_bb3_cmp36_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_171to171_bb3_cmp36_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_171to171_bb3_cmp36_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb3_cmp36),
	.data_out(rnode_171to171_bb3_cmp36_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_171to171_bb3_cmp36_0_reg_171_fifo.DEPTH = 3;
defparam rnode_171to171_bb3_cmp36_0_reg_171_fifo.DATA_WIDTH = 1;
defparam rnode_171to171_bb3_cmp36_0_reg_171_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_171to171_bb3_cmp36_0_reg_171_fifo.IMPL = "zl_reg";

assign rnode_171to171_bb3_cmp36_0_reg_171_inputs_ready_NO_SHIFT_REG = local_bb3_cmp36_valid_out_NO_SHIFT_REG;
assign local_bb3_cmp36_stall_in = rnode_171to171_bb3_cmp36_0_stall_out_reg_171_NO_SHIFT_REG;
assign rnode_171to171_bb3_cmp36_0_stall_in_0_reg_171_NO_SHIFT_REG = ((rnode_171to171_bb3_cmp36_0_stall_in_0_NO_SHIFT_REG & ~(rnode_171to171_bb3_cmp36_0_consumed_0_NO_SHIFT_REG)) | (rnode_171to171_bb3_cmp36_0_stall_in_1_NO_SHIFT_REG & ~(rnode_171to171_bb3_cmp36_0_consumed_1_NO_SHIFT_REG)));
assign rnode_171to171_bb3_cmp36_0_valid_out_0_NO_SHIFT_REG = (rnode_171to171_bb3_cmp36_0_valid_out_0_reg_171_NO_SHIFT_REG & ~(rnode_171to171_bb3_cmp36_0_consumed_0_NO_SHIFT_REG));
assign rnode_171to171_bb3_cmp36_0_valid_out_1_NO_SHIFT_REG = (rnode_171to171_bb3_cmp36_0_valid_out_0_reg_171_NO_SHIFT_REG & ~(rnode_171to171_bb3_cmp36_0_consumed_1_NO_SHIFT_REG));
assign rnode_171to171_bb3_cmp36_0_NO_SHIFT_REG = rnode_171to171_bb3_cmp36_0_reg_171_NO_SHIFT_REG;
assign rnode_171to171_bb3_cmp36_1_NO_SHIFT_REG = rnode_171to171_bb3_cmp36_0_reg_171_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_171to171_bb3_cmp36_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_171to171_bb3_cmp36_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_171to171_bb3_cmp36_0_consumed_0_NO_SHIFT_REG <= (rnode_171to171_bb3_cmp36_0_valid_out_0_reg_171_NO_SHIFT_REG & (rnode_171to171_bb3_cmp36_0_consumed_0_NO_SHIFT_REG | ~(rnode_171to171_bb3_cmp36_0_stall_in_0_NO_SHIFT_REG)) & rnode_171to171_bb3_cmp36_0_stall_in_0_reg_171_NO_SHIFT_REG);
		rnode_171to171_bb3_cmp36_0_consumed_1_NO_SHIFT_REG <= (rnode_171to171_bb3_cmp36_0_valid_out_0_reg_171_NO_SHIFT_REG & (rnode_171to171_bb3_cmp36_0_consumed_1_NO_SHIFT_REG | ~(rnode_171to171_bb3_cmp36_0_stall_in_1_NO_SHIFT_REG)) & rnode_171to171_bb3_cmp36_0_stall_in_0_reg_171_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 159
//  * capacity = 159
 logic rnode_171to330_bb3_cmp36_0_valid_out_NO_SHIFT_REG;
 logic rnode_171to330_bb3_cmp36_0_stall_in_NO_SHIFT_REG;
 logic rnode_171to330_bb3_cmp36_0_NO_SHIFT_REG;
 logic rnode_171to330_bb3_cmp36_0_reg_330_inputs_ready_NO_SHIFT_REG;
 logic rnode_171to330_bb3_cmp36_0_reg_330_NO_SHIFT_REG;
 logic rnode_171to330_bb3_cmp36_0_valid_out_reg_330_NO_SHIFT_REG;
 logic rnode_171to330_bb3_cmp36_0_stall_in_reg_330_NO_SHIFT_REG;
 logic rnode_171to330_bb3_cmp36_0_stall_out_reg_330_NO_SHIFT_REG;

acl_data_fifo rnode_171to330_bb3_cmp36_0_reg_330_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to330_bb3_cmp36_0_reg_330_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to330_bb3_cmp36_0_stall_in_reg_330_NO_SHIFT_REG),
	.valid_out(rnode_171to330_bb3_cmp36_0_valid_out_reg_330_NO_SHIFT_REG),
	.stall_out(rnode_171to330_bb3_cmp36_0_stall_out_reg_330_NO_SHIFT_REG),
	.data_in(rnode_171to171_bb3_cmp36_0_NO_SHIFT_REG),
	.data_out(rnode_171to330_bb3_cmp36_0_reg_330_NO_SHIFT_REG)
);

defparam rnode_171to330_bb3_cmp36_0_reg_330_fifo.DEPTH = 160;
defparam rnode_171to330_bb3_cmp36_0_reg_330_fifo.DATA_WIDTH = 1;
defparam rnode_171to330_bb3_cmp36_0_reg_330_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_171to330_bb3_cmp36_0_reg_330_fifo.IMPL = "ram";

assign rnode_171to330_bb3_cmp36_0_reg_330_inputs_ready_NO_SHIFT_REG = rnode_171to171_bb3_cmp36_0_valid_out_0_NO_SHIFT_REG;
assign rnode_171to171_bb3_cmp36_0_stall_in_0_NO_SHIFT_REG = rnode_171to330_bb3_cmp36_0_stall_out_reg_330_NO_SHIFT_REG;
assign rnode_171to330_bb3_cmp36_0_NO_SHIFT_REG = rnode_171to330_bb3_cmp36_0_reg_330_NO_SHIFT_REG;
assign rnode_171to330_bb3_cmp36_0_stall_in_reg_330_NO_SHIFT_REG = rnode_171to330_bb3_cmp36_0_stall_in_NO_SHIFT_REG;
assign rnode_171to330_bb3_cmp36_0_valid_out_NO_SHIFT_REG = rnode_171to330_bb3_cmp36_0_valid_out_reg_330_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp36_xor_stall_local;
wire local_bb3_cmp36_xor;
wire [96:0] rci_rcnode_330to331_rc0_t_119_0_reg_330;

assign local_bb3_cmp36_xor = (rnode_171to171_bb3_cmp36_1_NO_SHIFT_REG ^ 1'b1);
assign rci_rcnode_330to331_rc0_t_119_0_reg_330[31:0] = rcnode_1to330_rc8_t_119_0_NO_SHIFT_REG[31:0];
assign rci_rcnode_330to331_rc0_t_119_0_reg_330[63:32] = rcnode_1to330_rc8_t_119_0_NO_SHIFT_REG[63:32];
assign rci_rcnode_330to331_rc0_t_119_0_reg_330[64] = rnode_171to330_bb3_cmp36_0_NO_SHIFT_REG;
assign rci_rcnode_330to331_rc0_t_119_0_reg_330[96:65] = rnode_168to330_bb3_ld__0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_330to331_rc0_t_119_0_valid_out_0_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_stall_in_0_NO_SHIFT_REG;
 logic [96:0] rcnode_330to331_rc0_t_119_0_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_valid_out_1_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_stall_in_1_NO_SHIFT_REG;
 logic [96:0] rcnode_330to331_rc0_t_119_1_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_valid_out_2_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_stall_in_2_NO_SHIFT_REG;
 logic [96:0] rcnode_330to331_rc0_t_119_2_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_valid_out_3_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_stall_in_3_NO_SHIFT_REG;
 logic [96:0] rcnode_330to331_rc0_t_119_3_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_reg_331_inputs_ready_NO_SHIFT_REG;
 logic [96:0] rcnode_330to331_rc0_t_119_0_reg_331_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_valid_out_0_reg_331_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_stall_in_0_reg_331_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_IP_NO_SHIFT_REG;
 logic rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_NO_SHIFT_REG;

acl_data_fifo rcnode_330to331_rc0_t_119_0_reg_331_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_330to331_rc0_t_119_0_reg_331_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_330to331_rc0_t_119_0_stall_in_0_reg_331_NO_SHIFT_REG),
	.valid_out(rcnode_330to331_rc0_t_119_0_valid_out_0_reg_331_NO_SHIFT_REG),
	.stall_out(rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_330to331_rc0_t_119_0_reg_330),
	.data_out(rcnode_330to331_rc0_t_119_0_reg_331_NO_SHIFT_REG)
);

defparam rcnode_330to331_rc0_t_119_0_reg_331_fifo.DEPTH = 1;
defparam rcnode_330to331_rc0_t_119_0_reg_331_fifo.DATA_WIDTH = 97;
defparam rcnode_330to331_rc0_t_119_0_reg_331_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_330to331_rc0_t_119_0_reg_331_fifo.IMPL = "ll_reg";

assign rcnode_330to331_rc0_t_119_0_reg_331_inputs_ready_NO_SHIFT_REG = (rnode_171to330_bb3_cmp36_0_valid_out_NO_SHIFT_REG & rnode_168to330_bb3_ld__0_valid_out_NO_SHIFT_REG & rcnode_1to330_rc8_t_119_0_valid_out_NO_SHIFT_REG);
assign rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_NO_SHIFT_REG = (~(rcnode_330to331_rc0_t_119_0_reg_331_inputs_ready_NO_SHIFT_REG) | rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_IP_NO_SHIFT_REG);
assign rnode_171to330_bb3_cmp36_0_stall_in_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_NO_SHIFT_REG;
assign rnode_168to330_bb3_ld__0_stall_in_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_NO_SHIFT_REG;
assign rcnode_1to330_rc8_t_119_0_stall_in_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_stall_out_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_0_stall_in_0_reg_331_NO_SHIFT_REG = (rcnode_330to331_rc0_t_119_0_stall_in_0_NO_SHIFT_REG | rcnode_330to331_rc0_t_119_0_stall_in_1_NO_SHIFT_REG | rcnode_330to331_rc0_t_119_0_stall_in_2_NO_SHIFT_REG | rcnode_330to331_rc0_t_119_0_stall_in_3_NO_SHIFT_REG);
assign rcnode_330to331_rc0_t_119_0_valid_out_0_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_valid_out_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_0_valid_out_1_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_valid_out_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_0_valid_out_2_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_valid_out_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_0_valid_out_3_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_valid_out_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_0_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_1_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_2_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_reg_331_NO_SHIFT_REG;
assign rcnode_330to331_rc0_t_119_3_NO_SHIFT_REG = rcnode_330to331_rc0_t_119_0_reg_331_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__phi_decision45_or46_valid_out;
wire local_bb3__phi_decision45_or46_stall_in;
wire local_bb3__phi_decision45_or46_inputs_ready;
wire local_bb3__phi_decision45_or46_stall_local;
wire local_bb3__phi_decision45_or46;

assign local_bb3__phi_decision45_or46_inputs_ready = (rnode_170to171_var__u8_0_valid_out_0_NO_SHIFT_REG & rnode_171to171_bb3_cmp36_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3__phi_decision45_or46 = (rnode_170to171_var__u8_0_NO_SHIFT_REG | local_bb3_cmp36_xor);
assign local_bb3__phi_decision45_or46_valid_out = local_bb3__phi_decision45_or46_inputs_ready;
assign local_bb3__phi_decision45_or46_stall_local = local_bb3__phi_decision45_or46_stall_in;
assign rnode_170to171_var__u8_0_stall_in_0_NO_SHIFT_REG = (local_bb3__phi_decision45_or46_stall_local | ~(local_bb3__phi_decision45_or46_inputs_ready));
assign rnode_171to171_bb3_cmp36_0_stall_in_1_NO_SHIFT_REG = (local_bb3__phi_decision45_or46_stall_local | ~(local_bb3__phi_decision45_or46_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni1_stall_local;
wire [255:0] local_bb3_c0_eni1;

assign local_bb3_c0_eni1[31:0] = 32'bx;
assign local_bb3_c0_eni1[63:32] = rcnode_330to331_rc0_t_119_0_NO_SHIFT_REG[96:65];
assign local_bb3_c0_eni1[255:64] = 192'bx;

// This section implements a staging register.
// 
wire rstag_171to171_bb3__phi_decision45_or46_valid_out_0;
wire rstag_171to171_bb3__phi_decision45_or46_stall_in_0;
wire rstag_171to171_bb3__phi_decision45_or46_valid_out_1;
wire rstag_171to171_bb3__phi_decision45_or46_stall_in_1;
wire rstag_171to171_bb3__phi_decision45_or46_inputs_ready;
wire rstag_171to171_bb3__phi_decision45_or46_stall_local;
 reg rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG;
wire rstag_171to171_bb3__phi_decision45_or46_combined_valid;
 reg rstag_171to171_bb3__phi_decision45_or46_staging_reg_NO_SHIFT_REG;
wire rstag_171to171_bb3__phi_decision45_or46;
 reg rstag_171to171_bb3__phi_decision45_or46_consumed_0_NO_SHIFT_REG;
 reg rstag_171to171_bb3__phi_decision45_or46_consumed_1_NO_SHIFT_REG;

assign rstag_171to171_bb3__phi_decision45_or46_inputs_ready = local_bb3__phi_decision45_or46_valid_out;
assign rstag_171to171_bb3__phi_decision45_or46 = (rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG ? rstag_171to171_bb3__phi_decision45_or46_staging_reg_NO_SHIFT_REG : local_bb3__phi_decision45_or46);
assign rstag_171to171_bb3__phi_decision45_or46_combined_valid = (rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG | rstag_171to171_bb3__phi_decision45_or46_inputs_ready);
assign rstag_171to171_bb3__phi_decision45_or46_stall_local = ((rstag_171to171_bb3__phi_decision45_or46_stall_in_0 & ~(rstag_171to171_bb3__phi_decision45_or46_consumed_0_NO_SHIFT_REG)) | (rstag_171to171_bb3__phi_decision45_or46_stall_in_1 & ~(rstag_171to171_bb3__phi_decision45_or46_consumed_1_NO_SHIFT_REG)));
assign rstag_171to171_bb3__phi_decision45_or46_valid_out_0 = (rstag_171to171_bb3__phi_decision45_or46_combined_valid & ~(rstag_171to171_bb3__phi_decision45_or46_consumed_0_NO_SHIFT_REG));
assign rstag_171to171_bb3__phi_decision45_or46_valid_out_1 = (rstag_171to171_bb3__phi_decision45_or46_combined_valid & ~(rstag_171to171_bb3__phi_decision45_or46_consumed_1_NO_SHIFT_REG));
assign local_bb3__phi_decision45_or46_stall_in = (|rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_171to171_bb3__phi_decision45_or46_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_171to171_bb3__phi_decision45_or46_stall_local)
		begin
			if (~(rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG))
			begin
				rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG <= rstag_171to171_bb3__phi_decision45_or46_inputs_ready;
			end
		end
		else
		begin
			rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_171to171_bb3__phi_decision45_or46_staging_valid_NO_SHIFT_REG))
		begin
			rstag_171to171_bb3__phi_decision45_or46_staging_reg_NO_SHIFT_REG <= local_bb3__phi_decision45_or46;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_171to171_bb3__phi_decision45_or46_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_171to171_bb3__phi_decision45_or46_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_171to171_bb3__phi_decision45_or46_consumed_0_NO_SHIFT_REG <= (rstag_171to171_bb3__phi_decision45_or46_combined_valid & (rstag_171to171_bb3__phi_decision45_or46_consumed_0_NO_SHIFT_REG | ~(rstag_171to171_bb3__phi_decision45_or46_stall_in_0)) & rstag_171to171_bb3__phi_decision45_or46_stall_local);
		rstag_171to171_bb3__phi_decision45_or46_consumed_1_NO_SHIFT_REG <= (rstag_171to171_bb3__phi_decision45_or46_combined_valid & (rstag_171to171_bb3__phi_decision45_or46_consumed_1_NO_SHIFT_REG | ~(rstag_171to171_bb3__phi_decision45_or46_stall_in_1)) & rstag_171to171_bb3__phi_decision45_or46_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni2_stall_local;
wire [255:0] local_bb3_c0_eni2;

assign local_bb3_c0_eni2[63:0] = local_bb3_c0_eni1[63:0];
assign local_bb3_c0_eni2[95:64] = rnode_330to331_ld__0_NO_SHIFT_REG;
assign local_bb3_c0_eni2[255:96] = local_bb3_c0_eni1[255:96];

// This section implements a registered operation.
// 
wire local_bb3_ld__u12_inputs_ready;
 reg local_bb3_ld__u12_valid_out_NO_SHIFT_REG;
wire local_bb3_ld__u12_stall_in;
wire local_bb3_ld__u12_output_regs_ready;
wire local_bb3_ld__u12_fu_stall_out;
wire local_bb3_ld__u12_fu_valid_out;
wire [31:0] local_bb3_ld__u12_lsu_dataout;
 reg [31:0] local_bb3_ld__u12_NO_SHIFT_REG;
wire local_bb3_ld__u12_causedstall;

lsu_top lsu_local_bb3_ld__u12 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb3_ld__u12_fu_stall_out),
	.i_valid(local_bb3_ld__u12_inputs_ready),
	.i_address((rnode_170to171_bb3_arrayidx46_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_171to171_bb3__phi_decision45_or46),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb3_ld__u12_output_regs_ready)),
	.o_valid(local_bb3_ld__u12_fu_valid_out),
	.o_readdata(local_bb3_ld__u12_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb3_ld__u12_active),
	.avm_address(avm_local_bb3_ld__u12_address),
	.avm_read(avm_local_bb3_ld__u12_read),
	.avm_readdata(avm_local_bb3_ld__u12_readdata),
	.avm_write(avm_local_bb3_ld__u12_write),
	.avm_writeack(avm_local_bb3_ld__u12_writeack),
	.avm_burstcount(avm_local_bb3_ld__u12_burstcount),
	.avm_writedata(avm_local_bb3_ld__u12_writedata),
	.avm_byteenable(avm_local_bb3_ld__u12_byteenable),
	.avm_waitrequest(avm_local_bb3_ld__u12_waitrequest),
	.avm_readdatavalid(avm_local_bb3_ld__u12_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb3_ld__u12.AWIDTH = 33;
defparam lsu_local_bb3_ld__u12.WIDTH_BYTES = 4;
defparam lsu_local_bb3_ld__u12.MWIDTH_BYTES = 64;
defparam lsu_local_bb3_ld__u12.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb3_ld__u12.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb3_ld__u12.READ = 1;
defparam lsu_local_bb3_ld__u12.ATOMIC = 0;
defparam lsu_local_bb3_ld__u12.WIDTH = 32;
defparam lsu_local_bb3_ld__u12.MWIDTH = 512;
defparam lsu_local_bb3_ld__u12.ATOMIC_WIDTH = 3;
defparam lsu_local_bb3_ld__u12.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb3_ld__u12.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb3_ld__u12.MEMORY_SIDE_MEM_LATENCY = 132;
defparam lsu_local_bb3_ld__u12.USE_WRITE_ACK = 0;
defparam lsu_local_bb3_ld__u12.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb3_ld__u12.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb3_ld__u12.NUMBER_BANKS = 1;
defparam lsu_local_bb3_ld__u12.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb3_ld__u12.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb3_ld__u12.USEINPUTFIFO = 0;
defparam lsu_local_bb3_ld__u12.USECACHING = 1;
defparam lsu_local_bb3_ld__u12.CACHESIZE = 1024;
defparam lsu_local_bb3_ld__u12.USEOUTPUTFIFO = 1;
defparam lsu_local_bb3_ld__u12.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb3_ld__u12.HIGH_FMAX = 1;
defparam lsu_local_bb3_ld__u12.ADDRSPACE = 1;
defparam lsu_local_bb3_ld__u12.STYLE = "BURST-COALESCED";

assign local_bb3_ld__u12_inputs_ready = (rnode_170to171_bb3_arrayidx46_0_valid_out_NO_SHIFT_REG & rstag_171to171_bb3__phi_decision45_or46_valid_out_0);
assign local_bb3_ld__u12_output_regs_ready = (&(~(local_bb3_ld__u12_valid_out_NO_SHIFT_REG) | ~(local_bb3_ld__u12_stall_in)));
assign rnode_170to171_bb3_arrayidx46_0_stall_in_NO_SHIFT_REG = (local_bb3_ld__u12_fu_stall_out | ~(local_bb3_ld__u12_inputs_ready));
assign rstag_171to171_bb3__phi_decision45_or46_stall_in_0 = (local_bb3_ld__u12_fu_stall_out | ~(local_bb3_ld__u12_inputs_ready));
assign local_bb3_ld__u12_causedstall = (local_bb3_ld__u12_inputs_ready && (local_bb3_ld__u12_fu_stall_out && !(~(local_bb3_ld__u12_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_ld__u12_NO_SHIFT_REG <= 'x;
		local_bb3_ld__u12_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_ld__u12_output_regs_ready)
		begin
			local_bb3_ld__u12_NO_SHIFT_REG <= local_bb3_ld__u12_lsu_dataout;
			local_bb3_ld__u12_valid_out_NO_SHIFT_REG <= local_bb3_ld__u12_fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_ld__u12_stall_in))
			begin
				local_bb3_ld__u12_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_ld__u13_inputs_ready;
 reg local_bb3_ld__u13_valid_out_NO_SHIFT_REG;
wire local_bb3_ld__u13_stall_in;
wire local_bb3_ld__u13_output_regs_ready;
wire local_bb3_ld__u13_fu_stall_out;
wire local_bb3_ld__u13_fu_valid_out;
wire [31:0] local_bb3_ld__u13_lsu_dataout;
 reg [31:0] local_bb3_ld__u13_NO_SHIFT_REG;
wire local_bb3_ld__u13_causedstall;

lsu_top lsu_local_bb3_ld__u13 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb3_ld__u13_fu_stall_out),
	.i_valid(local_bb3_ld__u13_inputs_ready),
	.i_address((rnode_170to171_arrayidx43_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_171to171_bb3__phi_decision45_or46),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb3_ld__u13_output_regs_ready)),
	.o_valid(local_bb3_ld__u13_fu_valid_out),
	.o_readdata(local_bb3_ld__u13_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb3_ld__u13_active),
	.avm_address(avm_local_bb3_ld__u13_address),
	.avm_read(avm_local_bb3_ld__u13_read),
	.avm_readdata(avm_local_bb3_ld__u13_readdata),
	.avm_write(avm_local_bb3_ld__u13_write),
	.avm_writeack(avm_local_bb3_ld__u13_writeack),
	.avm_burstcount(avm_local_bb3_ld__u13_burstcount),
	.avm_writedata(avm_local_bb3_ld__u13_writedata),
	.avm_byteenable(avm_local_bb3_ld__u13_byteenable),
	.avm_waitrequest(avm_local_bb3_ld__u13_waitrequest),
	.avm_readdatavalid(avm_local_bb3_ld__u13_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb3_ld__u13.AWIDTH = 33;
defparam lsu_local_bb3_ld__u13.WIDTH_BYTES = 4;
defparam lsu_local_bb3_ld__u13.MWIDTH_BYTES = 64;
defparam lsu_local_bb3_ld__u13.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb3_ld__u13.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb3_ld__u13.READ = 1;
defparam lsu_local_bb3_ld__u13.ATOMIC = 0;
defparam lsu_local_bb3_ld__u13.WIDTH = 32;
defparam lsu_local_bb3_ld__u13.MWIDTH = 512;
defparam lsu_local_bb3_ld__u13.ATOMIC_WIDTH = 3;
defparam lsu_local_bb3_ld__u13.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb3_ld__u13.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb3_ld__u13.MEMORY_SIDE_MEM_LATENCY = 132;
defparam lsu_local_bb3_ld__u13.USE_WRITE_ACK = 0;
defparam lsu_local_bb3_ld__u13.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb3_ld__u13.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb3_ld__u13.NUMBER_BANKS = 1;
defparam lsu_local_bb3_ld__u13.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb3_ld__u13.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb3_ld__u13.USEINPUTFIFO = 0;
defparam lsu_local_bb3_ld__u13.USECACHING = 1;
defparam lsu_local_bb3_ld__u13.CACHESIZE = 1024;
defparam lsu_local_bb3_ld__u13.USEOUTPUTFIFO = 1;
defparam lsu_local_bb3_ld__u13.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb3_ld__u13.HIGH_FMAX = 1;
defparam lsu_local_bb3_ld__u13.ADDRSPACE = 1;
defparam lsu_local_bb3_ld__u13.STYLE = "BURST-COALESCED";

assign local_bb3_ld__u13_inputs_ready = (rnode_170to171_arrayidx43_0_valid_out_0_NO_SHIFT_REG & rstag_171to171_bb3__phi_decision45_or46_valid_out_1);
assign local_bb3_ld__u13_output_regs_ready = (&(~(local_bb3_ld__u13_valid_out_NO_SHIFT_REG) | ~(local_bb3_ld__u13_stall_in)));
assign rnode_170to171_arrayidx43_0_stall_in_0_NO_SHIFT_REG = (local_bb3_ld__u13_fu_stall_out | ~(local_bb3_ld__u13_inputs_ready));
assign rstag_171to171_bb3__phi_decision45_or46_stall_in_1 = (local_bb3_ld__u13_fu_stall_out | ~(local_bb3_ld__u13_inputs_ready));
assign local_bb3_ld__u13_causedstall = (local_bb3_ld__u13_inputs_ready && (local_bb3_ld__u13_fu_stall_out && !(~(local_bb3_ld__u13_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_ld__u13_NO_SHIFT_REG <= 'x;
		local_bb3_ld__u13_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_ld__u13_output_regs_ready)
		begin
			local_bb3_ld__u13_NO_SHIFT_REG <= local_bb3_ld__u13_lsu_dataout;
			local_bb3_ld__u13_valid_out_NO_SHIFT_REG <= local_bb3_ld__u13_fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_ld__u13_stall_in))
			begin
				local_bb3_ld__u13_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_331to331_bb3_ld__u12_valid_out;
wire rstag_331to331_bb3_ld__u12_stall_in;
wire rstag_331to331_bb3_ld__u12_inputs_ready;
wire rstag_331to331_bb3_ld__u12_stall_local;
 reg rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG;
wire rstag_331to331_bb3_ld__u12_combined_valid;
 reg [31:0] rstag_331to331_bb3_ld__u12_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_331to331_bb3_ld__u12;

assign rstag_331to331_bb3_ld__u12_inputs_ready = local_bb3_ld__u12_valid_out_NO_SHIFT_REG;
assign rstag_331to331_bb3_ld__u12 = (rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG ? rstag_331to331_bb3_ld__u12_staging_reg_NO_SHIFT_REG : local_bb3_ld__u12_NO_SHIFT_REG);
assign rstag_331to331_bb3_ld__u12_combined_valid = (rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG | rstag_331to331_bb3_ld__u12_inputs_ready);
assign rstag_331to331_bb3_ld__u12_valid_out = rstag_331to331_bb3_ld__u12_combined_valid;
assign rstag_331to331_bb3_ld__u12_stall_local = rstag_331to331_bb3_ld__u12_stall_in;
assign local_bb3_ld__u12_stall_in = (|rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_331to331_bb3_ld__u12_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_331to331_bb3_ld__u12_stall_local)
		begin
			if (~(rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG))
			begin
				rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG <= rstag_331to331_bb3_ld__u12_inputs_ready;
			end
		end
		else
		begin
			rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_331to331_bb3_ld__u12_staging_valid_NO_SHIFT_REG))
		begin
			rstag_331to331_bb3_ld__u12_staging_reg_NO_SHIFT_REG <= local_bb3_ld__u12_NO_SHIFT_REG;
		end
	end
end


// This section implements a staging register.
// 
wire rstag_331to331_bb3_ld__u13_valid_out;
wire rstag_331to331_bb3_ld__u13_stall_in;
wire rstag_331to331_bb3_ld__u13_inputs_ready;
wire rstag_331to331_bb3_ld__u13_stall_local;
 reg rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG;
wire rstag_331to331_bb3_ld__u13_combined_valid;
 reg [31:0] rstag_331to331_bb3_ld__u13_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_331to331_bb3_ld__u13;

assign rstag_331to331_bb3_ld__u13_inputs_ready = local_bb3_ld__u13_valid_out_NO_SHIFT_REG;
assign rstag_331to331_bb3_ld__u13 = (rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG ? rstag_331to331_bb3_ld__u13_staging_reg_NO_SHIFT_REG : local_bb3_ld__u13_NO_SHIFT_REG);
assign rstag_331to331_bb3_ld__u13_combined_valid = (rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG | rstag_331to331_bb3_ld__u13_inputs_ready);
assign rstag_331to331_bb3_ld__u13_valid_out = rstag_331to331_bb3_ld__u13_combined_valid;
assign rstag_331to331_bb3_ld__u13_stall_local = rstag_331to331_bb3_ld__u13_stall_in;
assign local_bb3_ld__u13_stall_in = (|rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_331to331_bb3_ld__u13_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_331to331_bb3_ld__u13_stall_local)
		begin
			if (~(rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG))
			begin
				rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG <= rstag_331to331_bb3_ld__u13_inputs_ready;
			end
		end
		else
		begin
			rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_331to331_bb3_ld__u13_staging_valid_NO_SHIFT_REG))
		begin
			rstag_331to331_bb3_ld__u13_staging_reg_NO_SHIFT_REG <= local_bb3_ld__u13_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni3_stall_local;
wire [255:0] local_bb3_c0_eni3;

assign local_bb3_c0_eni3[95:0] = local_bb3_c0_eni2[95:0];
assign local_bb3_c0_eni3[127:96] = rstag_331to331_bb3_ld__u13;
assign local_bb3_c0_eni3[255:128] = local_bb3_c0_eni2[255:128];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni4_stall_local;
wire [255:0] local_bb3_c0_eni4;

assign local_bb3_c0_eni4[127:0] = local_bb3_c0_eni3[127:0];
assign local_bb3_c0_eni4[159:128] = rstag_331to331_bb3_ld__u12;
assign local_bb3_c0_eni4[255:160] = local_bb3_c0_eni3[255:160];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni5_stall_local;
wire [255:0] local_bb3_c0_eni5;

assign local_bb3_c0_eni5[159:0] = local_bb3_c0_eni4[159:0];
assign local_bb3_c0_eni5[191:160] = rcnode_330to331_rc0_t_119_0_NO_SHIFT_REG[31:0];
assign local_bb3_c0_eni5[255:192] = local_bb3_c0_eni4[255:192];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni6_stall_local;
wire [255:0] local_bb3_c0_eni6;

assign local_bb3_c0_eni6[191:0] = local_bb3_c0_eni5[191:0];
assign local_bb3_c0_eni6[223:192] = rcnode_330to331_rc0_t_119_0_NO_SHIFT_REG[63:32];
assign local_bb3_c0_eni6[255:224] = local_bb3_c0_eni5[255:224];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni7_valid_out;
wire local_bb3_c0_eni7_stall_in;
wire local_bb3_c0_eni7_inputs_ready;
wire local_bb3_c0_eni7_stall_local;
wire [255:0] local_bb3_c0_eni7;

assign local_bb3_c0_eni7_inputs_ready = (rnode_330to331_ld__0_valid_out_0_NO_SHIFT_REG & rstag_331to331_bb3_ld__u13_valid_out & rcnode_330to331_rc0_t_119_0_valid_out_3_NO_SHIFT_REG & rstag_331to331_bb3_ld__u12_valid_out & rcnode_330to331_rc0_t_119_0_valid_out_0_NO_SHIFT_REG & rcnode_330to331_rc0_t_119_0_valid_out_1_NO_SHIFT_REG & rcnode_330to331_rc0_t_119_0_valid_out_2_NO_SHIFT_REG);
assign local_bb3_c0_eni7[223:0] = local_bb3_c0_eni6[223:0];
assign local_bb3_c0_eni7[224] = rcnode_330to331_rc0_t_119_0_NO_SHIFT_REG[64];
assign local_bb3_c0_eni7[255:225] = local_bb3_c0_eni6[255:225];
assign local_bb3_c0_eni7_valid_out = local_bb3_c0_eni7_inputs_ready;
assign local_bb3_c0_eni7_stall_local = local_bb3_c0_eni7_stall_in;
assign rnode_330to331_ld__0_stall_in_0_NO_SHIFT_REG = (local_bb3_c0_eni7_stall_local | ~(local_bb3_c0_eni7_inputs_ready));
assign rstag_331to331_bb3_ld__u13_stall_in = (local_bb3_c0_eni7_stall_local | ~(local_bb3_c0_eni7_inputs_ready));
assign rcnode_330to331_rc0_t_119_0_stall_in_3_NO_SHIFT_REG = (local_bb3_c0_eni7_stall_local | ~(local_bb3_c0_eni7_inputs_ready));
assign rstag_331to331_bb3_ld__u12_stall_in = (local_bb3_c0_eni7_stall_local | ~(local_bb3_c0_eni7_inputs_ready));
assign rcnode_330to331_rc0_t_119_0_stall_in_0_NO_SHIFT_REG = (local_bb3_c0_eni7_stall_local | ~(local_bb3_c0_eni7_inputs_ready));
assign rcnode_330to331_rc0_t_119_0_stall_in_1_NO_SHIFT_REG = (local_bb3_c0_eni7_stall_local | ~(local_bb3_c0_eni7_inputs_ready));
assign rcnode_330to331_rc0_t_119_0_stall_in_2_NO_SHIFT_REG = (local_bb3_c0_eni7_stall_local | ~(local_bb3_c0_eni7_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb3_c0_enter_c0_eni7_inputs_ready;
 reg local_bb3_c0_enter_c0_eni7_valid_out_0_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_0;
 reg local_bb3_c0_enter_c0_eni7_valid_out_1_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_1;
 reg local_bb3_c0_enter_c0_eni7_valid_out_2_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_2;
 reg local_bb3_c0_enter_c0_eni7_valid_out_3_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_3;
 reg local_bb3_c0_enter_c0_eni7_valid_out_4_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_4;
 reg local_bb3_c0_enter_c0_eni7_valid_out_5_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_5;
 reg local_bb3_c0_enter_c0_eni7_valid_out_6_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_6;
 reg local_bb3_c0_enter_c0_eni7_valid_out_7_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_stall_in_7;
wire local_bb3_c0_enter_c0_eni7_output_regs_ready;
 reg [255:0] local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG;
wire local_bb3_c0_enter_c0_eni7_input_accepted;
 reg local_bb3_c0_enter_c0_eni7_valid_bit_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi2_entry_stall;
wire local_bb3_c0_exit_c0_exi2_output_regs_ready;
wire [63:0] local_bb3_c0_exit_c0_exi2_valid_bits;
wire local_bb3_c0_exit_c0_exi2_valid_in;
wire local_bb3_c0_exit_c0_exi2_phases;
wire local_bb3_c0_enter_c0_eni7_inc_pipelined_thread;
wire local_bb3_c0_enter_c0_eni7_dec_pipelined_thread;
wire local_bb3_c0_enter_c0_eni7_causedstall;

assign local_bb3_c0_enter_c0_eni7_inputs_ready = local_bb3_c0_eni7_valid_out;
assign local_bb3_c0_enter_c0_eni7_output_regs_ready = 1'b1;
assign local_bb3_c0_enter_c0_eni7_input_accepted = (local_bb3_c0_enter_c0_eni7_inputs_ready && !(local_bb3_c0_exit_c0_exi2_entry_stall));
assign local_bb3_c0_enter_c0_eni7_inc_pipelined_thread = 1'b1;
assign local_bb3_c0_enter_c0_eni7_dec_pipelined_thread = ~(1'b0);
assign local_bb3_c0_eni7_stall_in = ((~(local_bb3_c0_enter_c0_eni7_inputs_ready) | local_bb3_c0_exit_c0_exi2_entry_stall) | ~(1'b1));
assign local_bb3_c0_enter_c0_eni7_causedstall = (1'b1 && ((~(local_bb3_c0_enter_c0_eni7_inputs_ready) | local_bb3_c0_exit_c0_exi2_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_c0_enter_c0_eni7_valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb3_c0_enter_c0_eni7_valid_bit_NO_SHIFT_REG <= local_bb3_c0_enter_c0_eni7_input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG <= 'x;
		local_bb3_c0_enter_c0_eni7_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_enter_c0_eni7_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_enter_c0_eni7_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_enter_c0_eni7_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_enter_c0_eni7_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_enter_c0_eni7_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_enter_c0_eni7_valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_enter_c0_eni7_valid_out_7_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_c0_enter_c0_eni7_output_regs_ready)
		begin
			local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG <= local_bb3_c0_eni7;
			local_bb3_c0_enter_c0_eni7_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_c0_enter_c0_eni7_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb3_c0_enter_c0_eni7_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb3_c0_enter_c0_eni7_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb3_c0_enter_c0_eni7_valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb3_c0_enter_c0_eni7_valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb3_c0_enter_c0_eni7_valid_out_6_NO_SHIFT_REG <= 1'b1;
			local_bb3_c0_enter_c0_eni7_valid_out_7_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_0))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_1))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_2))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_3))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_4))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_5))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_6))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_enter_c0_eni7_stall_in_7))
			begin
				local_bb3_c0_enter_c0_eni7_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_stall_local;
wire [31:0] local_bb3_c0_ene1;

assign local_bb3_c0_ene1 = local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene2_stall_local;
wire [31:0] local_bb3_c0_ene2;

assign local_bb3_c0_ene2 = local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG[95:64];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene3_stall_local;
wire [31:0] local_bb3_c0_ene3;

assign local_bb3_c0_ene3 = local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG[127:96];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene4_stall_local;
wire [31:0] local_bb3_c0_ene4;

assign local_bb3_c0_ene4 = local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG[159:128];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene5_valid_out;
wire local_bb3_c0_ene5_stall_in;
wire local_bb3_c0_ene5_inputs_ready;
wire local_bb3_c0_ene5_stall_local;
wire [31:0] local_bb3_c0_ene5;

assign local_bb3_c0_ene5_inputs_ready = local_bb3_c0_enter_c0_eni7_valid_out_4_NO_SHIFT_REG;
assign local_bb3_c0_ene5 = local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG[191:160];
assign local_bb3_c0_ene5_valid_out = 1'b1;
assign local_bb3_c0_enter_c0_eni7_stall_in_4 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene6_valid_out;
wire local_bb3_c0_ene6_stall_in;
wire local_bb3_c0_ene6_inputs_ready;
wire local_bb3_c0_ene6_stall_local;
wire [31:0] local_bb3_c0_ene6;

assign local_bb3_c0_ene6_inputs_ready = local_bb3_c0_enter_c0_eni7_valid_out_5_NO_SHIFT_REG;
assign local_bb3_c0_ene6 = local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG[223:192];
assign local_bb3_c0_ene6_valid_out = 1'b1;
assign local_bb3_c0_enter_c0_eni7_stall_in_5 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene7_valid_out;
wire local_bb3_c0_ene7_stall_in;
wire local_bb3_c0_ene7_inputs_ready;
wire local_bb3_c0_ene7_stall_local;
wire local_bb3_c0_ene7;

assign local_bb3_c0_ene7_inputs_ready = local_bb3_c0_enter_c0_eni7_valid_out_6_NO_SHIFT_REG;
assign local_bb3_c0_ene7 = local_bb3_c0_enter_c0_eni7_NO_SHIFT_REG[224];
assign local_bb3_c0_ene7_valid_out = 1'b1;
assign local_bb3_c0_enter_c0_eni7_stall_in_6 = 1'b0;

// This section implements an unregistered operation.
// 
wire SFC_1_VALID_332_332_0_valid_out;
wire SFC_1_VALID_332_332_0_stall_in;
wire SFC_1_VALID_332_332_0_inputs_ready;
wire SFC_1_VALID_332_332_0_stall_local;
wire SFC_1_VALID_332_332_0;

assign SFC_1_VALID_332_332_0_inputs_ready = local_bb3_c0_enter_c0_eni7_valid_out_7_NO_SHIFT_REG;
assign SFC_1_VALID_332_332_0 = local_bb3_c0_enter_c0_eni7_valid_bit_NO_SHIFT_REG;
assign SFC_1_VALID_332_332_0_valid_out = 1'b1;
assign local_bb3_c0_enter_c0_eni7_stall_in_7 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u14_stall_local;
wire [31:0] local_bb3_var__u14;

assign local_bb3_var__u14 = local_bb3_c0_ene1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u15_stall_local;
wire [31:0] local_bb3_var__u15;

assign local_bb3_var__u15 = local_bb3_c0_ene2;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u16_stall_local;
wire [31:0] local_bb3_var__u16;

assign local_bb3_var__u16 = local_bb3_c0_ene3;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u17_stall_local;
wire [31:0] local_bb3_var__u17;

assign local_bb3_var__u17 = local_bb3_c0_ene4;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene5_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_c0_ene5_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene5_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene5_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene5_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_c0_ene5_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_c0_ene5_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_c0_ene5_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_c0_ene5_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_c0_ene5_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene5),
	.data_out(rnode_332to333_bb3_c0_ene5_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_c0_ene5_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_c0_ene5_0_reg_333_fifo.DATA_WIDTH = 32;
defparam rnode_332to333_bb3_c0_ene5_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_c0_ene5_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_c0_ene5_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene5_stall_in = 1'b0;
assign rnode_332to333_bb3_c0_ene5_0_NO_SHIFT_REG = rnode_332to333_bb3_c0_ene5_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_c0_ene5_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene6_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_c0_ene6_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene6_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene6_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene6_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_c0_ene6_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_c0_ene6_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_c0_ene6_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_c0_ene6_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_c0_ene6_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene6),
	.data_out(rnode_332to333_bb3_c0_ene6_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_c0_ene6_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_c0_ene6_0_reg_333_fifo.DATA_WIDTH = 32;
defparam rnode_332to333_bb3_c0_ene6_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_c0_ene6_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_c0_ene6_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene6_stall_in = 1'b0;
assign rnode_332to333_bb3_c0_ene6_0_NO_SHIFT_REG = rnode_332to333_bb3_c0_ene6_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_c0_ene6_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene7_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene7_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene7_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene7_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene7_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_c0_ene7_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_c0_ene7_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_c0_ene7_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_c0_ene7_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_c0_ene7_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene7),
	.data_out(rnode_332to333_bb3_c0_ene7_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_c0_ene7_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_c0_ene7_0_reg_333_fifo.DATA_WIDTH = 1;
defparam rnode_332to333_bb3_c0_ene7_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_c0_ene7_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_c0_ene7_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene7_stall_in = 1'b0;
assign rnode_332to333_bb3_c0_ene7_0_NO_SHIFT_REG = rnode_332to333_bb3_c0_ene7_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_c0_ene7_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_332_333_0_inputs_ready;
 reg SFC_1_VALID_332_333_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_332_333_0_stall_in;
wire SFC_1_VALID_332_333_0_output_regs_ready;
 reg SFC_1_VALID_332_333_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_332_333_0_causedstall;

assign SFC_1_VALID_332_333_0_inputs_ready = 1'b1;
assign SFC_1_VALID_332_333_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_332_332_0_stall_in = 1'b0;
assign SFC_1_VALID_332_333_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_332_333_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_332_333_0_output_regs_ready)
		begin
			SFC_1_VALID_332_333_0_NO_SHIFT_REG <= SFC_1_VALID_332_332_0;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and2_i499_stall_local;
wire [31:0] local_bb3_and2_i499;

assign local_bb3_and2_i499 = (local_bb3_var__u14 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and12_i504_stall_local;
wire [31:0] local_bb3_and12_i504;

assign local_bb3_and12_i504 = (local_bb3_var__u14 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_xor_i496_stall_local;
wire [31:0] local_bb3_xor_i496;

assign local_bb3_xor_i496 = (local_bb3_var__u15 ^ 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i312_stall_local;
wire [31:0] local_bb3_shr_i312;

assign local_bb3_shr_i312 = (local_bb3_var__u16 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and5_i318_stall_local;
wire [31:0] local_bb3_and5_i318;

assign local_bb3_and5_i318 = (local_bb3_var__u16 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_shr2_i314_stall_local;
wire [31:0] local_bb3_shr2_i314;

assign local_bb3_shr2_i314 = (local_bb3_var__u17 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_xor_i316_stall_local;
wire [31:0] local_bb3_xor_i316;

assign local_bb3_xor_i316 = (local_bb3_var__u17 ^ local_bb3_var__u16);

// This section implements an unregistered operation.
// 
wire local_bb3_and6_i319_stall_local;
wire [31:0] local_bb3_and6_i319;

assign local_bb3_and6_i319 = (local_bb3_var__u17 & 32'h7FFFFF);

// Register node:
//  * latency = 52
//  * capacity = 52
 logic rnode_333to385_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to385_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_333to385_bb3_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_333to385_bb3_c0_ene5_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to385_bb3_c0_ene5_0_reg_385_NO_SHIFT_REG;
 logic rnode_333to385_bb3_c0_ene5_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_333to385_bb3_c0_ene5_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_333to385_bb3_c0_ene5_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_333to385_bb3_c0_ene5_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to385_bb3_c0_ene5_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to385_bb3_c0_ene5_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_333to385_bb3_c0_ene5_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_333to385_bb3_c0_ene5_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_333to385_bb3_c0_ene5_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_333to385_bb3_c0_ene5_0_reg_385_fifo.DEPTH = 52;
defparam rnode_333to385_bb3_c0_ene5_0_reg_385_fifo.DATA_WIDTH = 32;
defparam rnode_333to385_bb3_c0_ene5_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to385_bb3_c0_ene5_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_333to385_bb3_c0_ene5_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to385_bb3_c0_ene5_0_NO_SHIFT_REG = rnode_333to385_bb3_c0_ene5_0_reg_385_NO_SHIFT_REG;
assign rnode_333to385_bb3_c0_ene5_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_333to385_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 47
//  * capacity = 47
 logic rnode_333to380_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to380_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_333to380_bb3_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_333to380_bb3_c0_ene6_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to380_bb3_c0_ene6_0_reg_380_NO_SHIFT_REG;
 logic rnode_333to380_bb3_c0_ene6_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_333to380_bb3_c0_ene6_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_333to380_bb3_c0_ene6_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_333to380_bb3_c0_ene6_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to380_bb3_c0_ene6_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to380_bb3_c0_ene6_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_333to380_bb3_c0_ene6_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_333to380_bb3_c0_ene6_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_333to380_bb3_c0_ene6_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_333to380_bb3_c0_ene6_0_reg_380_fifo.DEPTH = 47;
defparam rnode_333to380_bb3_c0_ene6_0_reg_380_fifo.DATA_WIDTH = 32;
defparam rnode_333to380_bb3_c0_ene6_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to380_bb3_c0_ene6_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_333to380_bb3_c0_ene6_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to380_bb3_c0_ene6_0_NO_SHIFT_REG = rnode_333to380_bb3_c0_ene6_0_reg_380_NO_SHIFT_REG;
assign rnode_333to380_bb3_c0_ene6_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_333to380_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 54
//  * capacity = 54
 logic rnode_333to387_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to387_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_333to387_bb3_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_333to387_bb3_c0_ene7_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_333to387_bb3_c0_ene7_0_reg_387_NO_SHIFT_REG;
 logic rnode_333to387_bb3_c0_ene7_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_333to387_bb3_c0_ene7_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_333to387_bb3_c0_ene7_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_333to387_bb3_c0_ene7_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to387_bb3_c0_ene7_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to387_bb3_c0_ene7_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_333to387_bb3_c0_ene7_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_333to387_bb3_c0_ene7_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3_c0_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_333to387_bb3_c0_ene7_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_333to387_bb3_c0_ene7_0_reg_387_fifo.DEPTH = 54;
defparam rnode_333to387_bb3_c0_ene7_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_333to387_bb3_c0_ene7_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to387_bb3_c0_ene7_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_333to387_bb3_c0_ene7_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to387_bb3_c0_ene7_0_NO_SHIFT_REG = rnode_333to387_bb3_c0_ene7_0_reg_387_NO_SHIFT_REG;
assign rnode_333to387_bb3_c0_ene7_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_333to387_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_333_334_0_inputs_ready;
 reg SFC_1_VALID_333_334_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_333_334_0_stall_in;
wire SFC_1_VALID_333_334_0_output_regs_ready;
 reg SFC_1_VALID_333_334_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_333_334_0_causedstall;

assign SFC_1_VALID_333_334_0_inputs_ready = 1'b1;
assign SFC_1_VALID_333_334_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_332_333_0_stall_in = 1'b0;
assign SFC_1_VALID_333_334_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_333_334_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_333_334_0_output_regs_ready)
		begin
			SFC_1_VALID_333_334_0_NO_SHIFT_REG <= SFC_1_VALID_332_333_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_shr3_i500_stall_local;
wire [31:0] local_bb3_shr3_i500;

assign local_bb3_shr3_i500 = ((local_bb3_and2_i499 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and_i497_stall_local;
wire [31:0] local_bb3_and_i497;

assign local_bb3_and_i497 = (local_bb3_xor_i496 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and10_i503_stall_local;
wire [31:0] local_bb3_and10_i503;

assign local_bb3_and10_i503 = (local_bb3_xor_i496 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and_i313_stall_local;
wire [31:0] local_bb3_and_i313;

assign local_bb3_and_i313 = ((local_bb3_shr_i312 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_i324_stall_local;
wire local_bb3_lnot14_i324;

assign local_bb3_lnot14_i324 = ((local_bb3_and5_i318 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i346_stall_local;
wire [31:0] local_bb3_or_i346;

assign local_bb3_or_i346 = ((local_bb3_and5_i318 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_and3_i315_stall_local;
wire [31:0] local_bb3_and3_i315;

assign local_bb3_and3_i315 = ((local_bb3_shr2_i314 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_i325_stall_local;
wire local_bb3_lnot17_i325;

assign local_bb3_lnot17_i325 = ((local_bb3_and6_i319 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or47_i347_stall_local;
wire [31:0] local_bb3_or47_i347;

assign local_bb3_or47_i347 = ((local_bb3_and6_i319 & 32'h7FFFFF) | 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb3_c0_ene5_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_c0_ene5_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_c0_ene5_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3_c0_ene5_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_c0_ene5_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3_c0_ene5_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_c0_ene5_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_c0_ene5_0_valid_out_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_c0_ene5_0_stall_in_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_c0_ene5_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb3_c0_ene5_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb3_c0_ene5_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb3_c0_ene5_0_stall_in_0_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb3_c0_ene5_0_valid_out_0_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb3_c0_ene5_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in(rnode_333to385_bb3_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_385to386_bb3_c0_ene5_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb3_c0_ene5_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb3_c0_ene5_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_385to386_bb3_c0_ene5_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb3_c0_ene5_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb3_c0_ene5_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to385_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_c0_ene5_0_stall_in_0_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_c0_ene5_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_c0_ene5_0_NO_SHIFT_REG = rnode_385to386_bb3_c0_ene5_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_c0_ene5_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_c0_ene5_1_NO_SHIFT_REG = rnode_385to386_bb3_c0_ene5_0_reg_386_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_380to381_bb3_c0_ene6_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_c0_ene6_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_c0_ene6_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_380to381_bb3_c0_ene6_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_c0_ene6_1_NO_SHIFT_REG;
 logic rnode_380to381_bb3_c0_ene6_0_reg_381_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_c0_ene6_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_c0_ene6_0_valid_out_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_c0_ene6_0_stall_in_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_c0_ene6_0_stall_out_reg_381_NO_SHIFT_REG;

acl_data_fifo rnode_380to381_bb3_c0_ene6_0_reg_381_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_380to381_bb3_c0_ene6_0_reg_381_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_380to381_bb3_c0_ene6_0_stall_in_0_reg_381_NO_SHIFT_REG),
	.valid_out(rnode_380to381_bb3_c0_ene6_0_valid_out_0_reg_381_NO_SHIFT_REG),
	.stall_out(rnode_380to381_bb3_c0_ene6_0_stall_out_reg_381_NO_SHIFT_REG),
	.data_in(rnode_333to380_bb3_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_380to381_bb3_c0_ene6_0_reg_381_NO_SHIFT_REG)
);

defparam rnode_380to381_bb3_c0_ene6_0_reg_381_fifo.DEPTH = 1;
defparam rnode_380to381_bb3_c0_ene6_0_reg_381_fifo.DATA_WIDTH = 32;
defparam rnode_380to381_bb3_c0_ene6_0_reg_381_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_380to381_bb3_c0_ene6_0_reg_381_fifo.IMPL = "shift_reg";

assign rnode_380to381_bb3_c0_ene6_0_reg_381_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to380_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_c0_ene6_0_stall_in_0_reg_381_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_c0_ene6_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_380to381_bb3_c0_ene6_0_NO_SHIFT_REG = rnode_380to381_bb3_c0_ene6_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_c0_ene6_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_380to381_bb3_c0_ene6_1_NO_SHIFT_REG = rnode_380to381_bb3_c0_ene6_0_reg_381_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_c0_ene7_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene7_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_c0_ene7_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_c0_ene7_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_c0_ene7_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_c0_ene7_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_c0_ene7_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_333to387_bb3_c0_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb3_c0_ene7_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_c0_ene7_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_c0_ene7_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb3_c0_ene7_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_c0_ene7_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_c0_ene7_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to387_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_c0_ene7_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_c0_ene7_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_c0_ene7_0_NO_SHIFT_REG = rnode_387to388_bb3_c0_ene7_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_c0_ene7_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_c0_ene7_1_NO_SHIFT_REG = rnode_387to388_bb3_c0_ene7_0_reg_388_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_1_VALID_334_335_0_inputs_ready;
 reg SFC_1_VALID_334_335_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_334_335_0_stall_in;
wire SFC_1_VALID_334_335_0_output_regs_ready;
 reg SFC_1_VALID_334_335_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_334_335_0_causedstall;

assign SFC_1_VALID_334_335_0_inputs_ready = 1'b1;
assign SFC_1_VALID_334_335_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_333_334_0_stall_in = 1'b0;
assign SFC_1_VALID_334_335_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_334_335_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_334_335_0_output_regs_ready)
		begin
			SFC_1_VALID_334_335_0_NO_SHIFT_REG <= SFC_1_VALID_333_334_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_shr_i498_stall_local;
wire [31:0] local_bb3_shr_i498;

assign local_bb3_shr_i498 = ((local_bb3_and_i497 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp13_i505_stall_local;
wire local_bb3_cmp13_i505;

assign local_bb3_cmp13_i505 = ((local_bb3_and10_i503 & 32'hFFFF) > (local_bb3_and12_i504 & 32'hFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_i320_stall_local;
wire local_bb3_lnot_i320;

assign local_bb3_lnot_i320 = ((local_bb3_and_i313 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i322_stall_local;
wire local_bb3_cmp_i322;

assign local_bb3_cmp_i322 = ((local_bb3_and_i313 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u18_stall_local;
wire [31:0] local_bb3_var__u18;

assign local_bb3_var__u18 = ((local_bb3_and6_i319 & 32'h7FFFFF) | (local_bb3_and_i313 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_not_i343_stall_local;
wire local_bb3_lnot14_not_i343;

assign local_bb3_lnot14_not_i343 = (local_bb3_lnot14_i324 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_conv_i_i348_stall_local;
wire [63:0] local_bb3_conv_i_i348;

assign local_bb3_conv_i_i348[63:32] = 32'h0;
assign local_bb3_conv_i_i348[31:0] = ((local_bb3_or_i346 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot8_i321_stall_local;
wire local_bb3_lnot8_i321;

assign local_bb3_lnot8_i321 = ((local_bb3_and3_i315 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_i323_stall_local;
wire local_bb3_cmp11_i323;

assign local_bb3_cmp11_i323 = ((local_bb3_and3_i315 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u19_stall_local;
wire [31:0] local_bb3_var__u19;

assign local_bb3_var__u19 = ((local_bb3_and3_i315 & 32'hFF) | (local_bb3_and6_i319 & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_add_i357_stall_local;
wire [31:0] local_bb3_add_i357;

assign local_bb3_add_i357 = ((local_bb3_and3_i315 & 32'hFF) + (local_bb3_and_i313 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_not_i329_stall_local;
wire local_bb3_lnot17_not_i329;

assign local_bb3_lnot17_not_i329 = (local_bb3_lnot17_i325 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_conv1_i_i349_stall_local;
wire [63:0] local_bb3_conv1_i_i349;

assign local_bb3_conv1_i_i349[63:32] = 32'h0;
assign local_bb3_conv1_i_i349[31:0] = ((local_bb3_or47_i347 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u20_stall_local;
wire [31:0] local_bb3_var__u20;

assign local_bb3_var__u20 = rnode_385to386_bb3_c0_ene5_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to387_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_c0_ene5_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_c0_ene5_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_c0_ene5_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_c0_ene5_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_c0_ene5_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_c0_ene5_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_c0_ene5_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_c0_ene5_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_c0_ene5_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_c0_ene5_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_385to386_bb3_c0_ene5_1_NO_SHIFT_REG),
	.data_out(rnode_386to387_bb3_c0_ene5_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_c0_ene5_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_c0_ene5_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb3_c0_ene5_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_c0_ene5_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_c0_ene5_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_c0_ene5_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_c0_ene5_0_NO_SHIFT_REG = rnode_386to387_bb3_c0_ene5_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_c0_ene5_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u21_stall_local;
wire [31:0] local_bb3_var__u21;

assign local_bb3_var__u21 = rnode_380to381_bb3_c0_ene6_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_381to382_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_381to382_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3_c0_ene6_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_c0_ene6_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_c0_ene6_0_valid_out_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_c0_ene6_0_stall_in_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_c0_ene6_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_381to382_bb3_c0_ene6_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to382_bb3_c0_ene6_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to382_bb3_c0_ene6_0_stall_in_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_381to382_bb3_c0_ene6_0_valid_out_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_381to382_bb3_c0_ene6_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(rnode_380to381_bb3_c0_ene6_1_NO_SHIFT_REG),
	.data_out(rnode_381to382_bb3_c0_ene6_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_381to382_bb3_c0_ene6_0_reg_382_fifo.DEPTH = 1;
defparam rnode_381to382_bb3_c0_ene6_0_reg_382_fifo.DATA_WIDTH = 32;
defparam rnode_381to382_bb3_c0_ene6_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to382_bb3_c0_ene6_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_381to382_bb3_c0_ene6_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_380to381_bb3_c0_ene6_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_c0_ene6_0_NO_SHIFT_REG = rnode_381to382_bb3_c0_ene6_0_reg_382_NO_SHIFT_REG;
assign rnode_381to382_bb3_c0_ene6_0_stall_in_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_388to389_bb3_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_c0_ene7_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic rnode_388to389_bb3_c0_ene7_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_c0_ene7_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_c0_ene7_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_c0_ene7_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3_c0_ene7_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3_c0_ene7_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3_c0_ene7_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3_c0_ene7_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3_c0_ene7_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(rnode_387to388_bb3_c0_ene7_1_NO_SHIFT_REG),
	.data_out(rnode_388to389_bb3_c0_ene7_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3_c0_ene7_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3_c0_ene7_0_reg_389_fifo.DATA_WIDTH = 1;
defparam rnode_388to389_bb3_c0_ene7_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3_c0_ene7_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3_c0_ene7_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_c0_ene7_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_c0_ene7_0_NO_SHIFT_REG = rnode_388to389_bb3_c0_ene7_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3_c0_ene7_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_335_336_0_inputs_ready;
 reg SFC_1_VALID_335_336_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_335_336_0_stall_in;
wire SFC_1_VALID_335_336_0_output_regs_ready;
 reg SFC_1_VALID_335_336_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_335_336_0_causedstall;

assign SFC_1_VALID_335_336_0_inputs_ready = 1'b1;
assign SFC_1_VALID_335_336_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_334_335_0_stall_in = 1'b0;
assign SFC_1_VALID_335_336_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_335_336_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_335_336_0_output_regs_ready)
		begin
			SFC_1_VALID_335_336_0_NO_SHIFT_REG <= SFC_1_VALID_334_335_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i501_stall_local;
wire local_bb3_cmp_i501;

assign local_bb3_cmp_i501 = ((local_bb3_shr_i498 & 32'h7FFF) > (local_bb3_shr3_i500 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp8_i502_stall_local;
wire local_bb3_cmp8_i502;

assign local_bb3_cmp8_i502 = ((local_bb3_shr_i498 & 32'h7FFF) == (local_bb3_shr3_i500 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u22_stall_local;
wire local_bb3_var__u22;

assign local_bb3_var__u22 = ((local_bb3_var__u18 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__28_i344_stall_local;
wire local_bb3__28_i344;

assign local_bb3__28_i344 = (local_bb3_cmp_i322 & local_bb3_lnot14_not_i343);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_0_i375_stall_local;
wire local_bb3_reduction_0_i375;

assign local_bb3_reduction_0_i375 = (local_bb3_lnot_i320 | local_bb3_lnot8_i321);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge8_demorgan_i326_stall_local;
wire local_bb3_brmerge8_demorgan_i326;

assign local_bb3_brmerge8_demorgan_i326 = (local_bb3_cmp11_i323 & local_bb3_lnot17_i325);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_not_i330_stall_local;
wire local_bb3_cmp11_not_i330;

assign local_bb3_cmp11_not_i330 = (local_bb3_cmp11_i323 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u23_stall_local;
wire local_bb3_var__u23;

assign local_bb3_var__u23 = (local_bb3_cmp_i322 | local_bb3_cmp11_i323);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u24_stall_local;
wire local_bb3_var__u24;

assign local_bb3_var__u24 = ((local_bb3_var__u19 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and2_i13_stall_local;
wire [31:0] local_bb3_and2_i13;

assign local_bb3_and2_i13 = (local_bb3_var__u20 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and12_i18_stall_local;
wire [31:0] local_bb3_and12_i18;

assign local_bb3_and12_i18 = (local_bb3_var__u20 & 32'hFFFF);

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_387to392_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to392_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to392_bb3_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_387to392_bb3_c0_ene5_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to392_bb3_c0_ene5_0_reg_392_NO_SHIFT_REG;
 logic rnode_387to392_bb3_c0_ene5_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_387to392_bb3_c0_ene5_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_387to392_bb3_c0_ene5_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_387to392_bb3_c0_ene5_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to392_bb3_c0_ene5_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to392_bb3_c0_ene5_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_387to392_bb3_c0_ene5_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_387to392_bb3_c0_ene5_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_386to387_bb3_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_387to392_bb3_c0_ene5_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_387to392_bb3_c0_ene5_0_reg_392_fifo.DEPTH = 5;
defparam rnode_387to392_bb3_c0_ene5_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_387to392_bb3_c0_ene5_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to392_bb3_c0_ene5_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_387to392_bb3_c0_ene5_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to392_bb3_c0_ene5_0_NO_SHIFT_REG = rnode_387to392_bb3_c0_ene5_0_reg_392_NO_SHIFT_REG;
assign rnode_387to392_bb3_c0_ene5_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_387to392_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and2_i2_stall_local;
wire [31:0] local_bb3_and2_i2;

assign local_bb3_and2_i2 = (local_bb3_var__u21 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and12_i_stall_local;
wire [31:0] local_bb3_and12_i;

assign local_bb3_and12_i = (local_bb3_var__u21 & 32'hFFFF);

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_382to387_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_382to387_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_382to387_bb3_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_382to387_bb3_c0_ene6_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_382to387_bb3_c0_ene6_0_reg_387_NO_SHIFT_REG;
 logic rnode_382to387_bb3_c0_ene6_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_382to387_bb3_c0_ene6_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_382to387_bb3_c0_ene6_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_382to387_bb3_c0_ene6_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to387_bb3_c0_ene6_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to387_bb3_c0_ene6_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_382to387_bb3_c0_ene6_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_382to387_bb3_c0_ene6_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_381to382_bb3_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_382to387_bb3_c0_ene6_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_382to387_bb3_c0_ene6_0_reg_387_fifo.DEPTH = 5;
defparam rnode_382to387_bb3_c0_ene6_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_382to387_bb3_c0_ene6_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to387_bb3_c0_ene6_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_382to387_bb3_c0_ene6_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_382to387_bb3_c0_ene6_0_NO_SHIFT_REG = rnode_382to387_bb3_c0_ene6_0_reg_387_NO_SHIFT_REG;
assign rnode_382to387_bb3_c0_ene6_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_382to387_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_389to392_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to392_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_389to392_bb3_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_389to392_bb3_c0_ene7_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to392_bb3_c0_ene7_0_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb3_c0_ene7_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb3_c0_ene7_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb3_c0_ene7_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_389to392_bb3_c0_ene7_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to392_bb3_c0_ene7_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to392_bb3_c0_ene7_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_389to392_bb3_c0_ene7_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_389to392_bb3_c0_ene7_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_388to389_bb3_c0_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_389to392_bb3_c0_ene7_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_389to392_bb3_c0_ene7_0_reg_392_fifo.DEPTH = 3;
defparam rnode_389to392_bb3_c0_ene7_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_389to392_bb3_c0_ene7_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to392_bb3_c0_ene7_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_389to392_bb3_c0_ene7_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_389to392_bb3_c0_ene7_0_NO_SHIFT_REG = rnode_389to392_bb3_c0_ene7_0_reg_392_NO_SHIFT_REG;
assign rnode_389to392_bb3_c0_ene7_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_389to392_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_336_337_0_inputs_ready;
 reg SFC_1_VALID_336_337_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_336_337_0_stall_in;
wire SFC_1_VALID_336_337_0_output_regs_ready;
 reg SFC_1_VALID_336_337_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_336_337_0_causedstall;

assign SFC_1_VALID_336_337_0_inputs_ready = 1'b1;
assign SFC_1_VALID_336_337_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_335_336_0_stall_in = 1'b0;
assign SFC_1_VALID_336_337_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_336_337_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_336_337_0_output_regs_ready)
		begin
			SFC_1_VALID_336_337_0_NO_SHIFT_REG <= SFC_1_VALID_335_336_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3___i506_stall_local;
wire local_bb3___i506;

assign local_bb3___i506 = (local_bb3_cmp8_i502 & local_bb3_cmp13_i505);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge10_demorgan_i327_stall_local;
wire local_bb3_brmerge10_demorgan_i327;

assign local_bb3_brmerge10_demorgan_i327 = (local_bb3_brmerge8_demorgan_i326 & local_bb3_lnot_i320);

// This section implements an unregistered operation.
// 
wire local_bb3__mux9_mux_i328_stall_local;
wire local_bb3__mux9_mux_i328;

assign local_bb3__mux9_mux_i328 = (local_bb3_brmerge8_demorgan_i326 ^ local_bb3_cmp11_i323);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge3_i331_stall_local;
wire local_bb3_brmerge3_i331;

assign local_bb3_brmerge3_i331 = (local_bb3_var__u24 | local_bb3_cmp11_not_i330);

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_i333_stall_local;
wire local_bb3__mux_mux_i333;

assign local_bb3__mux_mux_i333 = (local_bb3_var__u24 | local_bb3_cmp11_i323);

// This section implements an unregistered operation.
// 
wire local_bb3__not_i335_stall_local;
wire local_bb3__not_i335;

assign local_bb3__not_i335 = (local_bb3_var__u24 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_shr3_i14_stall_local;
wire [31:0] local_bb3_shr3_i14;

assign local_bb3_shr3_i14 = ((local_bb3_and2_i13 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb3_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene5_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb3_c0_ene5_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene5_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene5_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene5_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3_c0_ene5_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3_c0_ene5_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3_c0_ene5_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3_c0_ene5_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3_c0_ene5_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_387to392_bb3_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb3_c0_ene5_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3_c0_ene5_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3_c0_ene5_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_392to393_bb3_c0_ene5_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3_c0_ene5_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3_c0_ene5_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_387to392_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_c0_ene5_0_NO_SHIFT_REG = rnode_392to393_bb3_c0_ene5_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_c0_ene5_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr3_i_stall_local;
wire [31:0] local_bb3_shr3_i;

assign local_bb3_shr3_i = ((local_bb3_and2_i2 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene6_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_c0_ene6_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene6_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene6_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_c0_ene6_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_c0_ene6_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_c0_ene6_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_c0_ene6_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_c0_ene6_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_c0_ene6_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_382to387_bb3_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb3_c0_ene6_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_c0_ene6_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_c0_ene6_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb3_c0_ene6_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_c0_ene6_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_c0_ene6_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_382to387_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_c0_ene6_0_NO_SHIFT_REG = rnode_387to388_bb3_c0_ene6_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_c0_ene6_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene7_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene7_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene7_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene7_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_c0_ene7_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3_c0_ene7_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3_c0_ene7_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3_c0_ene7_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3_c0_ene7_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3_c0_ene7_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_389to392_bb3_c0_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb3_c0_ene7_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3_c0_ene7_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3_c0_ene7_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb3_c0_ene7_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3_c0_ene7_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3_c0_ene7_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to392_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_c0_ene7_0_NO_SHIFT_REG = rnode_392to393_bb3_c0_ene7_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_c0_ene7_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_337_338_0_inputs_ready;
 reg SFC_1_VALID_337_338_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_337_338_0_stall_in;
wire SFC_1_VALID_337_338_0_output_regs_ready;
 reg SFC_1_VALID_337_338_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_337_338_0_causedstall;

assign SFC_1_VALID_337_338_0_inputs_ready = 1'b1;
assign SFC_1_VALID_337_338_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_336_337_0_stall_in = 1'b0;
assign SFC_1_VALID_337_338_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_337_338_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_337_338_0_output_regs_ready)
		begin
			SFC_1_VALID_337_338_0_NO_SHIFT_REG <= SFC_1_VALID_336_337_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_valid_out_1;
wire local_bb3_c0_ene1_stall_in_1;
wire local_bb3_var__u14_valid_out_2;
wire local_bb3_var__u14_stall_in_2;
wire local_bb3_xor_i496_valid_out_2;
wire local_bb3_xor_i496_stall_in_2;
wire local_bb3__21_i507_valid_out;
wire local_bb3__21_i507_stall_in;
wire local_bb3__21_i507_inputs_ready;
wire local_bb3__21_i507_stall_local;
wire local_bb3__21_i507;

assign local_bb3__21_i507_inputs_ready = (local_bb3_c0_enter_c0_eni7_valid_out_0_NO_SHIFT_REG & local_bb3_c0_enter_c0_eni7_valid_out_1_NO_SHIFT_REG);
assign local_bb3__21_i507 = (local_bb3_cmp_i501 | local_bb3___i506);
assign local_bb3_c0_ene1_valid_out_1 = 1'b1;
assign local_bb3_var__u14_valid_out_2 = 1'b1;
assign local_bb3_xor_i496_valid_out_2 = 1'b1;
assign local_bb3__21_i507_valid_out = 1'b1;
assign local_bb3_c0_enter_c0_eni7_stall_in_0 = 1'b0;
assign local_bb3_c0_enter_c0_eni7_stall_in_1 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__26_demorgan_i341_stall_local;
wire local_bb3__26_demorgan_i341;

assign local_bb3__26_demorgan_i341 = (local_bb3_cmp_i322 | local_bb3_brmerge10_demorgan_i327);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge5_i332_stall_local;
wire local_bb3_brmerge5_i332;

assign local_bb3_brmerge5_i332 = (local_bb3_brmerge3_i331 | local_bb3_lnot17_not_i329);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_3_i336_stall_local;
wire local_bb3_reduction_3_i336;

assign local_bb3_reduction_3_i336 = (local_bb3_cmp11_i323 & local_bb3__not_i335);

// This section implements a registered operation.
// 
wire SFC_1_VALID_338_339_0_inputs_ready;
 reg SFC_1_VALID_338_339_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_338_339_0_stall_in;
wire SFC_1_VALID_338_339_0_output_regs_ready;
 reg SFC_1_VALID_338_339_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_338_339_0_causedstall;

assign SFC_1_VALID_338_339_0_inputs_ready = 1'b1;
assign SFC_1_VALID_338_339_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_337_338_0_stall_in = 1'b0;
assign SFC_1_VALID_338_339_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_338_339_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_338_339_0_output_regs_ready)
		begin
			SFC_1_VALID_338_339_0_NO_SHIFT_REG <= SFC_1_VALID_337_338_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene1_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_c0_ene1_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene1_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene1_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_c0_ene1_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_c0_ene1_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_c0_ene1_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_c0_ene1_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_c0_ene1_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_c0_ene1_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene1),
	.data_out(rnode_332to333_bb3_c0_ene1_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_c0_ene1_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_c0_ene1_0_reg_333_fifo.DATA_WIDTH = 32;
defparam rnode_332to333_bb3_c0_ene1_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_c0_ene1_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_c0_ene1_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene1_stall_in_1 = 1'b0;
assign rnode_332to333_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_332to333_bb3_c0_ene1_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_c0_ene1_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_var__u14_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u14_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_var__u14_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u14_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u14_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_var__u14_1_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u14_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_var__u14_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u14_0_valid_out_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u14_0_stall_in_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u14_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_var__u14_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_var__u14_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_var__u14_0_stall_in_0_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_var__u14_0_valid_out_0_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_var__u14_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_var__u14),
	.data_out(rnode_332to333_bb3_var__u14_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_var__u14_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_var__u14_0_reg_333_fifo.DATA_WIDTH = 32;
defparam rnode_332to333_bb3_var__u14_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_var__u14_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_var__u14_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u14_stall_in_2 = 1'b0;
assign rnode_332to333_bb3_var__u14_0_stall_in_0_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_var__u14_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_var__u14_0_NO_SHIFT_REG = rnode_332to333_bb3_var__u14_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_var__u14_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_var__u14_1_NO_SHIFT_REG = rnode_332to333_bb3_var__u14_0_reg_333_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_xor_i496_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i496_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_xor_i496_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i496_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i496_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_xor_i496_1_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i496_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_xor_i496_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i496_0_valid_out_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i496_0_stall_in_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i496_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_xor_i496_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_xor_i496_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_xor_i496_0_stall_in_0_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_xor_i496_0_valid_out_0_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_xor_i496_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_xor_i496),
	.data_out(rnode_332to333_bb3_xor_i496_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_xor_i496_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_xor_i496_0_reg_333_fifo.DATA_WIDTH = 32;
defparam rnode_332to333_bb3_xor_i496_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_xor_i496_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_xor_i496_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_xor_i496_stall_in_2 = 1'b0;
assign rnode_332to333_bb3_xor_i496_0_stall_in_0_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_xor_i496_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_xor_i496_0_NO_SHIFT_REG = rnode_332to333_bb3_xor_i496_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_xor_i496_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_xor_i496_1_NO_SHIFT_REG = rnode_332to333_bb3_xor_i496_0_reg_333_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3__21_i507_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_1_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_valid_out_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_stall_in_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3__21_i507_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3__21_i507_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3__21_i507_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3__21_i507_0_stall_in_0_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3__21_i507_0_valid_out_0_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3__21_i507_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3__21_i507),
	.data_out(rnode_332to333_bb3__21_i507_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3__21_i507_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3__21_i507_0_reg_333_fifo.DATA_WIDTH = 1;
defparam rnode_332to333_bb3__21_i507_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3__21_i507_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3__21_i507_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__21_i507_stall_in = 1'b0;
assign rnode_332to333_bb3__21_i507_0_stall_in_0_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3__21_i507_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3__21_i507_0_NO_SHIFT_REG = rnode_332to333_bb3__21_i507_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3__21_i507_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3__21_i507_1_NO_SHIFT_REG = rnode_332to333_bb3__21_i507_0_reg_333_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_mux_i334_stall_local;
wire local_bb3__mux_mux_mux_i334;

assign local_bb3__mux_mux_mux_i334 = (local_bb3_brmerge5_i332 & local_bb3__mux_mux_i333);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_5_i337_stall_local;
wire local_bb3_reduction_5_i337;

assign local_bb3_reduction_5_i337 = (local_bb3_lnot14_i324 & local_bb3_reduction_3_i336);

// This section implements a registered operation.
// 
wire SFC_1_VALID_339_340_0_inputs_ready;
 reg SFC_1_VALID_339_340_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_339_340_0_stall_in;
wire SFC_1_VALID_339_340_0_output_regs_ready;
 reg SFC_1_VALID_339_340_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_339_340_0_causedstall;

assign SFC_1_VALID_339_340_0_inputs_ready = 1'b1;
assign SFC_1_VALID_339_340_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_338_339_0_stall_in = 1'b0;
assign SFC_1_VALID_339_340_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_339_340_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_339_340_0_output_regs_ready)
		begin
			SFC_1_VALID_339_340_0_NO_SHIFT_REG <= SFC_1_VALID_338_339_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 46
//  * capacity = 46
 logic rnode_333to379_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to379_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_333to379_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_333to379_bb3_c0_ene1_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to379_bb3_c0_ene1_0_reg_379_NO_SHIFT_REG;
 logic rnode_333to379_bb3_c0_ene1_0_valid_out_reg_379_NO_SHIFT_REG;
 logic rnode_333to379_bb3_c0_ene1_0_stall_in_reg_379_NO_SHIFT_REG;
 logic rnode_333to379_bb3_c0_ene1_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_333to379_bb3_c0_ene1_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to379_bb3_c0_ene1_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to379_bb3_c0_ene1_0_stall_in_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_333to379_bb3_c0_ene1_0_valid_out_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_333to379_bb3_c0_ene1_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3_c0_ene1_0_NO_SHIFT_REG),
	.data_out(rnode_333to379_bb3_c0_ene1_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_333to379_bb3_c0_ene1_0_reg_379_fifo.DEPTH = 46;
defparam rnode_333to379_bb3_c0_ene1_0_reg_379_fifo.DATA_WIDTH = 32;
defparam rnode_333to379_bb3_c0_ene1_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to379_bb3_c0_ene1_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_333to379_bb3_c0_ene1_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to379_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_333to379_bb3_c0_ene1_0_reg_379_NO_SHIFT_REG;
assign rnode_333to379_bb3_c0_ene1_0_stall_in_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_333to379_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__22_i508_stall_local;
wire [31:0] local_bb3__22_i508;

assign local_bb3__22_i508 = (rnode_332to333_bb3__21_i507_0_NO_SHIFT_REG ? rnode_332to333_bb3_var__u14_0_NO_SHIFT_REG : rnode_332to333_bb3_xor_i496_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3__23_i509_stall_local;
wire [31:0] local_bb3__23_i509;

assign local_bb3__23_i509 = (rnode_332to333_bb3__21_i507_1_NO_SHIFT_REG ? rnode_332to333_bb3_xor_i496_1_NO_SHIFT_REG : rnode_332to333_bb3_var__u14_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_6_i338_stall_local;
wire local_bb3_reduction_6_i338;

assign local_bb3_reduction_6_i338 = (local_bb3_var__u22 & local_bb3_reduction_5_i337);

// This section implements a registered operation.
// 
wire SFC_1_VALID_340_341_0_inputs_ready;
 reg SFC_1_VALID_340_341_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_340_341_0_stall_in;
wire SFC_1_VALID_340_341_0_output_regs_ready;
 reg SFC_1_VALID_340_341_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_340_341_0_causedstall;

assign SFC_1_VALID_340_341_0_inputs_ready = 1'b1;
assign SFC_1_VALID_340_341_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_339_340_0_stall_in = 1'b0;
assign SFC_1_VALID_340_341_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_340_341_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_340_341_0_output_regs_ready)
		begin
			SFC_1_VALID_340_341_0_NO_SHIFT_REG <= SFC_1_VALID_339_340_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_379to380_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_379to380_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_379to380_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_379to380_bb3_c0_ene1_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_379to380_bb3_c0_ene1_0_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_c0_ene1_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_c0_ene1_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_c0_ene1_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_379to380_bb3_c0_ene1_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_379to380_bb3_c0_ene1_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_379to380_bb3_c0_ene1_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_379to380_bb3_c0_ene1_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_379to380_bb3_c0_ene1_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(rnode_333to379_bb3_c0_ene1_0_NO_SHIFT_REG),
	.data_out(rnode_379to380_bb3_c0_ene1_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_379to380_bb3_c0_ene1_0_reg_380_fifo.DEPTH = 1;
defparam rnode_379to380_bb3_c0_ene1_0_reg_380_fifo.DATA_WIDTH = 32;
defparam rnode_379to380_bb3_c0_ene1_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_379to380_bb3_c0_ene1_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_379to380_bb3_c0_ene1_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to379_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_379to380_bb3_c0_ene1_0_reg_380_NO_SHIFT_REG;
assign rnode_379to380_bb3_c0_ene1_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr18_i512_stall_local;
wire [31:0] local_bb3_shr18_i512;

assign local_bb3_shr18_i512 = (local_bb3__22_i508 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shr16_i510_stall_local;
wire [31:0] local_bb3_shr16_i510;

assign local_bb3_shr16_i510 = (local_bb3__23_i509 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3__24_i339_stall_local;
wire local_bb3__24_i339;

assign local_bb3__24_i339 = (local_bb3_cmp_i322 ? local_bb3_reduction_6_i338 : local_bb3_brmerge10_demorgan_i327);

// This section implements a registered operation.
// 
wire SFC_1_VALID_341_342_0_inputs_ready;
 reg SFC_1_VALID_341_342_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_341_342_0_stall_in;
wire SFC_1_VALID_341_342_0_output_regs_ready;
 reg SFC_1_VALID_341_342_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_341_342_0_causedstall;

assign SFC_1_VALID_341_342_0_inputs_ready = 1'b1;
assign SFC_1_VALID_341_342_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_340_341_0_stall_in = 1'b0;
assign SFC_1_VALID_341_342_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_341_342_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_341_342_0_output_regs_ready)
		begin
			SFC_1_VALID_341_342_0_NO_SHIFT_REG <= SFC_1_VALID_340_341_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_var__u25_stall_local;
wire [31:0] local_bb3_var__u25;

assign local_bb3_var__u25 = rnode_379to380_bb3_c0_ene1_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_and19_i513_stall_local;
wire [31:0] local_bb3_and19_i513;

assign local_bb3_and19_i513 = ((local_bb3_shr18_i512 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_sub_i538_stall_local;
wire [31:0] local_bb3_sub_i538;

assign local_bb3_sub_i538 = ((local_bb3_shr16_i510 & 32'h1FF) - (local_bb3_shr18_i512 & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb3__25_i340_stall_local;
wire local_bb3__25_i340;

assign local_bb3__25_i340 = (local_bb3__24_i339 ? local_bb3_lnot14_i324 : local_bb3__mux_mux_mux_i334);

// This section implements a registered operation.
// 
wire SFC_1_VALID_342_343_0_inputs_ready;
 reg SFC_1_VALID_342_343_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_342_343_0_stall_in;
wire SFC_1_VALID_342_343_0_output_regs_ready;
 reg SFC_1_VALID_342_343_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_342_343_0_causedstall;

assign SFC_1_VALID_342_343_0_inputs_ready = 1'b1;
assign SFC_1_VALID_342_343_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_341_342_0_stall_in = 1'b0;
assign SFC_1_VALID_342_343_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_342_343_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_342_343_0_output_regs_ready)
		begin
			SFC_1_VALID_342_343_0_NO_SHIFT_REG <= SFC_1_VALID_341_342_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_shr2_i_stall_local;
wire [31:0] local_bb3_shr2_i;

assign local_bb3_shr2_i = (local_bb3_var__u25 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and6_i_stall_local;
wire [31:0] local_bb3_and6_i;

assign local_bb3_and6_i = (local_bb3_var__u25 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot23_i517_stall_local;
wire local_bb3_lnot23_i517;

assign local_bb3_lnot23_i517 = ((local_bb3_and19_i513 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp27_i519_stall_local;
wire local_bb3_cmp27_i519;

assign local_bb3_cmp27_i519 = ((local_bb3_and19_i513 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and69_i_stall_local;
wire [31:0] local_bb3_and69_i;

assign local_bb3_and69_i = (local_bb3_sub_i538 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3__27_i342_stall_local;
wire local_bb3__27_i342;

assign local_bb3__27_i342 = (local_bb3__26_demorgan_i341 ? local_bb3__25_i340 : local_bb3__mux9_mux_i328);

// This section implements a registered operation.
// 
wire SFC_1_VALID_343_344_0_inputs_ready;
 reg SFC_1_VALID_343_344_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_343_344_0_stall_in;
wire SFC_1_VALID_343_344_0_output_regs_ready;
 reg SFC_1_VALID_343_344_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_343_344_0_causedstall;

assign SFC_1_VALID_343_344_0_inputs_ready = 1'b1;
assign SFC_1_VALID_343_344_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_342_343_0_stall_in = 1'b0;
assign SFC_1_VALID_343_344_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_343_344_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_343_344_0_output_regs_ready)
		begin
			SFC_1_VALID_343_344_0_NO_SHIFT_REG <= SFC_1_VALID_342_343_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_or47_i_stall_local;
wire [31:0] local_bb3_or47_i;

assign local_bb3_or47_i = ((local_bb3_and6_i & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp70_i_stall_local;
wire local_bb3_cmp70_i;

assign local_bb3_cmp70_i = ((local_bb3_and69_i & 32'hFF) > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_xor_i316_valid_out;
wire local_bb3_xor_i316_stall_in;
wire local_bb3_add_i357_valid_out;
wire local_bb3_add_i357_stall_in;
wire local_bb3_conv_i_i348_valid_out;
wire local_bb3_conv_i_i348_stall_in;
wire local_bb3_conv1_i_i349_valid_out;
wire local_bb3_conv1_i_i349_stall_in;
wire local_bb3_reduction_0_i375_valid_out;
wire local_bb3_reduction_0_i375_stall_in;
wire local_bb3_var__u23_valid_out;
wire local_bb3_var__u23_stall_in;
wire local_bb3__29_i345_valid_out;
wire local_bb3__29_i345_stall_in;
wire local_bb3__29_i345_inputs_ready;
wire local_bb3__29_i345_stall_local;
wire local_bb3__29_i345;

assign local_bb3__29_i345_inputs_ready = (local_bb3_c0_enter_c0_eni7_valid_out_2_NO_SHIFT_REG & local_bb3_c0_enter_c0_eni7_valid_out_3_NO_SHIFT_REG);
assign local_bb3__29_i345 = (local_bb3__28_i344 | local_bb3__27_i342);
assign local_bb3_xor_i316_valid_out = 1'b1;
assign local_bb3_add_i357_valid_out = 1'b1;
assign local_bb3_conv_i_i348_valid_out = 1'b1;
assign local_bb3_conv1_i_i349_valid_out = 1'b1;
assign local_bb3_reduction_0_i375_valid_out = 1'b1;
assign local_bb3_var__u23_valid_out = 1'b1;
assign local_bb3__29_i345_valid_out = 1'b1;
assign local_bb3_c0_enter_c0_eni7_stall_in_2 = 1'b0;
assign local_bb3_c0_enter_c0_eni7_stall_in_3 = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_344_345_0_inputs_ready;
 reg SFC_1_VALID_344_345_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_344_345_0_stall_in;
wire SFC_1_VALID_344_345_0_output_regs_ready;
 reg SFC_1_VALID_344_345_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_344_345_0_causedstall;

assign SFC_1_VALID_344_345_0_inputs_ready = 1'b1;
assign SFC_1_VALID_344_345_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_343_344_0_stall_in = 1'b0;
assign SFC_1_VALID_344_345_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_344_345_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_344_345_0_output_regs_ready)
		begin
			SFC_1_VALID_344_345_0_NO_SHIFT_REG <= SFC_1_VALID_343_344_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_conv1_i_i_stall_local;
wire [63:0] local_bb3_conv1_i_i;

assign local_bb3_conv1_i_i[63:32] = 32'h0;
assign local_bb3_conv1_i_i[31:0] = ((local_bb3_or47_i & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3__22_i508_valid_out_1;
wire local_bb3__22_i508_stall_in_1;
wire local_bb3__23_i509_valid_out_1;
wire local_bb3__23_i509_stall_in_1;
wire local_bb3_shr16_i510_valid_out_1;
wire local_bb3_shr16_i510_stall_in_1;
wire local_bb3_lnot23_i517_valid_out;
wire local_bb3_lnot23_i517_stall_in;
wire local_bb3_cmp27_i519_valid_out;
wire local_bb3_cmp27_i519_stall_in;
wire local_bb3_align_0_i539_valid_out;
wire local_bb3_align_0_i539_stall_in;
wire local_bb3_align_0_i539_inputs_ready;
wire local_bb3_align_0_i539_stall_local;
wire [31:0] local_bb3_align_0_i539;

assign local_bb3_align_0_i539_inputs_ready = (rnode_332to333_bb3__21_i507_0_valid_out_0_NO_SHIFT_REG & rnode_332to333_bb3_var__u14_0_valid_out_0_NO_SHIFT_REG & rnode_332to333_bb3_xor_i496_0_valid_out_0_NO_SHIFT_REG & rnode_332to333_bb3__21_i507_0_valid_out_1_NO_SHIFT_REG & rnode_332to333_bb3_xor_i496_0_valid_out_1_NO_SHIFT_REG & rnode_332to333_bb3_var__u14_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_align_0_i539 = (local_bb3_cmp70_i ? 32'h1F : (local_bb3_and69_i & 32'hFF));
assign local_bb3__22_i508_valid_out_1 = 1'b1;
assign local_bb3__23_i509_valid_out_1 = 1'b1;
assign local_bb3_shr16_i510_valid_out_1 = 1'b1;
assign local_bb3_lnot23_i517_valid_out = 1'b1;
assign local_bb3_cmp27_i519_valid_out = 1'b1;
assign local_bb3_align_0_i539_valid_out = 1'b1;
assign rnode_332to333_bb3__21_i507_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_var__u14_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_xor_i496_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3__21_i507_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_xor_i496_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_var__u14_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_xor_i316_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i316_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_xor_i316_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i316_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_xor_i316_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i316_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i316_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_xor_i316_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_xor_i316_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_xor_i316_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_xor_i316_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_xor_i316_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_xor_i316_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_xor_i316),
	.data_out(rnode_332to333_bb3_xor_i316_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_xor_i316_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_xor_i316_0_reg_333_fifo.DATA_WIDTH = 32;
defparam rnode_332to333_bb3_xor_i316_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_xor_i316_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_xor_i316_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_xor_i316_stall_in = 1'b0;
assign rnode_332to333_bb3_xor_i316_0_NO_SHIFT_REG = rnode_332to333_bb3_xor_i316_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_xor_i316_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_xor_i316_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_add_i357_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_add_i357_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_add_i357_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_add_i357_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_332to333_bb3_add_i357_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_add_i357_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_add_i357_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_add_i357_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_add_i357_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_add_i357_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_add_i357_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_add_i357_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_add_i357_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in((local_bb3_add_i357 & 32'h1FF)),
	.data_out(rnode_332to333_bb3_add_i357_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_add_i357_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_add_i357_0_reg_333_fifo.DATA_WIDTH = 32;
defparam rnode_332to333_bb3_add_i357_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_add_i357_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_add_i357_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add_i357_stall_in = 1'b0;
assign rnode_332to333_bb3_add_i357_0_NO_SHIFT_REG = rnode_332to333_bb3_add_i357_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_add_i357_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_add_i357_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb3_mul_i_i350_inputs_ready;
 reg local_bb3_mul_i_i350_valid_out_0_NO_SHIFT_REG;
wire local_bb3_mul_i_i350_stall_in_0;
 reg local_bb3_mul_i_i350_valid_out_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i350_stall_in_1;
wire local_bb3_mul_i_i350_output_regs_ready;
wire [63:0] local_bb3_mul_i_i350;
 reg local_bb3_mul_i_i350_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_mul_i_i350_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i350_causedstall;

acl_int_mult int_module_local_bb3_mul_i_i350 (
	.clock(clock),
	.dataa(((local_bb3_conv1_i_i349 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb3_conv_i_i348 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb3_mul_i_i350_output_regs_ready),
	.result(local_bb3_mul_i_i350)
);

defparam int_module_local_bb3_mul_i_i350.INPUT1_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i350.INPUT2_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i350.OUTPUT_WIDTH = 64;
defparam int_module_local_bb3_mul_i_i350.LATENCY = 3;
defparam int_module_local_bb3_mul_i_i350.SIGNED = 0;

assign local_bb3_mul_i_i350_inputs_ready = 1'b1;
assign local_bb3_mul_i_i350_output_regs_ready = 1'b1;
assign local_bb3_conv1_i_i349_stall_in = 1'b0;
assign local_bb3_conv_i_i348_stall_in = 1'b0;
assign local_bb3_mul_i_i350_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i350_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i350_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i350_output_regs_ready)
		begin
			local_bb3_mul_i_i350_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i350_valid_pipe_1_NO_SHIFT_REG <= local_bb3_mul_i_i350_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i350_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i350_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i350_output_regs_ready)
		begin
			local_bb3_mul_i_i350_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i350_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_mul_i_i350_stall_in_0))
			begin
				local_bb3_mul_i_i350_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_mul_i_i350_stall_in_1))
			begin
				local_bb3_mul_i_i350_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_reduction_0_i375_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_reduction_0_i375_0_stall_in_NO_SHIFT_REG;
 logic rnode_332to333_bb3_reduction_0_i375_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_reduction_0_i375_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic rnode_332to333_bb3_reduction_0_i375_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_reduction_0_i375_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_reduction_0_i375_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_reduction_0_i375_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_reduction_0_i375_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_reduction_0_i375_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_reduction_0_i375_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_reduction_0_i375_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_reduction_0_i375_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_reduction_0_i375),
	.data_out(rnode_332to333_bb3_reduction_0_i375_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_reduction_0_i375_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_reduction_0_i375_0_reg_333_fifo.DATA_WIDTH = 1;
defparam rnode_332to333_bb3_reduction_0_i375_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_reduction_0_i375_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_reduction_0_i375_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_reduction_0_i375_stall_in = 1'b0;
assign rnode_332to333_bb3_reduction_0_i375_0_NO_SHIFT_REG = rnode_332to333_bb3_reduction_0_i375_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_reduction_0_i375_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_reduction_0_i375_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3_var__u23_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u23_0_stall_in_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u23_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u23_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u23_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u23_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u23_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3_var__u23_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3_var__u23_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3_var__u23_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3_var__u23_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3_var__u23_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3_var__u23_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3_var__u23),
	.data_out(rnode_332to333_bb3_var__u23_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3_var__u23_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3_var__u23_0_reg_333_fifo.DATA_WIDTH = 1;
defparam rnode_332to333_bb3_var__u23_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3_var__u23_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3_var__u23_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u23_stall_in = 1'b0;
assign rnode_332to333_bb3_var__u23_0_NO_SHIFT_REG = rnode_332to333_bb3_var__u23_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3_var__u23_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3_var__u23_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_332to333_bb3__29_i345_0_valid_out_NO_SHIFT_REG;
 logic rnode_332to333_bb3__29_i345_0_stall_in_NO_SHIFT_REG;
 logic rnode_332to333_bb3__29_i345_0_NO_SHIFT_REG;
 logic rnode_332to333_bb3__29_i345_0_reg_333_inputs_ready_NO_SHIFT_REG;
 logic rnode_332to333_bb3__29_i345_0_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3__29_i345_0_valid_out_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3__29_i345_0_stall_in_reg_333_NO_SHIFT_REG;
 logic rnode_332to333_bb3__29_i345_0_stall_out_reg_333_NO_SHIFT_REG;

acl_data_fifo rnode_332to333_bb3__29_i345_0_reg_333_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_332to333_bb3__29_i345_0_reg_333_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_332to333_bb3__29_i345_0_stall_in_reg_333_NO_SHIFT_REG),
	.valid_out(rnode_332to333_bb3__29_i345_0_valid_out_reg_333_NO_SHIFT_REG),
	.stall_out(rnode_332to333_bb3__29_i345_0_stall_out_reg_333_NO_SHIFT_REG),
	.data_in(local_bb3__29_i345),
	.data_out(rnode_332to333_bb3__29_i345_0_reg_333_NO_SHIFT_REG)
);

defparam rnode_332to333_bb3__29_i345_0_reg_333_fifo.DEPTH = 1;
defparam rnode_332to333_bb3__29_i345_0_reg_333_fifo.DATA_WIDTH = 1;
defparam rnode_332to333_bb3__29_i345_0_reg_333_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_332to333_bb3__29_i345_0_reg_333_fifo.IMPL = "shift_reg";

assign rnode_332to333_bb3__29_i345_0_reg_333_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__29_i345_stall_in = 1'b0;
assign rnode_332to333_bb3__29_i345_0_NO_SHIFT_REG = rnode_332to333_bb3__29_i345_0_reg_333_NO_SHIFT_REG;
assign rnode_332to333_bb3__29_i345_0_stall_in_reg_333_NO_SHIFT_REG = 1'b0;
assign rnode_332to333_bb3__29_i345_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_345_346_0_inputs_ready;
 reg SFC_1_VALID_345_346_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_345_346_0_stall_in;
wire SFC_1_VALID_345_346_0_output_regs_ready;
 reg SFC_1_VALID_345_346_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_345_346_0_causedstall;

assign SFC_1_VALID_345_346_0_inputs_ready = 1'b1;
assign SFC_1_VALID_345_346_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_344_345_0_stall_in = 1'b0;
assign SFC_1_VALID_345_346_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_345_346_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_345_346_0_output_regs_ready)
		begin
			SFC_1_VALID_345_346_0_NO_SHIFT_REG <= SFC_1_VALID_344_345_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_333to334_bb3__22_i508_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3__22_i508_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3__22_i508_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3__22_i508_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_333to334_bb3__22_i508_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3__22_i508_1_NO_SHIFT_REG;
 logic rnode_333to334_bb3__22_i508_0_reg_334_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3__22_i508_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3__22_i508_0_valid_out_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3__22_i508_0_stall_in_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3__22_i508_0_stall_out_reg_334_NO_SHIFT_REG;

acl_data_fifo rnode_333to334_bb3__22_i508_0_reg_334_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to334_bb3__22_i508_0_reg_334_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to334_bb3__22_i508_0_stall_in_0_reg_334_NO_SHIFT_REG),
	.valid_out(rnode_333to334_bb3__22_i508_0_valid_out_0_reg_334_NO_SHIFT_REG),
	.stall_out(rnode_333to334_bb3__22_i508_0_stall_out_reg_334_NO_SHIFT_REG),
	.data_in(local_bb3__22_i508),
	.data_out(rnode_333to334_bb3__22_i508_0_reg_334_NO_SHIFT_REG)
);

defparam rnode_333to334_bb3__22_i508_0_reg_334_fifo.DEPTH = 1;
defparam rnode_333to334_bb3__22_i508_0_reg_334_fifo.DATA_WIDTH = 32;
defparam rnode_333to334_bb3__22_i508_0_reg_334_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to334_bb3__22_i508_0_reg_334_fifo.IMPL = "shift_reg";

assign rnode_333to334_bb3__22_i508_0_reg_334_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__22_i508_stall_in_1 = 1'b0;
assign rnode_333to334_bb3__22_i508_0_stall_in_0_reg_334_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3__22_i508_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3__22_i508_0_NO_SHIFT_REG = rnode_333to334_bb3__22_i508_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3__22_i508_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3__22_i508_1_NO_SHIFT_REG = rnode_333to334_bb3__22_i508_0_reg_334_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_333to334_bb3__23_i509_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3__23_i509_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3__23_i509_1_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3__23_i509_2_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_reg_334_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3__23_i509_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_valid_out_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_stall_in_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3__23_i509_0_stall_out_reg_334_NO_SHIFT_REG;

acl_data_fifo rnode_333to334_bb3__23_i509_0_reg_334_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to334_bb3__23_i509_0_reg_334_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to334_bb3__23_i509_0_stall_in_0_reg_334_NO_SHIFT_REG),
	.valid_out(rnode_333to334_bb3__23_i509_0_valid_out_0_reg_334_NO_SHIFT_REG),
	.stall_out(rnode_333to334_bb3__23_i509_0_stall_out_reg_334_NO_SHIFT_REG),
	.data_in(local_bb3__23_i509),
	.data_out(rnode_333to334_bb3__23_i509_0_reg_334_NO_SHIFT_REG)
);

defparam rnode_333to334_bb3__23_i509_0_reg_334_fifo.DEPTH = 1;
defparam rnode_333to334_bb3__23_i509_0_reg_334_fifo.DATA_WIDTH = 32;
defparam rnode_333to334_bb3__23_i509_0_reg_334_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to334_bb3__23_i509_0_reg_334_fifo.IMPL = "shift_reg";

assign rnode_333to334_bb3__23_i509_0_reg_334_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__23_i509_stall_in_1 = 1'b0;
assign rnode_333to334_bb3__23_i509_0_stall_in_0_reg_334_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3__23_i509_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3__23_i509_0_NO_SHIFT_REG = rnode_333to334_bb3__23_i509_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3__23_i509_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3__23_i509_1_NO_SHIFT_REG = rnode_333to334_bb3__23_i509_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3__23_i509_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3__23_i509_2_NO_SHIFT_REG = rnode_333to334_bb3__23_i509_0_reg_334_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_333to335_bb3_shr16_i510_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_333to335_bb3_shr16_i510_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_333to335_bb3_shr16_i510_0_NO_SHIFT_REG;
 logic rnode_333to335_bb3_shr16_i510_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_333to335_bb3_shr16_i510_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_333to335_bb3_shr16_i510_1_NO_SHIFT_REG;
 logic rnode_333to335_bb3_shr16_i510_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to335_bb3_shr16_i510_0_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_shr16_i510_0_valid_out_0_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_shr16_i510_0_stall_in_0_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_shr16_i510_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_333to335_bb3_shr16_i510_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to335_bb3_shr16_i510_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to335_bb3_shr16_i510_0_stall_in_0_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_333to335_bb3_shr16_i510_0_valid_out_0_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_333to335_bb3_shr16_i510_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in((local_bb3_shr16_i510 & 32'h1FF)),
	.data_out(rnode_333to335_bb3_shr16_i510_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_333to335_bb3_shr16_i510_0_reg_335_fifo.DEPTH = 2;
defparam rnode_333to335_bb3_shr16_i510_0_reg_335_fifo.DATA_WIDTH = 32;
defparam rnode_333to335_bb3_shr16_i510_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to335_bb3_shr16_i510_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_333to335_bb3_shr16_i510_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr16_i510_stall_in_1 = 1'b0;
assign rnode_333to335_bb3_shr16_i510_0_stall_in_0_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_333to335_bb3_shr16_i510_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_333to335_bb3_shr16_i510_0_NO_SHIFT_REG = rnode_333to335_bb3_shr16_i510_0_reg_335_NO_SHIFT_REG;
assign rnode_333to335_bb3_shr16_i510_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_333to335_bb3_shr16_i510_1_NO_SHIFT_REG = rnode_333to335_bb3_shr16_i510_0_reg_335_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_333to334_bb3_lnot23_i517_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to334_bb3_lnot23_i517_0_stall_in_NO_SHIFT_REG;
 logic rnode_333to334_bb3_lnot23_i517_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3_lnot23_i517_0_reg_334_inputs_ready_NO_SHIFT_REG;
 logic rnode_333to334_bb3_lnot23_i517_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_lnot23_i517_0_valid_out_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_lnot23_i517_0_stall_in_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_lnot23_i517_0_stall_out_reg_334_NO_SHIFT_REG;

acl_data_fifo rnode_333to334_bb3_lnot23_i517_0_reg_334_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to334_bb3_lnot23_i517_0_reg_334_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to334_bb3_lnot23_i517_0_stall_in_reg_334_NO_SHIFT_REG),
	.valid_out(rnode_333to334_bb3_lnot23_i517_0_valid_out_reg_334_NO_SHIFT_REG),
	.stall_out(rnode_333to334_bb3_lnot23_i517_0_stall_out_reg_334_NO_SHIFT_REG),
	.data_in(local_bb3_lnot23_i517),
	.data_out(rnode_333to334_bb3_lnot23_i517_0_reg_334_NO_SHIFT_REG)
);

defparam rnode_333to334_bb3_lnot23_i517_0_reg_334_fifo.DEPTH = 1;
defparam rnode_333to334_bb3_lnot23_i517_0_reg_334_fifo.DATA_WIDTH = 1;
defparam rnode_333to334_bb3_lnot23_i517_0_reg_334_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to334_bb3_lnot23_i517_0_reg_334_fifo.IMPL = "shift_reg";

assign rnode_333to334_bb3_lnot23_i517_0_reg_334_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_lnot23_i517_stall_in = 1'b0;
assign rnode_333to334_bb3_lnot23_i517_0_NO_SHIFT_REG = rnode_333to334_bb3_lnot23_i517_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3_lnot23_i517_0_stall_in_reg_334_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_lnot23_i517_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_333to335_bb3_cmp27_i519_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_1_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_2_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_valid_out_0_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_stall_in_0_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_cmp27_i519_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_333to335_bb3_cmp27_i519_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to335_bb3_cmp27_i519_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to335_bb3_cmp27_i519_0_stall_in_0_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_333to335_bb3_cmp27_i519_0_valid_out_0_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_333to335_bb3_cmp27_i519_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in(local_bb3_cmp27_i519),
	.data_out(rnode_333to335_bb3_cmp27_i519_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_333to335_bb3_cmp27_i519_0_reg_335_fifo.DEPTH = 2;
defparam rnode_333to335_bb3_cmp27_i519_0_reg_335_fifo.DATA_WIDTH = 1;
defparam rnode_333to335_bb3_cmp27_i519_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to335_bb3_cmp27_i519_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_333to335_bb3_cmp27_i519_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp27_i519_stall_in = 1'b0;
assign rnode_333to335_bb3_cmp27_i519_0_stall_in_0_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_333to335_bb3_cmp27_i519_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_333to335_bb3_cmp27_i519_0_NO_SHIFT_REG = rnode_333to335_bb3_cmp27_i519_0_reg_335_NO_SHIFT_REG;
assign rnode_333to335_bb3_cmp27_i519_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_333to335_bb3_cmp27_i519_1_NO_SHIFT_REG = rnode_333to335_bb3_cmp27_i519_0_reg_335_NO_SHIFT_REG;
assign rnode_333to335_bb3_cmp27_i519_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_333to335_bb3_cmp27_i519_2_NO_SHIFT_REG = rnode_333to335_bb3_cmp27_i519_0_reg_335_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_333to334_bb3_align_0_i539_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_align_0_i539_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_align_0_i539_1_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_align_0_i539_2_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_align_0_i539_3_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_align_0_i539_4_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_reg_334_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_align_0_i539_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_valid_out_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_stall_in_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_align_0_i539_0_stall_out_reg_334_NO_SHIFT_REG;

acl_data_fifo rnode_333to334_bb3_align_0_i539_0_reg_334_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to334_bb3_align_0_i539_0_reg_334_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to334_bb3_align_0_i539_0_stall_in_0_reg_334_NO_SHIFT_REG),
	.valid_out(rnode_333to334_bb3_align_0_i539_0_valid_out_0_reg_334_NO_SHIFT_REG),
	.stall_out(rnode_333to334_bb3_align_0_i539_0_stall_out_reg_334_NO_SHIFT_REG),
	.data_in((local_bb3_align_0_i539 & 32'hFF)),
	.data_out(rnode_333to334_bb3_align_0_i539_0_reg_334_NO_SHIFT_REG)
);

defparam rnode_333to334_bb3_align_0_i539_0_reg_334_fifo.DEPTH = 1;
defparam rnode_333to334_bb3_align_0_i539_0_reg_334_fifo.DATA_WIDTH = 32;
defparam rnode_333to334_bb3_align_0_i539_0_reg_334_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to334_bb3_align_0_i539_0_reg_334_fifo.IMPL = "shift_reg";

assign rnode_333to334_bb3_align_0_i539_0_reg_334_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_align_0_i539_stall_in = 1'b0;
assign rnode_333to334_bb3_align_0_i539_0_stall_in_0_reg_334_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_align_0_i539_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3_align_0_i539_0_NO_SHIFT_REG = rnode_333to334_bb3_align_0_i539_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3_align_0_i539_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3_align_0_i539_1_NO_SHIFT_REG = rnode_333to334_bb3_align_0_i539_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3_align_0_i539_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3_align_0_i539_2_NO_SHIFT_REG = rnode_333to334_bb3_align_0_i539_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3_align_0_i539_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3_align_0_i539_3_NO_SHIFT_REG = rnode_333to334_bb3_align_0_i539_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3_align_0_i539_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3_align_0_i539_4_NO_SHIFT_REG = rnode_333to334_bb3_align_0_i539_0_reg_334_NO_SHIFT_REG;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_333to336_bb3_xor_i316_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to336_bb3_xor_i316_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_333to336_bb3_xor_i316_0_NO_SHIFT_REG;
 logic rnode_333to336_bb3_xor_i316_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to336_bb3_xor_i316_0_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3_xor_i316_0_valid_out_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3_xor_i316_0_stall_in_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3_xor_i316_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_333to336_bb3_xor_i316_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to336_bb3_xor_i316_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to336_bb3_xor_i316_0_stall_in_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_333to336_bb3_xor_i316_0_valid_out_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_333to336_bb3_xor_i316_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3_xor_i316_0_NO_SHIFT_REG),
	.data_out(rnode_333to336_bb3_xor_i316_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_333to336_bb3_xor_i316_0_reg_336_fifo.DEPTH = 3;
defparam rnode_333to336_bb3_xor_i316_0_reg_336_fifo.DATA_WIDTH = 32;
defparam rnode_333to336_bb3_xor_i316_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to336_bb3_xor_i316_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_333to336_bb3_xor_i316_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_xor_i316_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to336_bb3_xor_i316_0_NO_SHIFT_REG = rnode_333to336_bb3_xor_i316_0_reg_336_NO_SHIFT_REG;
assign rnode_333to336_bb3_xor_i316_0_stall_in_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_333to336_bb3_xor_i316_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_333to334_bb3_add_i357_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to334_bb3_add_i357_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_add_i357_0_NO_SHIFT_REG;
 logic rnode_333to334_bb3_add_i357_0_reg_334_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_333to334_bb3_add_i357_0_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_add_i357_0_valid_out_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_add_i357_0_stall_in_reg_334_NO_SHIFT_REG;
 logic rnode_333to334_bb3_add_i357_0_stall_out_reg_334_NO_SHIFT_REG;

acl_data_fifo rnode_333to334_bb3_add_i357_0_reg_334_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to334_bb3_add_i357_0_reg_334_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to334_bb3_add_i357_0_stall_in_reg_334_NO_SHIFT_REG),
	.valid_out(rnode_333to334_bb3_add_i357_0_valid_out_reg_334_NO_SHIFT_REG),
	.stall_out(rnode_333to334_bb3_add_i357_0_stall_out_reg_334_NO_SHIFT_REG),
	.data_in((rnode_332to333_bb3_add_i357_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_333to334_bb3_add_i357_0_reg_334_NO_SHIFT_REG)
);

defparam rnode_333to334_bb3_add_i357_0_reg_334_fifo.DEPTH = 1;
defparam rnode_333to334_bb3_add_i357_0_reg_334_fifo.DATA_WIDTH = 32;
defparam rnode_333to334_bb3_add_i357_0_reg_334_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to334_bb3_add_i357_0_reg_334_fifo.IMPL = "shift_reg";

assign rnode_333to334_bb3_add_i357_0_reg_334_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_add_i357_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_add_i357_0_NO_SHIFT_REG = rnode_333to334_bb3_add_i357_0_reg_334_NO_SHIFT_REG;
assign rnode_333to334_bb3_add_i357_0_stall_in_reg_334_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_add_i357_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_conv3_i_i351_stall_local;
wire [31:0] local_bb3_conv3_i_i351;
wire [63:0] local_bb3_conv3_i_i351$ps;

assign local_bb3_conv3_i_i351$ps = (local_bb3_mul_i_i350 & 64'hFFFFFFFFFFFF);
assign local_bb3_conv3_i_i351 = local_bb3_conv3_i_i351$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_var__u26_stall_local;
wire [63:0] local_bb3_var__u26;

assign local_bb3_var__u26 = ((local_bb3_mul_i_i350 & 64'hFFFFFFFFFFFF) >> 64'h18);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_333to336_bb3_reduction_0_i375_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to336_bb3_reduction_0_i375_0_stall_in_NO_SHIFT_REG;
 logic rnode_333to336_bb3_reduction_0_i375_0_NO_SHIFT_REG;
 logic rnode_333to336_bb3_reduction_0_i375_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic rnode_333to336_bb3_reduction_0_i375_0_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3_reduction_0_i375_0_valid_out_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3_reduction_0_i375_0_stall_in_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3_reduction_0_i375_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_333to336_bb3_reduction_0_i375_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to336_bb3_reduction_0_i375_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to336_bb3_reduction_0_i375_0_stall_in_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_333to336_bb3_reduction_0_i375_0_valid_out_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_333to336_bb3_reduction_0_i375_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3_reduction_0_i375_0_NO_SHIFT_REG),
	.data_out(rnode_333to336_bb3_reduction_0_i375_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_333to336_bb3_reduction_0_i375_0_reg_336_fifo.DEPTH = 3;
defparam rnode_333to336_bb3_reduction_0_i375_0_reg_336_fifo.DATA_WIDTH = 1;
defparam rnode_333to336_bb3_reduction_0_i375_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to336_bb3_reduction_0_i375_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_333to336_bb3_reduction_0_i375_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_reduction_0_i375_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to336_bb3_reduction_0_i375_0_NO_SHIFT_REG = rnode_333to336_bb3_reduction_0_i375_0_reg_336_NO_SHIFT_REG;
assign rnode_333to336_bb3_reduction_0_i375_0_stall_in_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_333to336_bb3_reduction_0_i375_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_333to335_bb3_var__u23_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to335_bb3_var__u23_0_stall_in_NO_SHIFT_REG;
 logic rnode_333to335_bb3_var__u23_0_NO_SHIFT_REG;
 logic rnode_333to335_bb3_var__u23_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic rnode_333to335_bb3_var__u23_0_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_var__u23_0_valid_out_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_var__u23_0_stall_in_reg_335_NO_SHIFT_REG;
 logic rnode_333to335_bb3_var__u23_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_333to335_bb3_var__u23_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to335_bb3_var__u23_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to335_bb3_var__u23_0_stall_in_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_333to335_bb3_var__u23_0_valid_out_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_333to335_bb3_var__u23_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3_var__u23_0_NO_SHIFT_REG),
	.data_out(rnode_333to335_bb3_var__u23_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_333to335_bb3_var__u23_0_reg_335_fifo.DEPTH = 2;
defparam rnode_333to335_bb3_var__u23_0_reg_335_fifo.DATA_WIDTH = 1;
defparam rnode_333to335_bb3_var__u23_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to335_bb3_var__u23_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_333to335_bb3_var__u23_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3_var__u23_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to335_bb3_var__u23_0_NO_SHIFT_REG = rnode_333to335_bb3_var__u23_0_reg_335_NO_SHIFT_REG;
assign rnode_333to335_bb3_var__u23_0_stall_in_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_333to335_bb3_var__u23_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_333to336_bb3__29_i345_0_valid_out_NO_SHIFT_REG;
 logic rnode_333to336_bb3__29_i345_0_stall_in_NO_SHIFT_REG;
 logic rnode_333to336_bb3__29_i345_0_NO_SHIFT_REG;
 logic rnode_333to336_bb3__29_i345_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic rnode_333to336_bb3__29_i345_0_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3__29_i345_0_valid_out_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3__29_i345_0_stall_in_reg_336_NO_SHIFT_REG;
 logic rnode_333to336_bb3__29_i345_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_333to336_bb3__29_i345_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_333to336_bb3__29_i345_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_333to336_bb3__29_i345_0_stall_in_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_333to336_bb3__29_i345_0_valid_out_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_333to336_bb3__29_i345_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in(rnode_332to333_bb3__29_i345_0_NO_SHIFT_REG),
	.data_out(rnode_333to336_bb3__29_i345_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_333to336_bb3__29_i345_0_reg_336_fifo.DEPTH = 3;
defparam rnode_333to336_bb3__29_i345_0_reg_336_fifo.DATA_WIDTH = 1;
defparam rnode_333to336_bb3__29_i345_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_333to336_bb3__29_i345_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_333to336_bb3__29_i345_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_332to333_bb3__29_i345_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to336_bb3__29_i345_0_NO_SHIFT_REG = rnode_333to336_bb3__29_i345_0_reg_336_NO_SHIFT_REG;
assign rnode_333to336_bb3__29_i345_0_stall_in_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_333to336_bb3__29_i345_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_346_347_0_inputs_ready;
 reg SFC_1_VALID_346_347_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_346_347_0_stall_in;
wire SFC_1_VALID_346_347_0_output_regs_ready;
 reg SFC_1_VALID_346_347_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_346_347_0_causedstall;

assign SFC_1_VALID_346_347_0_inputs_ready = 1'b1;
assign SFC_1_VALID_346_347_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_345_346_0_stall_in = 1'b0;
assign SFC_1_VALID_346_347_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_346_347_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_346_347_0_output_regs_ready)
		begin
			SFC_1_VALID_346_347_0_NO_SHIFT_REG <= SFC_1_VALID_345_346_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and21_i515_stall_local;
wire [31:0] local_bb3_and21_i515;

assign local_bb3_and21_i515 = (rnode_333to334_bb3__22_i508_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and20_i514_valid_out;
wire local_bb3_and20_i514_stall_in;
wire local_bb3_and20_i514_inputs_ready;
wire local_bb3_and20_i514_stall_local;
wire [31:0] local_bb3_and20_i514;

assign local_bb3_and20_i514_inputs_ready = rnode_333to334_bb3__23_i509_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_and20_i514 = (rnode_333to334_bb3__23_i509_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb3_and20_i514_valid_out = 1'b1;
assign rnode_333to334_bb3__23_i509_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and35_i520_valid_out;
wire local_bb3_and35_i520_stall_in;
wire local_bb3_and35_i520_inputs_ready;
wire local_bb3_and35_i520_stall_local;
wire [31:0] local_bb3_and35_i520;

assign local_bb3_and35_i520_inputs_ready = rnode_333to334_bb3__23_i509_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_and35_i520 = (rnode_333to334_bb3__23_i509_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb3_and35_i520_valid_out = 1'b1;
assign rnode_333to334_bb3__23_i509_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_xor36_i_stall_local;
wire [31:0] local_bb3_xor36_i;

assign local_bb3_xor36_i = (rnode_333to334_bb3__23_i509_2_NO_SHIFT_REG ^ rnode_333to334_bb3__22_i508_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_and17_i511_stall_local;
wire [31:0] local_bb3_and17_i511;

assign local_bb3_and17_i511 = ((rnode_333to335_bb3_shr16_i510_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_335to337_bb3_shr16_i510_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to337_bb3_shr16_i510_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_shr16_i510_0_NO_SHIFT_REG;
 logic rnode_335to337_bb3_shr16_i510_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_shr16_i510_0_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_shr16_i510_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_shr16_i510_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_shr16_i510_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_335to337_bb3_shr16_i510_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to337_bb3_shr16_i510_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to337_bb3_shr16_i510_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_335to337_bb3_shr16_i510_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_335to337_bb3_shr16_i510_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((rnode_333to335_bb3_shr16_i510_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_335to337_bb3_shr16_i510_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_335to337_bb3_shr16_i510_0_reg_337_fifo.DEPTH = 2;
defparam rnode_335to337_bb3_shr16_i510_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_335to337_bb3_shr16_i510_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to337_bb3_shr16_i510_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_335to337_bb3_shr16_i510_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to335_bb3_shr16_i510_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_shr16_i510_0_NO_SHIFT_REG = rnode_335to337_bb3_shr16_i510_0_reg_337_NO_SHIFT_REG;
assign rnode_335to337_bb3_shr16_i510_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_shr16_i510_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and94_i_stall_local;
wire [31:0] local_bb3_and94_i;

assign local_bb3_and94_i = ((rnode_333to334_bb3_align_0_i539_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb3_and96_i_stall_local;
wire [31:0] local_bb3_and96_i;

assign local_bb3_and96_i = ((rnode_333to334_bb3_align_0_i539_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and116_i_stall_local;
wire [31:0] local_bb3_and116_i;

assign local_bb3_and116_i = ((rnode_333to334_bb3_align_0_i539_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_and131_i_stall_local;
wire [31:0] local_bb3_and131_i;

assign local_bb3_and131_i = ((rnode_333to334_bb3_align_0_i539_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb3_and150_i_stall_local;
wire [31:0] local_bb3_and150_i;

assign local_bb3_and150_i = ((rnode_333to334_bb3_align_0_i539_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_xor_i316_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_xor_i316_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_xor_i316_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_xor_i316_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_xor_i316_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_xor_i316_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_xor_i316_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_xor_i316_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_xor_i316_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_xor_i316_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_xor_i316_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_xor_i316_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_xor_i316_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(rnode_333to336_bb3_xor_i316_0_NO_SHIFT_REG),
	.data_out(rnode_336to337_bb3_xor_i316_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_xor_i316_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_xor_i316_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_336to337_bb3_xor_i316_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_xor_i316_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_xor_i316_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to336_bb3_xor_i316_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_xor_i316_0_NO_SHIFT_REG = rnode_336to337_bb3_xor_i316_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_xor_i316_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_xor_i316_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_334to335_bb3_add_i357_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_add_i357_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_add_i357_1_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_add_i357_2_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_add_i357_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_valid_out_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_stall_in_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_add_i357_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_334to335_bb3_add_i357_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_334to335_bb3_add_i357_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_334to335_bb3_add_i357_0_stall_in_0_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_334to335_bb3_add_i357_0_valid_out_0_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_334to335_bb3_add_i357_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in((rnode_333to334_bb3_add_i357_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_334to335_bb3_add_i357_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_334to335_bb3_add_i357_0_reg_335_fifo.DEPTH = 1;
defparam rnode_334to335_bb3_add_i357_0_reg_335_fifo.DATA_WIDTH = 32;
defparam rnode_334to335_bb3_add_i357_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_334to335_bb3_add_i357_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_334to335_bb3_add_i357_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to334_bb3_add_i357_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_add_i357_0_stall_in_0_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_add_i357_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_add_i357_0_NO_SHIFT_REG = rnode_334to335_bb3_add_i357_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_add_i357_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_add_i357_1_NO_SHIFT_REG = rnode_334to335_bb3_add_i357_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_add_i357_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_add_i357_2_NO_SHIFT_REG = rnode_334to335_bb3_add_i357_0_reg_335_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i16_i354_stall_local;
wire [31:0] local_bb3_shr_i16_i354;

assign local_bb3_shr_i16_i354 = (local_bb3_conv3_i_i351 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i18_i356_stall_local;
wire [31:0] local_bb3_shl1_i18_i356;

assign local_bb3_shl1_i18_i356 = (local_bb3_conv3_i_i351 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u27_stall_local;
wire [31:0] local_bb3_var__u27;

assign local_bb3_var__u27 = (local_bb3_conv3_i_i351 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i_i364_stall_local;
wire [31:0] local_bb3_shl1_i_i364;

assign local_bb3_shl1_i_i364 = (local_bb3_conv3_i_i351 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb3__tr_i352_stall_local;
wire [31:0] local_bb3__tr_i352;
wire [63:0] local_bb3__tr_i352$ps;

assign local_bb3__tr_i352$ps = (local_bb3_var__u26 & 64'hFFFFFF);
assign local_bb3__tr_i352 = local_bb3__tr_i352$ps[31:0];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_reduction_0_i375_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_reduction_0_i375_0_stall_in_NO_SHIFT_REG;
 logic rnode_336to337_bb3_reduction_0_i375_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_reduction_0_i375_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to337_bb3_reduction_0_i375_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_reduction_0_i375_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_reduction_0_i375_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_reduction_0_i375_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_reduction_0_i375_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_reduction_0_i375_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_reduction_0_i375_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_reduction_0_i375_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_reduction_0_i375_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(rnode_333to336_bb3_reduction_0_i375_0_NO_SHIFT_REG),
	.data_out(rnode_336to337_bb3_reduction_0_i375_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_reduction_0_i375_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_reduction_0_i375_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_336to337_bb3_reduction_0_i375_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_reduction_0_i375_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_reduction_0_i375_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to336_bb3_reduction_0_i375_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_reduction_0_i375_0_NO_SHIFT_REG = rnode_336to337_bb3_reduction_0_i375_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_reduction_0_i375_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_reduction_0_i375_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_335to336_bb3_var__u23_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u23_0_stall_in_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u23_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u23_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u23_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u23_0_valid_out_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u23_0_stall_in_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u23_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_335to336_bb3_var__u23_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to336_bb3_var__u23_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to336_bb3_var__u23_0_stall_in_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_335to336_bb3_var__u23_0_valid_out_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_335to336_bb3_var__u23_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in(rnode_333to335_bb3_var__u23_0_NO_SHIFT_REG),
	.data_out(rnode_335to336_bb3_var__u23_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_335to336_bb3_var__u23_0_reg_336_fifo.DEPTH = 1;
defparam rnode_335to336_bb3_var__u23_0_reg_336_fifo.DATA_WIDTH = 1;
defparam rnode_335to336_bb3_var__u23_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to336_bb3_var__u23_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_335to336_bb3_var__u23_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to335_bb3_var__u23_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3_var__u23_0_NO_SHIFT_REG = rnode_335to336_bb3_var__u23_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3_var__u23_0_stall_in_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3_var__u23_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3__29_i345_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3__29_i345_0_stall_in_NO_SHIFT_REG;
 logic rnode_336to337_bb3__29_i345_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3__29_i345_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to337_bb3__29_i345_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__29_i345_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__29_i345_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__29_i345_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3__29_i345_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3__29_i345_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3__29_i345_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3__29_i345_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3__29_i345_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(rnode_333to336_bb3__29_i345_0_NO_SHIFT_REG),
	.data_out(rnode_336to337_bb3__29_i345_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3__29_i345_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3__29_i345_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_336to337_bb3__29_i345_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3__29_i345_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3__29_i345_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_333to336_bb3__29_i345_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__29_i345_0_NO_SHIFT_REG = rnode_336to337_bb3__29_i345_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3__29_i345_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__29_i345_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_347_348_0_inputs_ready;
 reg SFC_1_VALID_347_348_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_347_348_0_stall_in;
wire SFC_1_VALID_347_348_0_output_regs_ready;
 reg SFC_1_VALID_347_348_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_347_348_0_causedstall;

assign SFC_1_VALID_347_348_0_inputs_ready = 1'b1;
assign SFC_1_VALID_347_348_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_346_347_0_stall_in = 1'b0;
assign SFC_1_VALID_347_348_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_347_348_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_347_348_0_output_regs_ready)
		begin
			SFC_1_VALID_347_348_0_NO_SHIFT_REG <= SFC_1_VALID_346_347_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_lnot33_not_i524_stall_local;
wire local_bb3_lnot33_not_i524;

assign local_bb3_lnot33_not_i524 = ((local_bb3_and21_i515 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or65_i_stall_local;
wire [31:0] local_bb3_or65_i;

assign local_bb3_or65_i = ((local_bb3_and21_i515 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_334to335_bb3_and20_i514_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and20_i514_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_and20_i514_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and20_i514_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and20_i514_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_and20_i514_1_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and20_i514_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_and20_i514_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and20_i514_0_valid_out_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and20_i514_0_stall_in_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and20_i514_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_334to335_bb3_and20_i514_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_334to335_bb3_and20_i514_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_334to335_bb3_and20_i514_0_stall_in_0_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_334to335_bb3_and20_i514_0_valid_out_0_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_334to335_bb3_and20_i514_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in((local_bb3_and20_i514 & 32'h7FFFFF)),
	.data_out(rnode_334to335_bb3_and20_i514_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_334to335_bb3_and20_i514_0_reg_335_fifo.DEPTH = 1;
defparam rnode_334to335_bb3_and20_i514_0_reg_335_fifo.DATA_WIDTH = 32;
defparam rnode_334to335_bb3_and20_i514_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_334to335_bb3_and20_i514_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_334to335_bb3_and20_i514_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and20_i514_stall_in = 1'b0;
assign rnode_334to335_bb3_and20_i514_0_stall_in_0_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_and20_i514_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_and20_i514_0_NO_SHIFT_REG = rnode_334to335_bb3_and20_i514_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_and20_i514_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_and20_i514_1_NO_SHIFT_REG = rnode_334to335_bb3_and20_i514_0_reg_335_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_334to335_bb3_and35_i520_0_valid_out_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and35_i520_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_and35_i520_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and35_i520_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_and35_i520_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and35_i520_0_valid_out_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and35_i520_0_stall_in_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and35_i520_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_334to335_bb3_and35_i520_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_334to335_bb3_and35_i520_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_334to335_bb3_and35_i520_0_stall_in_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_334to335_bb3_and35_i520_0_valid_out_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_334to335_bb3_and35_i520_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in((local_bb3_and35_i520 & 32'h80000000)),
	.data_out(rnode_334to335_bb3_and35_i520_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_334to335_bb3_and35_i520_0_reg_335_fifo.DEPTH = 1;
defparam rnode_334to335_bb3_and35_i520_0_reg_335_fifo.DATA_WIDTH = 32;
defparam rnode_334to335_bb3_and35_i520_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_334to335_bb3_and35_i520_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_334to335_bb3_and35_i520_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and35_i520_stall_in = 1'b0;
assign rnode_334to335_bb3_and35_i520_0_NO_SHIFT_REG = rnode_334to335_bb3_and35_i520_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_and35_i520_0_stall_in_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_and35_i520_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp38_i_stall_local;
wire local_bb3_cmp38_i;

assign local_bb3_cmp38_i = ($signed(local_bb3_xor36_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb3_xor36_lobit_i_stall_local;
wire [31:0] local_bb3_xor36_lobit_i;

assign local_bb3_xor36_lobit_i = ($signed(local_bb3_xor36_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_and37_lobit_i_stall_local;
wire [31:0] local_bb3_and37_lobit_i;

assign local_bb3_and37_lobit_i = (local_bb3_xor36_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_i516_stall_local;
wire local_bb3_lnot_i516;

assign local_bb3_lnot_i516 = ((local_bb3_and17_i511 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_i518_stall_local;
wire local_bb3_cmp25_i518;

assign local_bb3_cmp25_i518 = ((local_bb3_and17_i511 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp97_i_stall_local;
wire local_bb3_cmp97_i;

assign local_bb3_cmp97_i = ((local_bb3_and96_i & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp117_i_stall_local;
wire local_bb3_cmp117_i;

assign local_bb3_cmp117_i = ((local_bb3_and116_i & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp132_not_i_stall_local;
wire local_bb3_cmp132_not_i;

assign local_bb3_cmp132_not_i = ((local_bb3_and131_i & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_Pivot20_i550_stall_local;
wire local_bb3_Pivot20_i550;

assign local_bb3_Pivot20_i550 = ((local_bb3_and150_i & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_SwitchLeaf_i551_stall_local;
wire local_bb3_SwitchLeaf_i551;

assign local_bb3_SwitchLeaf_i551 = ((local_bb3_and150_i & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and4_i317_stall_local;
wire [31:0] local_bb3_and4_i317;

assign local_bb3_and4_i317 = (rnode_336to337_bb3_xor_i316_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_inc_i360_stall_local;
wire [31:0] local_bb3_inc_i360;

assign local_bb3_inc_i360 = ((rnode_334to335_bb3_add_i357_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp50_not_i365_stall_local;
wire local_bb3_cmp50_not_i365;

assign local_bb3_cmp50_not_i365 = ((rnode_334to335_bb3_add_i357_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i_i362_stall_local;
wire [31:0] local_bb3_shr_i_i362;

assign local_bb3_shr_i_i362 = ((local_bb3_var__u27 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i15_i353_stall_local;
wire [31:0] local_bb3_shl_i15_i353;

assign local_bb3_shl_i15_i353 = ((local_bb3__tr_i352 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb3_and48_i358_stall_local;
wire [31:0] local_bb3_and48_i358;

assign local_bb3_and48_i358 = ((local_bb3__tr_i352 & 32'hFFFFFF) & 32'h800000);

// This section implements a registered operation.
// 
wire SFC_1_VALID_348_349_0_inputs_ready;
 reg SFC_1_VALID_348_349_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_348_349_0_stall_in;
wire SFC_1_VALID_348_349_0_output_regs_ready;
 reg SFC_1_VALID_348_349_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_348_349_0_causedstall;

assign SFC_1_VALID_348_349_0_inputs_ready = 1'b1;
assign SFC_1_VALID_348_349_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_347_348_0_stall_in = 1'b0;
assign SFC_1_VALID_348_349_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_348_349_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_348_349_0_output_regs_ready)
		begin
			SFC_1_VALID_348_349_0_NO_SHIFT_REG <= SFC_1_VALID_347_348_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_shl66_i_stall_local;
wire [31:0] local_bb3_shl66_i;

assign local_bb3_shl66_i = ((local_bb3_or65_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot30_i522_stall_local;
wire local_bb3_lnot30_i522;

assign local_bb3_lnot30_i522 = ((rnode_334to335_bb3_and20_i514_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i534_stall_local;
wire [31:0] local_bb3_or_i534;

assign local_bb3_or_i534 = ((rnode_334to335_bb3_and20_i514_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_335to337_bb3_and35_i520_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and35_i520_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_and35_i520_0_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and35_i520_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_and35_i520_0_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and35_i520_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and35_i520_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and35_i520_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_335to337_bb3_and35_i520_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to337_bb3_and35_i520_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to337_bb3_and35_i520_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_335to337_bb3_and35_i520_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_335to337_bb3_and35_i520_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((rnode_334to335_bb3_and35_i520_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_335to337_bb3_and35_i520_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_335to337_bb3_and35_i520_0_reg_337_fifo.DEPTH = 2;
defparam rnode_335to337_bb3_and35_i520_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_335to337_bb3_and35_i520_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to337_bb3_and35_i520_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_335to337_bb3_and35_i520_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_and35_i520_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_and35_i520_0_NO_SHIFT_REG = rnode_335to337_bb3_and35_i520_0_reg_337_NO_SHIFT_REG;
assign rnode_335to337_bb3_and35_i520_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_and35_i520_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_not_i521_stall_local;
wire local_bb3_cmp25_not_i521;

assign local_bb3_cmp25_not_i521 = (local_bb3_cmp25_i518 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u28_stall_local;
wire local_bb3_var__u28;

assign local_bb3_var__u28 = (local_bb3_cmp25_i518 | rnode_333to335_bb3_cmp27_i519_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i17_i355_stall_local;
wire [31:0] local_bb3_or_i17_i355;

assign local_bb3_or_i17_i355 = ((local_bb3_shl_i15_i353 & 32'hFFFF00) | (local_bb3_shr_i16_i354 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool49_i359_stall_local;
wire local_bb3_tobool49_i359;

assign local_bb3_tobool49_i359 = ((local_bb3_and48_i358 & 32'h800000) == 32'h0);

// This section implements a registered operation.
// 
wire SFC_1_VALID_349_350_0_inputs_ready;
 reg SFC_1_VALID_349_350_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_349_350_0_stall_in;
wire SFC_1_VALID_349_350_0_output_regs_ready;
 reg SFC_1_VALID_349_350_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_349_350_0_causedstall;

assign SFC_1_VALID_349_350_0_inputs_ready = 1'b1;
assign SFC_1_VALID_349_350_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_348_349_0_stall_in = 1'b0;
assign SFC_1_VALID_349_350_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_349_350_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_349_350_0_output_regs_ready)
		begin
			SFC_1_VALID_349_350_0_NO_SHIFT_REG <= SFC_1_VALID_348_349_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__28_i537_stall_local;
wire [31:0] local_bb3__28_i537;

assign local_bb3__28_i537 = (rnode_333to334_bb3_lnot23_i517_0_NO_SHIFT_REG ? 32'h0 : ((local_bb3_shl66_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot30_not_i526_stall_local;
wire local_bb3_lnot30_not_i526;

assign local_bb3_lnot30_not_i526 = (local_bb3_lnot30_i522 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i535_stall_local;
wire [31:0] local_bb3_shl_i535;

assign local_bb3_shl_i535 = ((local_bb3_or_i534 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_337to338_bb3_and35_i520_0_valid_out_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and35_i520_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_and35_i520_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and35_i520_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_and35_i520_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and35_i520_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and35_i520_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and35_i520_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_337to338_bb3_and35_i520_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to338_bb3_and35_i520_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to338_bb3_and35_i520_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_337to338_bb3_and35_i520_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_337to338_bb3_and35_i520_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in((rnode_335to337_bb3_and35_i520_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_337to338_bb3_and35_i520_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_337to338_bb3_and35_i520_0_reg_338_fifo.DEPTH = 1;
defparam rnode_337to338_bb3_and35_i520_0_reg_338_fifo.DATA_WIDTH = 32;
defparam rnode_337to338_bb3_and35_i520_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to338_bb3_and35_i520_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_337to338_bb3_and35_i520_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_335to337_bb3_and35_i520_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_and35_i520_0_NO_SHIFT_REG = rnode_337to338_bb3_and35_i520_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3_and35_i520_0_stall_in_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_and35_i520_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_or_cond_i523_stall_local;
wire local_bb3_or_cond_i523;

assign local_bb3_or_cond_i523 = (local_bb3_lnot30_i522 | local_bb3_cmp25_not_i521);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i_i361_stall_local;
wire [31:0] local_bb3_shl_i_i361;

assign local_bb3_shl_i_i361 = ((local_bb3_or_i17_i355 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__31_i366_stall_local;
wire local_bb3__31_i366;

assign local_bb3__31_i366 = (local_bb3_tobool49_i359 & local_bb3_cmp50_not_i365);

// This section implements a registered operation.
// 
wire SFC_1_VALID_350_351_0_inputs_ready;
 reg SFC_1_VALID_350_351_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_350_351_0_stall_in;
wire SFC_1_VALID_350_351_0_output_regs_ready;
 reg SFC_1_VALID_350_351_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_350_351_0_causedstall;

assign SFC_1_VALID_350_351_0_inputs_ready = 1'b1;
assign SFC_1_VALID_350_351_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_349_350_0_stall_in = 1'b0;
assign SFC_1_VALID_350_351_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_350_351_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_350_351_0_output_regs_ready)
		begin
			SFC_1_VALID_350_351_0_NO_SHIFT_REG <= SFC_1_VALID_349_350_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and73_i_stall_local;
wire [31:0] local_bb3_and73_i;

assign local_bb3_and73_i = ((local_bb3__28_i537 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb3_and76_i_stall_local;
wire [31:0] local_bb3_and76_i;

assign local_bb3_and76_i = ((local_bb3__28_i537 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb3_and79_i_stall_local;
wire [31:0] local_bb3_and79_i;

assign local_bb3_and79_i = ((local_bb3__28_i537 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb3_shr95_i_stall_local;
wire [31:0] local_bb3_shr95_i;

assign local_bb3_shr95_i = ((local_bb3__28_i537 & 32'h7FFFFF8) >> (local_bb3_and94_i & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb3_and91_i_stall_local;
wire [31:0] local_bb3_and91_i;

assign local_bb3_and91_i = ((local_bb3__28_i537 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb3_and88_i541_stall_local;
wire [31:0] local_bb3_and88_i541;

assign local_bb3_and88_i541 = ((local_bb3__28_i537 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb3_and85_i_stall_local;
wire [31:0] local_bb3_and85_i;

assign local_bb3_and85_i = ((local_bb3__28_i537 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u29_stall_local;
wire [31:0] local_bb3_var__u29;

assign local_bb3_var__u29 = ((local_bb3__28_i537 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb3_or_cond_not_i527_stall_local;
wire local_bb3_or_cond_not_i527;

assign local_bb3_or_cond_not_i527 = (local_bb3_cmp25_i518 & local_bb3_lnot30_not_i526);

// This section implements an unregistered operation.
// 
wire local_bb3__27_i536_stall_local;
wire [31:0] local_bb3__27_i536;

assign local_bb3__27_i536 = (local_bb3_lnot_i516 ? 32'h0 : ((local_bb3_shl_i535 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_8_i531_stall_local;
wire local_bb3_reduction_8_i531;

assign local_bb3_reduction_8_i531 = (rnode_333to335_bb3_cmp27_i519_1_NO_SHIFT_REG & local_bb3_or_cond_i523);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i_i363_stall_local;
wire [31:0] local_bb3_or_i_i363;

assign local_bb3_or_i_i363 = ((local_bb3_shl_i_i361 & 32'h1FFFFFE) | (local_bb3_shr_i_i362 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__32_i367_stall_local;
wire [31:0] local_bb3__32_i367;

assign local_bb3__32_i367 = (local_bb3__31_i366 ? (local_bb3_shl1_i_i364 & 32'hFFFFFE00) : (local_bb3_shl1_i18_i356 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__36_i371_stall_local;
wire [31:0] local_bb3__36_i371;

assign local_bb3__36_i371 = (local_bb3__31_i366 ? (rnode_334to335_bb3_add_i357_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements a registered operation.
// 
wire SFC_1_VALID_351_352_0_inputs_ready;
 reg SFC_1_VALID_351_352_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_351_352_0_stall_in;
wire SFC_1_VALID_351_352_0_output_regs_ready;
 reg SFC_1_VALID_351_352_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_351_352_0_causedstall;

assign SFC_1_VALID_351_352_0_inputs_ready = 1'b1;
assign SFC_1_VALID_351_352_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_350_351_0_stall_in = 1'b0;
assign SFC_1_VALID_351_352_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_351_352_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_351_352_0_output_regs_ready)
		begin
			SFC_1_VALID_351_352_0_NO_SHIFT_REG <= SFC_1_VALID_350_351_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and73_tr_i_stall_local;
wire [7:0] local_bb3_and73_tr_i;
wire [31:0] local_bb3_and73_tr_i$ps;

assign local_bb3_and73_tr_i$ps = (local_bb3_and73_i & 32'hFFFFFF);
assign local_bb3_and73_tr_i = local_bb3_and73_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb3_cmp77_i540_stall_local;
wire local_bb3_cmp77_i540;

assign local_bb3_cmp77_i540 = ((local_bb3_and76_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp80_i_stall_local;
wire local_bb3_cmp80_i;

assign local_bb3_cmp80_i = ((local_bb3_and79_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and143_i_stall_local;
wire [31:0] local_bb3_and143_i;

assign local_bb3_and143_i = (local_bb3_shr95_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_shr151_i_stall_local;
wire [31:0] local_bb3_shr151_i;

assign local_bb3_shr151_i = (local_bb3_shr95_i >> (local_bb3_and150_i & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u30_stall_local;
wire [31:0] local_bb3_var__u30;

assign local_bb3_var__u30 = (local_bb3_shr95_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and147_i_stall_local;
wire [31:0] local_bb3_and147_i;

assign local_bb3_and147_i = (local_bb3_shr95_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp92_i_stall_local;
wire local_bb3_cmp92_i;

assign local_bb3_cmp92_i = ((local_bb3_and91_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp89_i_stall_local;
wire local_bb3_cmp89_i;

assign local_bb3_cmp89_i = ((local_bb3_and88_i541 & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp86_i_stall_local;
wire local_bb3_cmp86_i;

assign local_bb3_cmp86_i = ((local_bb3_and85_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u31_stall_local;
wire local_bb3_var__u31;

assign local_bb3_var__u31 = ((local_bb3_var__u29 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__34_i369_stall_local;
wire [31:0] local_bb3__34_i369;

assign local_bb3__34_i369 = (local_bb3__31_i366 ? (local_bb3_or_i_i363 & 32'h1FFFFFF) : (local_bb3_or_i17_i355 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__33_i368_stall_local;
wire [31:0] local_bb3__33_i368;

assign local_bb3__33_i368 = (local_bb3_tobool49_i359 ? (local_bb3__32_i367 & 32'hFFFFFF00) : (local_bb3_shl1_i18_i356 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__37_i372_stall_local;
wire [31:0] local_bb3__37_i372;

assign local_bb3__37_i372 = (local_bb3_tobool49_i359 ? (local_bb3__36_i371 & 32'h1FF) : (local_bb3_inc_i360 & 32'h3FF));

// This section implements a registered operation.
// 
wire SFC_1_VALID_352_353_0_inputs_ready;
 reg SFC_1_VALID_352_353_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_352_353_0_stall_in;
wire SFC_1_VALID_352_353_0_output_regs_ready;
 reg SFC_1_VALID_352_353_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_352_353_0_causedstall;

assign SFC_1_VALID_352_353_0_inputs_ready = 1'b1;
assign SFC_1_VALID_352_353_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_351_352_0_stall_in = 1'b0;
assign SFC_1_VALID_352_353_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_352_353_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_352_353_0_output_regs_ready)
		begin
			SFC_1_VALID_352_353_0_NO_SHIFT_REG <= SFC_1_VALID_351_352_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_frombool75_i_stall_local;
wire [7:0] local_bb3_frombool75_i;

assign local_bb3_frombool75_i = (local_bb3_and73_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u32_stall_local;
wire [31:0] local_bb3_var__u32;

assign local_bb3_var__u32 = ((local_bb3_and147_i & 32'h3FFFFFFF) | local_bb3_shr95_i);

// This section implements an unregistered operation.
// 
wire local_bb3__31_v_i545_stall_local;
wire local_bb3__31_v_i545;

assign local_bb3__31_v_i545 = (local_bb3_cmp97_i ? local_bb3_cmp80_i : local_bb3_cmp92_i);

// This section implements an unregistered operation.
// 
wire local_bb3__30_v_i543_stall_local;
wire local_bb3__30_v_i543;

assign local_bb3__30_v_i543 = (local_bb3_cmp97_i ? local_bb3_cmp77_i540 : local_bb3_cmp89_i);

// This section implements an unregistered operation.
// 
wire local_bb3_frombool110_i_stall_local;
wire [7:0] local_bb3_frombool110_i;

assign local_bb3_frombool110_i[7:1] = 7'h0;
assign local_bb3_frombool110_i[0] = local_bb3_cmp86_i;

// This section implements an unregistered operation.
// 
wire local_bb3_or108_i_stall_local;
wire [31:0] local_bb3_or108_i;

assign local_bb3_or108_i[31:1] = 31'h0;
assign local_bb3_or108_i[0] = local_bb3_var__u31;

// This section implements an unregistered operation.
// 
wire local_bb3__35_i370_stall_local;
wire [31:0] local_bb3__35_i370;

assign local_bb3__35_i370 = (local_bb3_tobool49_i359 ? (local_bb3__34_i369 & 32'h1FFFFFF) : (local_bb3_or_i17_i355 & 32'hFFFFFF));

// This section implements a registered operation.
// 
wire SFC_1_VALID_353_354_0_inputs_ready;
 reg SFC_1_VALID_353_354_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_353_354_0_stall_in;
wire SFC_1_VALID_353_354_0_output_regs_ready;
 reg SFC_1_VALID_353_354_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_353_354_0_causedstall;

assign SFC_1_VALID_353_354_0_inputs_ready = 1'b1;
assign SFC_1_VALID_353_354_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_352_353_0_stall_in = 1'b0;
assign SFC_1_VALID_353_354_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_353_354_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_353_354_0_output_regs_ready)
		begin
			SFC_1_VALID_353_354_0_NO_SHIFT_REG <= SFC_1_VALID_352_353_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_or1606_i_stall_local;
wire [31:0] local_bb3_or1606_i;

assign local_bb3_or1606_i = (local_bb3_var__u32 | (local_bb3_and143_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__31_i546_stall_local;
wire [7:0] local_bb3__31_i546;

assign local_bb3__31_i546[7:1] = 7'h0;
assign local_bb3__31_i546[0] = local_bb3__31_v_i545;

// This section implements an unregistered operation.
// 
wire local_bb3__30_i544_stall_local;
wire [7:0] local_bb3__30_i544;

assign local_bb3__30_i544[7:1] = 7'h0;
assign local_bb3__30_i544[0] = local_bb3__30_v_i543;

// This section implements an unregistered operation.
// 
wire local_bb3__29_i542_stall_local;
wire [7:0] local_bb3__29_i542;

assign local_bb3__29_i542 = (local_bb3_cmp97_i ? (local_bb3_frombool75_i & 8'h1) : (local_bb3_frombool110_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__32_i547_stall_local;
wire [31:0] local_bb3__32_i547;

assign local_bb3__32_i547 = (local_bb3_cmp97_i ? 32'h0 : (local_bb3_or108_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and75_i378_stall_local;
wire [31:0] local_bb3_and75_i378;

assign local_bb3_and75_i378 = ((local_bb3__35_i370 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3__33_i368_valid_out;
wire local_bb3__33_i368_stall_in;
wire local_bb3__37_i372_valid_out;
wire local_bb3__37_i372_stall_in;
wire local_bb3_and75_i378_valid_out;
wire local_bb3_and75_i378_stall_in;
wire local_bb3_and83_i384_valid_out;
wire local_bb3_and83_i384_stall_in;
wire local_bb3_and83_i384_inputs_ready;
wire local_bb3_and83_i384_stall_local;
wire [31:0] local_bb3_and83_i384;

assign local_bb3_and83_i384_inputs_ready = (local_bb3_mul_i_i350_valid_out_0_NO_SHIFT_REG & local_bb3_mul_i_i350_valid_out_1_NO_SHIFT_REG & rnode_334to335_bb3_add_i357_0_valid_out_1_NO_SHIFT_REG & rnode_334to335_bb3_add_i357_0_valid_out_0_NO_SHIFT_REG & rnode_334to335_bb3_add_i357_0_valid_out_2_NO_SHIFT_REG);
assign local_bb3_and83_i384 = ((local_bb3__35_i370 & 32'h1FFFFFF) & 32'h1);
assign local_bb3__33_i368_valid_out = 1'b1;
assign local_bb3__37_i372_valid_out = 1'b1;
assign local_bb3_and75_i378_valid_out = 1'b1;
assign local_bb3_and83_i384_valid_out = 1'b1;
assign local_bb3_mul_i_i350_stall_in_0 = 1'b0;
assign local_bb3_mul_i_i350_stall_in_1 = 1'b0;
assign rnode_334to335_bb3_add_i357_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_add_i357_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_add_i357_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_354_355_0_inputs_ready;
 reg SFC_1_VALID_354_355_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_354_355_0_stall_in;
wire SFC_1_VALID_354_355_0_output_regs_ready;
 reg SFC_1_VALID_354_355_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_354_355_0_causedstall;

assign SFC_1_VALID_354_355_0_inputs_ready = 1'b1;
assign SFC_1_VALID_354_355_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_353_354_0_stall_in = 1'b0;
assign SFC_1_VALID_354_355_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_354_355_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_354_355_0_output_regs_ready)
		begin
			SFC_1_VALID_354_355_0_NO_SHIFT_REG <= SFC_1_VALID_353_354_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_or163_i_stall_local;
wire [31:0] local_bb3_or163_i;

assign local_bb3_or163_i = (local_bb3_or1606_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or1247_i_stall_local;
wire [7:0] local_bb3_or1247_i;

assign local_bb3_or1247_i = ((local_bb3__30_i544 & 8'h1) | (local_bb3__29_i542 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__33_i549_stall_local;
wire [7:0] local_bb3__33_i549;

assign local_bb3__33_i549 = (local_bb3_cmp117_i ? (local_bb3__29_i542 & 8'h1) : (local_bb3__31_i546 & 8'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_335to336_bb3__33_i368_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3__33_i368_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__33_i368_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3__33_i368_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_335to336_bb3__33_i368_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__33_i368_1_NO_SHIFT_REG;
 logic rnode_335to336_bb3__33_i368_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__33_i368_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__33_i368_0_valid_out_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__33_i368_0_stall_in_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__33_i368_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_335to336_bb3__33_i368_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to336_bb3__33_i368_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to336_bb3__33_i368_0_stall_in_0_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_335to336_bb3__33_i368_0_valid_out_0_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_335to336_bb3__33_i368_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in((local_bb3__33_i368 & 32'hFFFFFF00)),
	.data_out(rnode_335to336_bb3__33_i368_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_335to336_bb3__33_i368_0_reg_336_fifo.DEPTH = 1;
defparam rnode_335to336_bb3__33_i368_0_reg_336_fifo.DATA_WIDTH = 32;
defparam rnode_335to336_bb3__33_i368_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to336_bb3__33_i368_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_335to336_bb3__33_i368_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__33_i368_stall_in = 1'b0;
assign rnode_335to336_bb3__33_i368_0_stall_in_0_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3__33_i368_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3__33_i368_0_NO_SHIFT_REG = rnode_335to336_bb3__33_i368_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3__33_i368_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3__33_i368_1_NO_SHIFT_REG = rnode_335to336_bb3__33_i368_0_reg_336_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_335to336_bb3__37_i372_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__37_i372_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__37_i372_1_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__37_i372_2_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__37_i372_3_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3__37_i372_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_valid_out_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_stall_in_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__37_i372_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_335to336_bb3__37_i372_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to336_bb3__37_i372_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to336_bb3__37_i372_0_stall_in_0_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_335to336_bb3__37_i372_0_valid_out_0_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_335to336_bb3__37_i372_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in((local_bb3__37_i372 & 32'h3FF)),
	.data_out(rnode_335to336_bb3__37_i372_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_335to336_bb3__37_i372_0_reg_336_fifo.DEPTH = 1;
defparam rnode_335to336_bb3__37_i372_0_reg_336_fifo.DATA_WIDTH = 32;
defparam rnode_335to336_bb3__37_i372_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to336_bb3__37_i372_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_335to336_bb3__37_i372_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__37_i372_stall_in = 1'b0;
assign rnode_335to336_bb3__37_i372_0_stall_in_0_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3__37_i372_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3__37_i372_0_NO_SHIFT_REG = rnode_335to336_bb3__37_i372_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3__37_i372_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3__37_i372_1_NO_SHIFT_REG = rnode_335to336_bb3__37_i372_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3__37_i372_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3__37_i372_2_NO_SHIFT_REG = rnode_335to336_bb3__37_i372_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3__37_i372_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3__37_i372_3_NO_SHIFT_REG = rnode_335to336_bb3__37_i372_0_reg_336_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_335to337_bb3_and75_i378_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and75_i378_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_and75_i378_0_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and75_i378_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_and75_i378_0_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and75_i378_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and75_i378_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and75_i378_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_335to337_bb3_and75_i378_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to337_bb3_and75_i378_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to337_bb3_and75_i378_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_335to337_bb3_and75_i378_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_335to337_bb3_and75_i378_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((local_bb3_and75_i378 & 32'h7FFFFF)),
	.data_out(rnode_335to337_bb3_and75_i378_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_335to337_bb3_and75_i378_0_reg_337_fifo.DEPTH = 2;
defparam rnode_335to337_bb3_and75_i378_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_335to337_bb3_and75_i378_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to337_bb3_and75_i378_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_335to337_bb3_and75_i378_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and75_i378_stall_in = 1'b0;
assign rnode_335to337_bb3_and75_i378_0_NO_SHIFT_REG = rnode_335to337_bb3_and75_i378_0_reg_337_NO_SHIFT_REG;
assign rnode_335to337_bb3_and75_i378_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_and75_i378_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_335to336_bb3_and83_i384_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to336_bb3_and83_i384_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3_and83_i384_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3_and83_i384_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3_and83_i384_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_and83_i384_0_valid_out_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_and83_i384_0_stall_in_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_and83_i384_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_335to336_bb3_and83_i384_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to336_bb3_and83_i384_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to336_bb3_and83_i384_0_stall_in_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_335to336_bb3_and83_i384_0_valid_out_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_335to336_bb3_and83_i384_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in((local_bb3_and83_i384 & 32'h1)),
	.data_out(rnode_335to336_bb3_and83_i384_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_335to336_bb3_and83_i384_0_reg_336_fifo.DEPTH = 1;
defparam rnode_335to336_bb3_and83_i384_0_reg_336_fifo.DATA_WIDTH = 32;
defparam rnode_335to336_bb3_and83_i384_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to336_bb3_and83_i384_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_335to336_bb3_and83_i384_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and83_i384_stall_in = 1'b0;
assign rnode_335to336_bb3_and83_i384_0_NO_SHIFT_REG = rnode_335to336_bb3_and83_i384_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3_and83_i384_0_stall_in_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3_and83_i384_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_355_356_0_inputs_ready;
 reg SFC_1_VALID_355_356_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_355_356_0_stall_in;
wire SFC_1_VALID_355_356_0_output_regs_ready;
 reg SFC_1_VALID_355_356_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_355_356_0_causedstall;

assign SFC_1_VALID_355_356_0_inputs_ready = 1'b1;
assign SFC_1_VALID_355_356_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_354_355_0_stall_in = 1'b0;
assign SFC_1_VALID_355_356_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_355_356_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_355_356_0_output_regs_ready)
		begin
			SFC_1_VALID_355_356_0_NO_SHIFT_REG <= SFC_1_VALID_354_355_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__37_v_i552_stall_local;
wire [31:0] local_bb3__37_v_i552;

assign local_bb3__37_v_i552 = (local_bb3_Pivot20_i550 ? 32'h0 : (local_bb3_or163_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or124_i548_stall_local;
wire [31:0] local_bb3_or124_i548;

assign local_bb3_or124_i548[31:8] = 24'h0;
assign local_bb3_or124_i548[7:0] = (local_bb3_or1247_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u33_stall_local;
wire [7:0] local_bb3_var__u33;

assign local_bb3_var__u33 = ((local_bb3__33_i549 & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp77_i383_stall_local;
wire local_bb3_cmp77_i383;

assign local_bb3_cmp77_i383 = ((rnode_335to336_bb3__33_i368_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u34_stall_local;
wire local_bb3_var__u34;

assign local_bb3_var__u34 = ($signed((rnode_335to336_bb3__33_i368_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp53_i373_stall_local;
wire local_bb3_cmp53_i373;

assign local_bb3_cmp53_i373 = ((rnode_335to336_bb3__37_i372_0_NO_SHIFT_REG & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp68_i377_valid_out;
wire local_bb3_cmp68_i377_stall_in;
wire local_bb3_cmp68_i377_inputs_ready;
wire local_bb3_cmp68_i377_stall_local;
wire local_bb3_cmp68_i377;

assign local_bb3_cmp68_i377_inputs_ready = rnode_335to336_bb3__37_i372_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_cmp68_i377 = ((rnode_335to336_bb3__37_i372_1_NO_SHIFT_REG & 32'h3FF) < 32'h80);
assign local_bb3_cmp68_i377_valid_out = 1'b1;
assign rnode_335to336_bb3__37_i372_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_sub_i379_stall_local;
wire [31:0] local_bb3_sub_i379;

assign local_bb3_sub_i379 = ((rnode_335to336_bb3__37_i372_2_NO_SHIFT_REG & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp71_not_i394_valid_out;
wire local_bb3_cmp71_not_i394_stall_in;
wire local_bb3_cmp71_not_i394_inputs_ready;
wire local_bb3_cmp71_not_i394_stall_local;
wire local_bb3_cmp71_not_i394;

assign local_bb3_cmp71_not_i394_inputs_ready = rnode_335to336_bb3__37_i372_0_valid_out_3_NO_SHIFT_REG;
assign local_bb3_cmp71_not_i394 = ((rnode_335to336_bb3__37_i372_3_NO_SHIFT_REG & 32'h3FF) != 32'h7F);
assign local_bb3_cmp71_not_i394_valid_out = 1'b1;
assign rnode_335to336_bb3__37_i372_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_tobool84_i385_stall_local;
wire local_bb3_tobool84_i385;

assign local_bb3_tobool84_i385 = ((rnode_335to336_bb3_and83_i384_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements a registered operation.
// 
wire SFC_1_VALID_356_357_0_inputs_ready;
 reg SFC_1_VALID_356_357_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_356_357_0_stall_in;
wire SFC_1_VALID_356_357_0_output_regs_ready;
 reg SFC_1_VALID_356_357_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_356_357_0_causedstall;

assign SFC_1_VALID_356_357_0_inputs_ready = 1'b1;
assign SFC_1_VALID_356_357_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_355_356_0_stall_in = 1'b0;
assign SFC_1_VALID_356_357_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_356_357_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_356_357_0_output_regs_ready)
		begin
			SFC_1_VALID_356_357_0_NO_SHIFT_REG <= SFC_1_VALID_355_356_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__39_v_i553_stall_local;
wire [31:0] local_bb3__39_v_i553;

assign local_bb3__39_v_i553 = (local_bb3_SwitchLeaf_i551 ? (local_bb3_var__u30 & 32'h1) : (local_bb3__37_v_i552 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or125_i_stall_local;
wire [31:0] local_bb3_or125_i;

assign local_bb3_or125_i = (local_bb3_cmp117_i ? 32'h0 : (local_bb3_or124_i548 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_conv136_i_stall_local;
wire [31:0] local_bb3_conv136_i;

assign local_bb3_conv136_i[31:8] = 24'h0;
assign local_bb3_conv136_i[7:0] = (local_bb3_var__u33 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or581_i374_valid_out;
wire local_bb3_or581_i374_stall_in;
wire local_bb3_or581_i374_inputs_ready;
wire local_bb3_or581_i374_stall_local;
wire local_bb3_or581_i374;

assign local_bb3_or581_i374_inputs_ready = (rnode_335to336_bb3_var__u23_0_valid_out_NO_SHIFT_REG & rnode_335to336_bb3__37_i372_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3_or581_i374 = (rnode_335to336_bb3_var__u23_0_NO_SHIFT_REG | local_bb3_cmp53_i373);
assign local_bb3_or581_i374_valid_out = 1'b1;
assign rnode_335to336_bb3_var__u23_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3__37_i372_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_cmp68_i377_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp68_i377_0_stall_in_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp68_i377_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp68_i377_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp68_i377_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp68_i377_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp68_i377_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp68_i377_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_cmp68_i377_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_cmp68_i377_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_cmp68_i377_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_cmp68_i377_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_cmp68_i377_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(local_bb3_cmp68_i377),
	.data_out(rnode_336to337_bb3_cmp68_i377_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_cmp68_i377_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_cmp68_i377_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_336to337_bb3_cmp68_i377_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_cmp68_i377_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_cmp68_i377_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp68_i377_stall_in = 1'b0;
assign rnode_336to337_bb3_cmp68_i377_0_NO_SHIFT_REG = rnode_336to337_bb3_cmp68_i377_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_cmp68_i377_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_cmp68_i377_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and74_i380_stall_local;
wire [31:0] local_bb3_and74_i380;

assign local_bb3_and74_i380 = ((local_bb3_sub_i379 & 32'hFF800000) + 32'h40800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_cmp71_not_i394_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp71_not_i394_0_stall_in_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp71_not_i394_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp71_not_i394_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp71_not_i394_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp71_not_i394_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp71_not_i394_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_cmp71_not_i394_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_cmp71_not_i394_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_cmp71_not_i394_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_cmp71_not_i394_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_cmp71_not_i394_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_cmp71_not_i394_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(local_bb3_cmp71_not_i394),
	.data_out(rnode_336to337_bb3_cmp71_not_i394_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_cmp71_not_i394_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_cmp71_not_i394_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_336to337_bb3_cmp71_not_i394_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_cmp71_not_i394_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_cmp71_not_i394_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp71_not_i394_stall_in = 1'b0;
assign rnode_336to337_bb3_cmp71_not_i394_0_NO_SHIFT_REG = rnode_336to337_bb3_cmp71_not_i394_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_cmp71_not_i394_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_cmp71_not_i394_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__39_i386_stall_local;
wire local_bb3__39_i386;

assign local_bb3__39_i386 = (local_bb3_tobool84_i385 & local_bb3_var__u34);

// This section implements a registered operation.
// 
wire SFC_1_VALID_357_358_0_inputs_ready;
 reg SFC_1_VALID_357_358_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_357_358_0_stall_in;
wire SFC_1_VALID_357_358_0_output_regs_ready;
 reg SFC_1_VALID_357_358_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_357_358_0_causedstall;

assign SFC_1_VALID_357_358_0_inputs_ready = 1'b1;
assign SFC_1_VALID_357_358_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_356_357_0_stall_in = 1'b0;
assign SFC_1_VALID_357_358_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_357_358_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_357_358_0_output_regs_ready)
		begin
			SFC_1_VALID_357_358_0_NO_SHIFT_REG <= SFC_1_VALID_356_357_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_reduction_3_i554_stall_local;
wire [31:0] local_bb3_reduction_3_i554;

assign local_bb3_reduction_3_i554 = ((local_bb3__32_i547 & 32'h1) | (local_bb3_or125_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or137_i_stall_local;
wire [31:0] local_bb3_or137_i;

assign local_bb3_or137_i = (local_bb3_cmp132_not_i ? (local_bb3_conv136_i & 32'h1) : 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_or581_i374_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_1_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_valid_out_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_stall_in_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_or581_i374_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_or581_i374_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_or581_i374_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_or581_i374_0_stall_in_0_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_or581_i374_0_valid_out_0_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_or581_i374_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(local_bb3_or581_i374),
	.data_out(rnode_336to337_bb3_or581_i374_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_or581_i374_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_or581_i374_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_336to337_bb3_or581_i374_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_or581_i374_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_or581_i374_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or581_i374_stall_in = 1'b0;
assign rnode_336to337_bb3_or581_i374_0_stall_in_0_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_or581_i374_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3_or581_i374_0_NO_SHIFT_REG = rnode_336to337_bb3_or581_i374_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_or581_i374_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3_or581_i374_1_NO_SHIFT_REG = rnode_336to337_bb3_or581_i374_0_reg_337_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u35_stall_local;
wire [31:0] local_bb3_var__u35;

assign local_bb3_var__u35[31:1] = 31'h0;
assign local_bb3_var__u35[0] = rnode_336to337_bb3_cmp68_i377_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i381_valid_out;
wire local_bb3_shl_i381_stall_in;
wire local_bb3_shl_i381_inputs_ready;
wire local_bb3_shl_i381_stall_local;
wire [31:0] local_bb3_shl_i381;

assign local_bb3_shl_i381_inputs_ready = rnode_335to336_bb3__37_i372_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_shl_i381 = ((local_bb3_and74_i380 & 32'hFF800000) & 32'h7F800000);
assign local_bb3_shl_i381_valid_out = 1'b1;
assign rnode_335to336_bb3__37_i372_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__40_i387_valid_out;
wire local_bb3__40_i387_stall_in;
wire local_bb3__40_i387_inputs_ready;
wire local_bb3__40_i387_stall_local;
wire local_bb3__40_i387;

assign local_bb3__40_i387_inputs_ready = (rnode_335to336_bb3__33_i368_0_valid_out_0_NO_SHIFT_REG & rnode_335to336_bb3__33_i368_0_valid_out_1_NO_SHIFT_REG & rnode_335to336_bb3_and83_i384_0_valid_out_NO_SHIFT_REG);
assign local_bb3__40_i387 = (local_bb3_cmp77_i383 | local_bb3__39_i386);
assign local_bb3__40_i387_valid_out = 1'b1;
assign rnode_335to336_bb3__33_i368_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3__33_i368_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3_and83_i384_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_358_359_0_inputs_ready;
 reg SFC_1_VALID_358_359_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_358_359_0_stall_in;
wire SFC_1_VALID_358_359_0_output_regs_ready;
 reg SFC_1_VALID_358_359_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_358_359_0_causedstall;

assign SFC_1_VALID_358_359_0_inputs_ready = 1'b1;
assign SFC_1_VALID_358_359_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_357_358_0_stall_in = 1'b0;
assign SFC_1_VALID_358_359_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_358_359_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_358_359_0_output_regs_ready)
		begin
			SFC_1_VALID_358_359_0_NO_SHIFT_REG <= SFC_1_VALID_357_358_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_reduction_5_i556_stall_local;
wire [31:0] local_bb3_reduction_5_i556;

assign local_bb3_reduction_5_i556 = (local_bb3_shr151_i | (local_bb3_reduction_3_i554 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_4_i555_stall_local;
wire [31:0] local_bb3_reduction_4_i555;

assign local_bb3_reduction_4_i555 = ((local_bb3_or137_i & 32'h1) | (local_bb3__39_v_i553 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_2_i376_stall_local;
wire local_bb3_reduction_2_i376;

assign local_bb3_reduction_2_i376 = (rnode_336to337_bb3_reduction_0_i375_0_NO_SHIFT_REG | rnode_336to337_bb3_or581_i374_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_cond111_i402_stall_local;
wire [31:0] local_bb3_cond111_i402;

assign local_bb3_cond111_i402 = (rnode_336to337_bb3_or581_i374_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_shl_i381_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_shl_i381_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_shl_i381_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_shl_i381_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_shl_i381_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_shl_i381_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_shl_i381_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_shl_i381_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_shl_i381_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_shl_i381_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_shl_i381_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_shl_i381_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_shl_i381_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((local_bb3_shl_i381 & 32'h7F800000)),
	.data_out(rnode_336to337_bb3_shl_i381_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_shl_i381_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_shl_i381_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_336to337_bb3_shl_i381_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_shl_i381_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_shl_i381_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shl_i381_stall_in = 1'b0;
assign rnode_336to337_bb3_shl_i381_0_NO_SHIFT_REG = rnode_336to337_bb3_shl_i381_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_shl_i381_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_shl_i381_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3__40_i387_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3__40_i387_0_stall_in_NO_SHIFT_REG;
 logic rnode_336to337_bb3__40_i387_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3__40_i387_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to337_bb3__40_i387_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__40_i387_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__40_i387_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__40_i387_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3__40_i387_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3__40_i387_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3__40_i387_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3__40_i387_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3__40_i387_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(local_bb3__40_i387),
	.data_out(rnode_336to337_bb3__40_i387_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3__40_i387_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3__40_i387_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_336to337_bb3__40_i387_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3__40_i387_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3__40_i387_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__40_i387_stall_in = 1'b0;
assign rnode_336to337_bb3__40_i387_0_NO_SHIFT_REG = rnode_336to337_bb3__40_i387_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3__40_i387_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__40_i387_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_359_360_0_inputs_ready;
 reg SFC_1_VALID_359_360_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_359_360_0_stall_in;
wire SFC_1_VALID_359_360_0_output_regs_ready;
 reg SFC_1_VALID_359_360_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_359_360_0_causedstall;

assign SFC_1_VALID_359_360_0_inputs_ready = 1'b1;
assign SFC_1_VALID_359_360_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_358_359_0_stall_in = 1'b0;
assign SFC_1_VALID_359_360_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_359_360_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_359_360_0_output_regs_ready)
		begin
			SFC_1_VALID_359_360_0_NO_SHIFT_REG <= SFC_1_VALID_358_359_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_reduction_6_i557_stall_local;
wire [31:0] local_bb3_reduction_6_i557;

assign local_bb3_reduction_6_i557 = ((local_bb3_reduction_4_i555 & 32'h1) | local_bb3_reduction_5_i556);

// This section implements an unregistered operation.
// 
wire local_bb3_conv101_i397_stall_local;
wire [31:0] local_bb3_conv101_i397;

assign local_bb3_conv101_i397[31:1] = 31'h0;
assign local_bb3_conv101_i397[0] = local_bb3_reduction_2_i376;

// This section implements an unregistered operation.
// 
wire local_bb3_or76_i382_stall_local;
wire [31:0] local_bb3_or76_i382;

assign local_bb3_or76_i382 = ((rnode_336to337_bb3_shl_i381_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_335to337_bb3_and75_i378_0_NO_SHIFT_REG & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cond_i388_stall_local;
wire [31:0] local_bb3_cond_i388;

assign local_bb3_cond_i388[31:1] = 31'h0;
assign local_bb3_cond_i388[0] = rnode_336to337_bb3__40_i387_0_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_1_VALID_360_361_0_inputs_ready;
 reg SFC_1_VALID_360_361_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_360_361_0_stall_in;
wire SFC_1_VALID_360_361_0_output_regs_ready;
 reg SFC_1_VALID_360_361_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_360_361_0_causedstall;

assign SFC_1_VALID_360_361_0_inputs_ready = 1'b1;
assign SFC_1_VALID_360_361_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_359_360_0_stall_in = 1'b0;
assign SFC_1_VALID_360_361_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_360_361_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_360_361_0_output_regs_ready)
		begin
			SFC_1_VALID_360_361_0_NO_SHIFT_REG <= SFC_1_VALID_359_360_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_lnot33_not_i524_valid_out;
wire local_bb3_lnot33_not_i524_stall_in;
wire local_bb3_cmp38_i_valid_out;
wire local_bb3_cmp38_i_stall_in;
wire local_bb3_and37_lobit_i_valid_out;
wire local_bb3_and37_lobit_i_stall_in;
wire local_bb3_xor189_i_valid_out;
wire local_bb3_xor189_i_stall_in;
wire local_bb3_xor189_i_inputs_ready;
wire local_bb3_xor189_i_stall_local;
wire [31:0] local_bb3_xor189_i;

assign local_bb3_xor189_i_inputs_ready = (rnode_333to334_bb3__22_i508_0_valid_out_0_NO_SHIFT_REG & rnode_333to334_bb3_lnot23_i517_0_valid_out_NO_SHIFT_REG & rnode_333to334_bb3_align_0_i539_0_valid_out_0_NO_SHIFT_REG & rnode_333to334_bb3_align_0_i539_0_valid_out_4_NO_SHIFT_REG & rnode_333to334_bb3_align_0_i539_0_valid_out_1_NO_SHIFT_REG & rnode_333to334_bb3_align_0_i539_0_valid_out_2_NO_SHIFT_REG & rnode_333to334_bb3_align_0_i539_0_valid_out_3_NO_SHIFT_REG & rnode_333to334_bb3__23_i509_0_valid_out_2_NO_SHIFT_REG & rnode_333to334_bb3__22_i508_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_xor189_i = (local_bb3_reduction_6_i557 ^ local_bb3_xor36_lobit_i);
assign local_bb3_lnot33_not_i524_valid_out = 1'b1;
assign local_bb3_cmp38_i_valid_out = 1'b1;
assign local_bb3_and37_lobit_i_valid_out = 1'b1;
assign local_bb3_xor189_i_valid_out = 1'b1;
assign rnode_333to334_bb3__22_i508_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_lnot23_i517_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_align_0_i539_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_align_0_i539_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_align_0_i539_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_align_0_i539_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3_align_0_i539_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3__23_i509_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_333to334_bb3__22_i508_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_add87_i389_stall_local;
wire [31:0] local_bb3_add87_i389;

assign local_bb3_add87_i389 = ((local_bb3_cond_i388 & 32'h1) + (local_bb3_or76_i382 & 32'h7FFFFFFF));

// This section implements a registered operation.
// 
wire SFC_1_VALID_361_362_0_inputs_ready;
 reg SFC_1_VALID_361_362_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_361_362_0_stall_in;
wire SFC_1_VALID_361_362_0_output_regs_ready;
 reg SFC_1_VALID_361_362_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_361_362_0_causedstall;

assign SFC_1_VALID_361_362_0_inputs_ready = 1'b1;
assign SFC_1_VALID_361_362_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_360_361_0_stall_in = 1'b0;
assign SFC_1_VALID_361_362_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_361_362_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_361_362_0_output_regs_ready)
		begin
			SFC_1_VALID_361_362_0_NO_SHIFT_REG <= SFC_1_VALID_360_361_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_334to335_bb3_lnot33_not_i524_0_valid_out_NO_SHIFT_REG;
 logic rnode_334to335_bb3_lnot33_not_i524_0_stall_in_NO_SHIFT_REG;
 logic rnode_334to335_bb3_lnot33_not_i524_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_lnot33_not_i524_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic rnode_334to335_bb3_lnot33_not_i524_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_lnot33_not_i524_0_valid_out_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_lnot33_not_i524_0_stall_in_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_lnot33_not_i524_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_334to335_bb3_lnot33_not_i524_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_334to335_bb3_lnot33_not_i524_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_334to335_bb3_lnot33_not_i524_0_stall_in_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_334to335_bb3_lnot33_not_i524_0_valid_out_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_334to335_bb3_lnot33_not_i524_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in(local_bb3_lnot33_not_i524),
	.data_out(rnode_334to335_bb3_lnot33_not_i524_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_334to335_bb3_lnot33_not_i524_0_reg_335_fifo.DEPTH = 1;
defparam rnode_334to335_bb3_lnot33_not_i524_0_reg_335_fifo.DATA_WIDTH = 1;
defparam rnode_334to335_bb3_lnot33_not_i524_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_334to335_bb3_lnot33_not_i524_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_334to335_bb3_lnot33_not_i524_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_lnot33_not_i524_stall_in = 1'b0;
assign rnode_334to335_bb3_lnot33_not_i524_0_NO_SHIFT_REG = rnode_334to335_bb3_lnot33_not_i524_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_lnot33_not_i524_0_stall_in_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_lnot33_not_i524_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_334to335_bb3_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_valid_out_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_stall_in_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_cmp38_i_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_334to335_bb3_cmp38_i_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_334to335_bb3_cmp38_i_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_334to335_bb3_cmp38_i_0_stall_in_0_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_334to335_bb3_cmp38_i_0_valid_out_0_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_334to335_bb3_cmp38_i_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in(local_bb3_cmp38_i),
	.data_out(rnode_334to335_bb3_cmp38_i_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_334to335_bb3_cmp38_i_0_reg_335_fifo.DEPTH = 1;
defparam rnode_334to335_bb3_cmp38_i_0_reg_335_fifo.DATA_WIDTH = 1;
defparam rnode_334to335_bb3_cmp38_i_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_334to335_bb3_cmp38_i_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_334to335_bb3_cmp38_i_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp38_i_stall_in = 1'b0;
assign rnode_334to335_bb3_cmp38_i_0_stall_in_0_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_cmp38_i_0_NO_SHIFT_REG = rnode_334to335_bb3_cmp38_i_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_cmp38_i_1_NO_SHIFT_REG = rnode_334to335_bb3_cmp38_i_0_reg_335_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_334to335_bb3_and37_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and37_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_and37_lobit_i_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and37_lobit_i_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_and37_lobit_i_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and37_lobit_i_0_valid_out_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and37_lobit_i_0_stall_in_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_and37_lobit_i_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_334to335_bb3_and37_lobit_i_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_334to335_bb3_and37_lobit_i_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_334to335_bb3_and37_lobit_i_0_stall_in_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_334to335_bb3_and37_lobit_i_0_valid_out_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_334to335_bb3_and37_lobit_i_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in((local_bb3_and37_lobit_i & 32'h1)),
	.data_out(rnode_334to335_bb3_and37_lobit_i_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_334to335_bb3_and37_lobit_i_0_reg_335_fifo.DEPTH = 1;
defparam rnode_334to335_bb3_and37_lobit_i_0_reg_335_fifo.DATA_WIDTH = 32;
defparam rnode_334to335_bb3_and37_lobit_i_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_334to335_bb3_and37_lobit_i_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_334to335_bb3_and37_lobit_i_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and37_lobit_i_stall_in = 1'b0;
assign rnode_334to335_bb3_and37_lobit_i_0_NO_SHIFT_REG = rnode_334to335_bb3_and37_lobit_i_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_and37_lobit_i_0_stall_in_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_and37_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_334to335_bb3_xor189_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_334to335_bb3_xor189_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_xor189_i_0_NO_SHIFT_REG;
 logic rnode_334to335_bb3_xor189_i_0_reg_335_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_334to335_bb3_xor189_i_0_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_xor189_i_0_valid_out_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_xor189_i_0_stall_in_reg_335_NO_SHIFT_REG;
 logic rnode_334to335_bb3_xor189_i_0_stall_out_reg_335_NO_SHIFT_REG;

acl_data_fifo rnode_334to335_bb3_xor189_i_0_reg_335_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_334to335_bb3_xor189_i_0_reg_335_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_334to335_bb3_xor189_i_0_stall_in_reg_335_NO_SHIFT_REG),
	.valid_out(rnode_334to335_bb3_xor189_i_0_valid_out_reg_335_NO_SHIFT_REG),
	.stall_out(rnode_334to335_bb3_xor189_i_0_stall_out_reg_335_NO_SHIFT_REG),
	.data_in(local_bb3_xor189_i),
	.data_out(rnode_334to335_bb3_xor189_i_0_reg_335_NO_SHIFT_REG)
);

defparam rnode_334to335_bb3_xor189_i_0_reg_335_fifo.DEPTH = 1;
defparam rnode_334to335_bb3_xor189_i_0_reg_335_fifo.DATA_WIDTH = 32;
defparam rnode_334to335_bb3_xor189_i_0_reg_335_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_334to335_bb3_xor189_i_0_reg_335_fifo.IMPL = "shift_reg";

assign rnode_334to335_bb3_xor189_i_0_reg_335_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_xor189_i_stall_in = 1'b0;
assign rnode_334to335_bb3_xor189_i_0_NO_SHIFT_REG = rnode_334to335_bb3_xor189_i_0_reg_335_NO_SHIFT_REG;
assign rnode_334to335_bb3_xor189_i_0_stall_in_reg_335_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_xor189_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and88_i390_stall_local;
wire [31:0] local_bb3_and88_i390;

assign local_bb3_and88_i390 = (local_bb3_add87_i389 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and90_i392_stall_local;
wire [31:0] local_bb3_and90_i392;

assign local_bb3_and90_i392 = (local_bb3_add87_i389 & 32'h800000);

// This section implements a registered operation.
// 
wire SFC_1_VALID_362_363_0_inputs_ready;
 reg SFC_1_VALID_362_363_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_362_363_0_stall_in;
wire SFC_1_VALID_362_363_0_output_regs_ready;
 reg SFC_1_VALID_362_363_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_362_363_0_causedstall;

assign SFC_1_VALID_362_363_0_inputs_ready = 1'b1;
assign SFC_1_VALID_362_363_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_361_362_0_stall_in = 1'b0;
assign SFC_1_VALID_362_363_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_362_363_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_362_363_0_output_regs_ready)
		begin
			SFC_1_VALID_362_363_0_NO_SHIFT_REG <= SFC_1_VALID_361_362_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_brmerge_not_i525_stall_local;
wire local_bb3_brmerge_not_i525;

assign local_bb3_brmerge_not_i525 = (rnode_333to335_bb3_cmp27_i519_0_NO_SHIFT_REG & rnode_334to335_bb3_lnot33_not_i524_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_335to337_bb3_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_2_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_valid_out_0_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_stall_in_0_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_cmp38_i_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_335to337_bb3_cmp38_i_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to337_bb3_cmp38_i_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to337_bb3_cmp38_i_0_stall_in_0_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_335to337_bb3_cmp38_i_0_valid_out_0_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_335to337_bb3_cmp38_i_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(rnode_334to335_bb3_cmp38_i_1_NO_SHIFT_REG),
	.data_out(rnode_335to337_bb3_cmp38_i_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_335to337_bb3_cmp38_i_0_reg_337_fifo.DEPTH = 2;
defparam rnode_335to337_bb3_cmp38_i_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_335to337_bb3_cmp38_i_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to337_bb3_cmp38_i_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_335to337_bb3_cmp38_i_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_334to335_bb3_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_cmp38_i_0_stall_in_0_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_335to337_bb3_cmp38_i_0_NO_SHIFT_REG = rnode_335to337_bb3_cmp38_i_0_reg_337_NO_SHIFT_REG;
assign rnode_335to337_bb3_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_335to337_bb3_cmp38_i_1_NO_SHIFT_REG = rnode_335to337_bb3_cmp38_i_0_reg_337_NO_SHIFT_REG;
assign rnode_335to337_bb3_cmp38_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_335to337_bb3_cmp38_i_2_NO_SHIFT_REG = rnode_335to337_bb3_cmp38_i_0_reg_337_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_add_i558_stall_local;
wire [31:0] local_bb3_add_i558;

assign local_bb3_add_i558 = ((local_bb3__27_i536 & 32'h7FFFFF8) | (rnode_334to335_bb3_and37_lobit_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or89_i391_stall_local;
wire [31:0] local_bb3_or89_i391;

assign local_bb3_or89_i391 = ((local_bb3_and88_i390 & 32'h7FFFFFFF) | (local_bb3_and4_i317 & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp91_i393_stall_local;
wire local_bb3_cmp91_i393;

assign local_bb3_cmp91_i393 = ((local_bb3_and90_i392 & 32'h800000) == 32'h0);

// This section implements a registered operation.
// 
wire SFC_1_VALID_363_364_0_inputs_ready;
 reg SFC_1_VALID_363_364_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_363_364_0_stall_in;
wire SFC_1_VALID_363_364_0_output_regs_ready;
 reg SFC_1_VALID_363_364_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_363_364_0_causedstall;

assign SFC_1_VALID_363_364_0_inputs_ready = 1'b1;
assign SFC_1_VALID_363_364_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_362_363_0_stall_in = 1'b0;
assign SFC_1_VALID_363_364_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_363_364_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_363_364_0_output_regs_ready)
		begin
			SFC_1_VALID_363_364_0_NO_SHIFT_REG <= SFC_1_VALID_362_363_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__24_i528_stall_local;
wire local_bb3__24_i528;

assign local_bb3__24_i528 = (local_bb3_or_cond_not_i527 | local_bb3_brmerge_not_i525);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge_not_not_i529_stall_local;
wire local_bb3_brmerge_not_not_i529;

assign local_bb3_brmerge_not_not_i529 = (local_bb3_brmerge_not_i525 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_not_cmp38_i_stall_local;
wire local_bb3_not_cmp38_i;

assign local_bb3_not_cmp38_i = (rnode_335to337_bb3_cmp38_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_add193_i_stall_local;
wire [31:0] local_bb3_add193_i;

assign local_bb3_add193_i = ((local_bb3_add_i558 & 32'h7FFFFF9) + rnode_334to335_bb3_xor189_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge14_i395_stall_local;
wire local_bb3_brmerge14_i395;

assign local_bb3_brmerge14_i395 = (local_bb3_cmp91_i393 | rnode_336to337_bb3_cmp71_not_i394_0_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_1_VALID_364_365_0_inputs_ready;
 reg SFC_1_VALID_364_365_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_364_365_0_stall_in;
wire SFC_1_VALID_364_365_0_output_regs_ready;
 reg SFC_1_VALID_364_365_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_364_365_0_causedstall;

assign SFC_1_VALID_364_365_0_inputs_ready = 1'b1;
assign SFC_1_VALID_364_365_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_363_364_0_stall_in = 1'b0;
assign SFC_1_VALID_364_365_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_364_365_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_364_365_0_output_regs_ready)
		begin
			SFC_1_VALID_364_365_0_NO_SHIFT_REG <= SFC_1_VALID_363_364_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_reduction_7_i530_stall_local;
wire local_bb3_reduction_7_i530;

assign local_bb3_reduction_7_i530 = (local_bb3_cmp25_i518 & local_bb3_brmerge_not_not_i529);

// This section implements an unregistered operation.
// 
wire local_bb3_conv99_i396_stall_local;
wire [31:0] local_bb3_conv99_i396;

assign local_bb3_conv99_i396 = (local_bb3_brmerge14_i395 ? (local_bb3_var__u35 & 32'h1) : 32'h0);

// This section implements a registered operation.
// 
wire SFC_1_VALID_365_366_0_inputs_ready;
 reg SFC_1_VALID_365_366_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_365_366_0_stall_in;
wire SFC_1_VALID_365_366_0_output_regs_ready;
 reg SFC_1_VALID_365_366_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_365_366_0_causedstall;

assign SFC_1_VALID_365_366_0_inputs_ready = 1'b1;
assign SFC_1_VALID_365_366_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_364_365_0_stall_in = 1'b0;
assign SFC_1_VALID_365_366_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_365_366_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_365_366_0_output_regs_ready)
		begin
			SFC_1_VALID_365_366_0_NO_SHIFT_REG <= SFC_1_VALID_364_365_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_reduction_9_i532_stall_local;
wire local_bb3_reduction_9_i532;

assign local_bb3_reduction_9_i532 = (local_bb3_reduction_7_i530 & local_bb3_reduction_8_i531);

// This section implements an unregistered operation.
// 
wire local_bb3_or102_i398_stall_local;
wire [31:0] local_bb3_or102_i398;

assign local_bb3_or102_i398 = ((local_bb3_conv99_i396 & 32'h1) | (local_bb3_conv101_i397 & 32'h1));

// This section implements a registered operation.
// 
wire SFC_1_VALID_366_367_0_inputs_ready;
 reg SFC_1_VALID_366_367_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_366_367_0_stall_in;
wire SFC_1_VALID_366_367_0_output_regs_ready;
 reg SFC_1_VALID_366_367_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_366_367_0_causedstall;

assign SFC_1_VALID_366_367_0_inputs_ready = 1'b1;
assign SFC_1_VALID_366_367_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_365_366_0_stall_in = 1'b0;
assign SFC_1_VALID_366_367_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_366_367_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_366_367_0_output_regs_ready)
		begin
			SFC_1_VALID_366_367_0_NO_SHIFT_REG <= SFC_1_VALID_365_366_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and17_i511_valid_out_2;
wire local_bb3_and17_i511_stall_in_2;
wire local_bb3_var__u28_valid_out;
wire local_bb3_var__u28_stall_in;
wire local_bb3_add193_i_valid_out;
wire local_bb3_add193_i_stall_in;
wire local_bb3__26_i533_valid_out;
wire local_bb3__26_i533_stall_in;
wire local_bb3__26_i533_inputs_ready;
wire local_bb3__26_i533_stall_local;
wire local_bb3__26_i533;

assign local_bb3__26_i533_inputs_ready = (rnode_333to335_bb3_shr16_i510_0_valid_out_0_NO_SHIFT_REG & rnode_333to335_bb3_cmp27_i519_0_valid_out_2_NO_SHIFT_REG & rnode_334to335_bb3_and37_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_334to335_bb3_xor189_i_0_valid_out_NO_SHIFT_REG & rnode_334to335_bb3_and20_i514_0_valid_out_0_NO_SHIFT_REG & rnode_333to335_bb3_cmp27_i519_0_valid_out_0_NO_SHIFT_REG & rnode_334to335_bb3_lnot33_not_i524_0_valid_out_NO_SHIFT_REG & rnode_333to335_bb3_cmp27_i519_0_valid_out_1_NO_SHIFT_REG & rnode_334to335_bb3_and20_i514_0_valid_out_1_NO_SHIFT_REG & rnode_334to335_bb3_cmp38_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3__26_i533 = (local_bb3_reduction_9_i532 ? rnode_334to335_bb3_cmp38_i_0_NO_SHIFT_REG : local_bb3__24_i528);
assign local_bb3_and17_i511_valid_out_2 = 1'b1;
assign local_bb3_var__u28_valid_out = 1'b1;
assign local_bb3_add193_i_valid_out = 1'b1;
assign local_bb3__26_i533_valid_out = 1'b1;
assign rnode_333to335_bb3_shr16_i510_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_333to335_bb3_cmp27_i519_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_and37_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_xor189_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_and20_i514_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_333to335_bb3_cmp27_i519_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_lnot33_not_i524_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_333to335_bb3_cmp27_i519_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_and20_i514_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_334to335_bb3_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_tobool103_i399_stall_local;
wire local_bb3_tobool103_i399;

assign local_bb3_tobool103_i399 = ((local_bb3_or102_i398 & 32'h1) != 32'h0);

// This section implements a registered operation.
// 
wire SFC_1_VALID_367_368_0_inputs_ready;
 reg SFC_1_VALID_367_368_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_367_368_0_stall_in;
wire SFC_1_VALID_367_368_0_output_regs_ready;
 reg SFC_1_VALID_367_368_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_367_368_0_causedstall;

assign SFC_1_VALID_367_368_0_inputs_ready = 1'b1;
assign SFC_1_VALID_367_368_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_366_367_0_stall_in = 1'b0;
assign SFC_1_VALID_367_368_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_367_368_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_367_368_0_output_regs_ready)
		begin
			SFC_1_VALID_367_368_0_NO_SHIFT_REG <= SFC_1_VALID_366_367_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_335to337_bb3_and17_i511_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and17_i511_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_and17_i511_0_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and17_i511_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to337_bb3_and17_i511_0_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and17_i511_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and17_i511_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_335to337_bb3_and17_i511_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_335to337_bb3_and17_i511_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to337_bb3_and17_i511_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to337_bb3_and17_i511_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_335to337_bb3_and17_i511_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_335to337_bb3_and17_i511_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((local_bb3_and17_i511 & 32'hFF)),
	.data_out(rnode_335to337_bb3_and17_i511_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_335to337_bb3_and17_i511_0_reg_337_fifo.DEPTH = 2;
defparam rnode_335to337_bb3_and17_i511_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_335to337_bb3_and17_i511_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to337_bb3_and17_i511_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_335to337_bb3_and17_i511_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and17_i511_stall_in_2 = 1'b0;
assign rnode_335to337_bb3_and17_i511_0_NO_SHIFT_REG = rnode_335to337_bb3_and17_i511_0_reg_337_NO_SHIFT_REG;
assign rnode_335to337_bb3_and17_i511_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_and17_i511_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_335to336_bb3_var__u28_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u28_0_stall_in_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u28_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u28_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u28_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u28_0_valid_out_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u28_0_stall_in_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_var__u28_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_335to336_bb3_var__u28_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to336_bb3_var__u28_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to336_bb3_var__u28_0_stall_in_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_335to336_bb3_var__u28_0_valid_out_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_335to336_bb3_var__u28_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in(local_bb3_var__u28),
	.data_out(rnode_335to336_bb3_var__u28_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_335to336_bb3_var__u28_0_reg_336_fifo.DEPTH = 1;
defparam rnode_335to336_bb3_var__u28_0_reg_336_fifo.DATA_WIDTH = 1;
defparam rnode_335to336_bb3_var__u28_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to336_bb3_var__u28_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_335to336_bb3_var__u28_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u28_stall_in = 1'b0;
assign rnode_335to336_bb3_var__u28_0_NO_SHIFT_REG = rnode_335to336_bb3_var__u28_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3_var__u28_0_stall_in_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3_var__u28_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_335to336_bb3_add193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3_add193_i_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3_add193_i_1_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3_add193_i_2_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3_add193_i_3_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_335to336_bb3_add193_i_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_valid_out_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_stall_in_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3_add193_i_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_335to336_bb3_add193_i_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to336_bb3_add193_i_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to336_bb3_add193_i_0_stall_in_0_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_335to336_bb3_add193_i_0_valid_out_0_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_335to336_bb3_add193_i_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in(local_bb3_add193_i),
	.data_out(rnode_335to336_bb3_add193_i_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_335to336_bb3_add193_i_0_reg_336_fifo.DEPTH = 1;
defparam rnode_335to336_bb3_add193_i_0_reg_336_fifo.DATA_WIDTH = 32;
defparam rnode_335to336_bb3_add193_i_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to336_bb3_add193_i_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_335to336_bb3_add193_i_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add193_i_stall_in = 1'b0;
assign rnode_335to336_bb3_add193_i_0_stall_in_0_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3_add193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3_add193_i_0_NO_SHIFT_REG = rnode_335to336_bb3_add193_i_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3_add193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3_add193_i_1_NO_SHIFT_REG = rnode_335to336_bb3_add193_i_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3_add193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3_add193_i_2_NO_SHIFT_REG = rnode_335to336_bb3_add193_i_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3_add193_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3_add193_i_3_NO_SHIFT_REG = rnode_335to336_bb3_add193_i_0_reg_336_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_335to336_bb3__26_i533_0_valid_out_NO_SHIFT_REG;
 logic rnode_335to336_bb3__26_i533_0_stall_in_NO_SHIFT_REG;
 logic rnode_335to336_bb3__26_i533_0_NO_SHIFT_REG;
 logic rnode_335to336_bb3__26_i533_0_reg_336_inputs_ready_NO_SHIFT_REG;
 logic rnode_335to336_bb3__26_i533_0_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__26_i533_0_valid_out_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__26_i533_0_stall_in_reg_336_NO_SHIFT_REG;
 logic rnode_335to336_bb3__26_i533_0_stall_out_reg_336_NO_SHIFT_REG;

acl_data_fifo rnode_335to336_bb3__26_i533_0_reg_336_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_335to336_bb3__26_i533_0_reg_336_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_335to336_bb3__26_i533_0_stall_in_reg_336_NO_SHIFT_REG),
	.valid_out(rnode_335to336_bb3__26_i533_0_valid_out_reg_336_NO_SHIFT_REG),
	.stall_out(rnode_335to336_bb3__26_i533_0_stall_out_reg_336_NO_SHIFT_REG),
	.data_in(local_bb3__26_i533),
	.data_out(rnode_335to336_bb3__26_i533_0_reg_336_NO_SHIFT_REG)
);

defparam rnode_335to336_bb3__26_i533_0_reg_336_fifo.DEPTH = 1;
defparam rnode_335to336_bb3__26_i533_0_reg_336_fifo.DATA_WIDTH = 1;
defparam rnode_335to336_bb3__26_i533_0_reg_336_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_335to336_bb3__26_i533_0_reg_336_fifo.IMPL = "shift_reg";

assign rnode_335to336_bb3__26_i533_0_reg_336_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__26_i533_stall_in = 1'b0;
assign rnode_335to336_bb3__26_i533_0_NO_SHIFT_REG = rnode_335to336_bb3__26_i533_0_reg_336_NO_SHIFT_REG;
assign rnode_335to336_bb3__26_i533_0_stall_in_reg_336_NO_SHIFT_REG = 1'b0;
assign rnode_335to336_bb3__26_i533_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cond107_i400_stall_local;
wire [31:0] local_bb3_cond107_i400;

assign local_bb3_cond107_i400 = (local_bb3_tobool103_i399 ? (local_bb3_and4_i317 & 32'h80000000) : 32'hFFFFFFFF);

// This section implements a registered operation.
// 
wire SFC_1_VALID_368_369_0_inputs_ready;
 reg SFC_1_VALID_368_369_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_368_369_0_stall_in;
wire SFC_1_VALID_368_369_0_output_regs_ready;
 reg SFC_1_VALID_368_369_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_368_369_0_causedstall;

assign SFC_1_VALID_368_369_0_inputs_ready = 1'b1;
assign SFC_1_VALID_368_369_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_367_368_0_stall_in = 1'b0;
assign SFC_1_VALID_368_369_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_368_369_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_368_369_0_output_regs_ready)
		begin
			SFC_1_VALID_368_369_0_NO_SHIFT_REG <= SFC_1_VALID_367_368_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_var__u28_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_var__u28_0_stall_in_NO_SHIFT_REG;
 logic rnode_336to337_bb3_var__u28_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_var__u28_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to337_bb3_var__u28_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_var__u28_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_var__u28_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_var__u28_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_var__u28_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_var__u28_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_var__u28_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_var__u28_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_var__u28_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in(rnode_335to336_bb3_var__u28_0_NO_SHIFT_REG),
	.data_out(rnode_336to337_bb3_var__u28_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_var__u28_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_var__u28_0_reg_337_fifo.DATA_WIDTH = 1;
defparam rnode_336to337_bb3_var__u28_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_var__u28_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_var__u28_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3_var__u28_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_var__u28_0_NO_SHIFT_REG = rnode_336to337_bb3_var__u28_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_var__u28_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_var__u28_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and194_i_valid_out;
wire local_bb3_and194_i_stall_in;
wire local_bb3_and194_i_inputs_ready;
wire local_bb3_and194_i_stall_local;
wire [31:0] local_bb3_and194_i;

assign local_bb3_and194_i_inputs_ready = rnode_335to336_bb3_add193_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_and194_i = (rnode_335to336_bb3_add193_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb3_and194_i_valid_out = 1'b1;
assign rnode_335to336_bb3_add193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and196_i_valid_out;
wire local_bb3_and196_i_stall_in;
wire local_bb3_and196_i_inputs_ready;
wire local_bb3_and196_i_stall_local;
wire [31:0] local_bb3_and196_i;

assign local_bb3_and196_i_inputs_ready = rnode_335to336_bb3_add193_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_and196_i = (rnode_335to336_bb3_add193_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb3_and196_i_valid_out = 1'b1;
assign rnode_335to336_bb3_add193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and199_i_valid_out;
wire local_bb3_and199_i_stall_in;
wire local_bb3_and199_i_inputs_ready;
wire local_bb3_and199_i_stall_local;
wire [31:0] local_bb3_and199_i;

assign local_bb3_and199_i_inputs_ready = rnode_335to336_bb3_add193_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_and199_i = (rnode_335to336_bb3_add193_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb3_and199_i_valid_out = 1'b1;
assign rnode_335to336_bb3_add193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and202_i_stall_local;
wire [31:0] local_bb3_and202_i;

assign local_bb3_and202_i = (rnode_335to336_bb3_add193_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_336to338_bb3__26_i533_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to338_bb3__26_i533_0_stall_in_NO_SHIFT_REG;
 logic rnode_336to338_bb3__26_i533_0_NO_SHIFT_REG;
 logic rnode_336to338_bb3__26_i533_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic rnode_336to338_bb3__26_i533_0_reg_338_NO_SHIFT_REG;
 logic rnode_336to338_bb3__26_i533_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_336to338_bb3__26_i533_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_336to338_bb3__26_i533_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_336to338_bb3__26_i533_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to338_bb3__26_i533_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to338_bb3__26_i533_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_336to338_bb3__26_i533_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_336to338_bb3__26_i533_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(rnode_335to336_bb3__26_i533_0_NO_SHIFT_REG),
	.data_out(rnode_336to338_bb3__26_i533_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_336to338_bb3__26_i533_0_reg_338_fifo.DEPTH = 2;
defparam rnode_336to338_bb3__26_i533_0_reg_338_fifo.DATA_WIDTH = 1;
defparam rnode_336to338_bb3__26_i533_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to338_bb3__26_i533_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_336to338_bb3__26_i533_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_335to336_bb3__26_i533_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to338_bb3__26_i533_0_NO_SHIFT_REG = rnode_336to338_bb3__26_i533_0_reg_338_NO_SHIFT_REG;
assign rnode_336to338_bb3__26_i533_0_stall_in_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_336to338_bb3__26_i533_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and108_i401_stall_local;
wire [31:0] local_bb3_and108_i401;

assign local_bb3_and108_i401 = (local_bb3_cond107_i400 & local_bb3_or89_i391);

// This section implements a registered operation.
// 
wire SFC_1_VALID_369_370_0_inputs_ready;
 reg SFC_1_VALID_369_370_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_369_370_0_stall_in;
wire SFC_1_VALID_369_370_0_output_regs_ready;
 reg SFC_1_VALID_369_370_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_369_370_0_causedstall;

assign SFC_1_VALID_369_370_0_inputs_ready = 1'b1;
assign SFC_1_VALID_369_370_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_368_369_0_stall_in = 1'b0;
assign SFC_1_VALID_369_370_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_369_370_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_369_370_0_output_regs_ready)
		begin
			SFC_1_VALID_369_370_0_NO_SHIFT_REG <= SFC_1_VALID_368_369_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_337to338_bb3_var__u28_0_valid_out_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u28_0_stall_in_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u28_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u28_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u28_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u28_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u28_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u28_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_337to338_bb3_var__u28_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to338_bb3_var__u28_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to338_bb3_var__u28_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_337to338_bb3_var__u28_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_337to338_bb3_var__u28_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(rnode_336to337_bb3_var__u28_0_NO_SHIFT_REG),
	.data_out(rnode_337to338_bb3_var__u28_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_337to338_bb3_var__u28_0_reg_338_fifo.DEPTH = 1;
defparam rnode_337to338_bb3_var__u28_0_reg_338_fifo.DATA_WIDTH = 1;
defparam rnode_337to338_bb3_var__u28_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to338_bb3_var__u28_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_337to338_bb3_var__u28_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3_var__u28_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_var__u28_0_NO_SHIFT_REG = rnode_337to338_bb3_var__u28_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3_var__u28_0_stall_in_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_var__u28_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_and194_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and194_i_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and194_i_1_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and194_i_2_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and194_i_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_valid_out_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_stall_in_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and194_i_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_and194_i_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_and194_i_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_and194_i_0_stall_in_0_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_and194_i_0_valid_out_0_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_and194_i_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((local_bb3_and194_i & 32'hFFFFFFF)),
	.data_out(rnode_336to337_bb3_and194_i_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_and194_i_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_and194_i_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_336to337_bb3_and194_i_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_and194_i_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_and194_i_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and194_i_stall_in = 1'b0;
assign rnode_336to337_bb3_and194_i_0_stall_in_0_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and194_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3_and194_i_0_NO_SHIFT_REG = rnode_336to337_bb3_and194_i_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_and194_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3_and194_i_1_NO_SHIFT_REG = rnode_336to337_bb3_and194_i_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_and194_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3_and194_i_2_NO_SHIFT_REG = rnode_336to337_bb3_and194_i_0_reg_337_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_and196_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and196_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and196_i_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and196_i_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and196_i_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and196_i_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and196_i_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and196_i_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_and196_i_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_and196_i_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_and196_i_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_and196_i_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_and196_i_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((local_bb3_and196_i & 32'h1F)),
	.data_out(rnode_336to337_bb3_and196_i_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_and196_i_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_and196_i_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_336to337_bb3_and196_i_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_and196_i_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_and196_i_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and196_i_stall_in = 1'b0;
assign rnode_336to337_bb3_and196_i_0_NO_SHIFT_REG = rnode_336to337_bb3_and196_i_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_and196_i_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and196_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3_and199_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and199_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and199_i_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and199_i_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3_and199_i_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and199_i_0_valid_out_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and199_i_0_stall_in_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3_and199_i_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3_and199_i_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3_and199_i_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3_and199_i_0_stall_in_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3_and199_i_0_valid_out_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3_and199_i_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((local_bb3_and199_i & 32'h1)),
	.data_out(rnode_336to337_bb3_and199_i_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3_and199_i_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3_and199_i_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_336to337_bb3_and199_i_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3_and199_i_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3_and199_i_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and199_i_stall_in = 1'b0;
assign rnode_336to337_bb3_and199_i_0_NO_SHIFT_REG = rnode_336to337_bb3_and199_i_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3_and199_i_0_stall_in_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and199_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i_i559_stall_local;
wire [31:0] local_bb3_shr_i_i559;

assign local_bb3_shr_i_i559 = ((local_bb3_and202_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb3__26_i533_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_2_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_valid_out_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_stall_in_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3__26_i533_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb3__26_i533_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb3__26_i533_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb3__26_i533_0_stall_in_0_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb3__26_i533_0_valid_out_0_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb3__26_i533_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in(rnode_336to338_bb3__26_i533_0_NO_SHIFT_REG),
	.data_out(rnode_338to339_bb3__26_i533_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb3__26_i533_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb3__26_i533_0_reg_339_fifo.DATA_WIDTH = 1;
defparam rnode_338to339_bb3__26_i533_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb3__26_i533_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_338to339_bb3__26_i533_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_336to338_bb3__26_i533_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__26_i533_0_stall_in_0_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__26_i533_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3__26_i533_0_NO_SHIFT_REG = rnode_338to339_bb3__26_i533_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3__26_i533_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3__26_i533_1_NO_SHIFT_REG = rnode_338to339_bb3__26_i533_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3__26_i533_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3__26_i533_2_NO_SHIFT_REG = rnode_338to339_bb3__26_i533_0_reg_339_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or112_i403_stall_local;
wire [31:0] local_bb3_or112_i403;

assign local_bb3_or112_i403 = (local_bb3_and108_i401 | (local_bb3_cond111_i402 & 32'h7F800000));

// This section implements a registered operation.
// 
wire SFC_1_VALID_370_371_0_inputs_ready;
 reg SFC_1_VALID_370_371_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_370_371_0_stall_in;
wire SFC_1_VALID_370_371_0_output_regs_ready;
 reg SFC_1_VALID_370_371_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_370_371_0_causedstall;

assign SFC_1_VALID_370_371_0_inputs_ready = 1'b1;
assign SFC_1_VALID_370_371_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_369_370_0_stall_in = 1'b0;
assign SFC_1_VALID_370_371_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_370_371_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_370_371_0_output_regs_ready)
		begin
			SFC_1_VALID_370_371_0_NO_SHIFT_REG <= SFC_1_VALID_369_370_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_shr217_i_stall_local;
wire [31:0] local_bb3_shr217_i;

assign local_bb3_shr217_i = ((rnode_336to337_bb3_and194_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__pre_i573_stall_local;
wire [31:0] local_bb3__pre_i573;

assign local_bb3__pre_i573 = ((rnode_336to337_bb3_and196_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i_i560_stall_local;
wire [31:0] local_bb3_or_i_i560;

assign local_bb3_or_i_i560 = ((local_bb3_shr_i_i559 & 32'h3FFFFFF) | (local_bb3_and202_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cond293_i_stall_local;
wire [31:0] local_bb3_cond293_i;

assign local_bb3_cond293_i = (rnode_338to339_bb3__26_i533_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u36_stall_local;
wire [31:0] local_bb3_var__u36;

assign local_bb3_var__u36[31:1] = 31'h0;
assign local_bb3_var__u36[0] = rnode_338to339_bb3__26_i533_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u37_valid_out;
wire local_bb3_var__u37_stall_in;
wire local_bb3_var__u37_inputs_ready;
wire local_bb3_var__u37_stall_local;
wire [31:0] local_bb3_var__u37;

assign local_bb3_var__u37_inputs_ready = (rnode_336to337_bb3_xor_i316_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3__29_i345_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3_or581_i374_0_valid_out_1_NO_SHIFT_REG & rnode_336to337_bb3_or581_i374_0_valid_out_0_NO_SHIFT_REG & rnode_336to337_bb3_reduction_0_i375_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3_cmp68_i377_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3_cmp71_not_i394_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3_shl_i381_0_valid_out_NO_SHIFT_REG & rnode_335to337_bb3_and75_i378_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3__40_i387_0_valid_out_NO_SHIFT_REG);
assign local_bb3_var__u37 = (rnode_336to337_bb3__29_i345_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb3_or112_i403);
assign local_bb3_var__u37_valid_out = 1'b1;
assign rnode_336to337_bb3_xor_i316_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__29_i345_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_or581_i374_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_or581_i374_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_reduction_0_i375_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_cmp68_i377_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_cmp71_not_i394_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_shl_i381_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_and75_i378_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__40_i387_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_371_372_0_inputs_ready;
 reg SFC_1_VALID_371_372_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_371_372_0_stall_in;
wire SFC_1_VALID_371_372_0_output_regs_ready;
 reg SFC_1_VALID_371_372_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_371_372_0_causedstall;

assign SFC_1_VALID_371_372_0_inputs_ready = 1'b1;
assign SFC_1_VALID_371_372_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_370_371_0_stall_in = 1'b0;
assign SFC_1_VALID_371_372_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_371_372_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_371_372_0_output_regs_ready)
		begin
			SFC_1_VALID_371_372_0_NO_SHIFT_REG <= SFC_1_VALID_370_371_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_or220_i_stall_local;
wire [31:0] local_bb3_or220_i;

assign local_bb3_or220_i = ((local_bb3_shr217_i & 32'h7FFFFFF) | (rnode_336to337_bb3_and199_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool214_i_stall_local;
wire local_bb3_tobool214_i;

assign local_bb3_tobool214_i = ((local_bb3__pre_i573 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_shr1_i_i561_stall_local;
wire [31:0] local_bb3_shr1_i_i561;

assign local_bb3_shr1_i_i561 = ((local_bb3_or_i_i560 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext_i590_stall_local;
wire [31:0] local_bb3_lnot_ext_i590;

assign local_bb3_lnot_ext_i590 = ((local_bb3_var__u36 & 32'h1) ^ 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_337to338_bb3_var__u37_0_valid_out_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u37_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_var__u37_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u37_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_var__u37_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u37_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u37_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_var__u37_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_337to338_bb3_var__u37_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to338_bb3_var__u37_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to338_bb3_var__u37_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_337to338_bb3_var__u37_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_337to338_bb3_var__u37_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(local_bb3_var__u37),
	.data_out(rnode_337to338_bb3_var__u37_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_337to338_bb3_var__u37_0_reg_338_fifo.DEPTH = 1;
defparam rnode_337to338_bb3_var__u37_0_reg_338_fifo.DATA_WIDTH = 32;
defparam rnode_337to338_bb3_var__u37_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to338_bb3_var__u37_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_337to338_bb3_var__u37_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u37_stall_in = 1'b0;
assign rnode_337to338_bb3_var__u37_0_NO_SHIFT_REG = rnode_337to338_bb3_var__u37_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3_var__u37_0_stall_in_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_var__u37_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_372_373_0_inputs_ready;
 reg SFC_1_VALID_372_373_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_372_373_0_stall_in;
wire SFC_1_VALID_372_373_0_output_regs_ready;
 reg SFC_1_VALID_372_373_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_372_373_0_causedstall;

assign SFC_1_VALID_372_373_0_inputs_ready = 1'b1;
assign SFC_1_VALID_372_373_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_371_372_0_stall_in = 1'b0;
assign SFC_1_VALID_372_373_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_372_373_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_372_373_0_output_regs_ready)
		begin
			SFC_1_VALID_372_373_0_NO_SHIFT_REG <= SFC_1_VALID_371_372_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__40_demorgan_i574_stall_local;
wire local_bb3__40_demorgan_i574;

assign local_bb3__40_demorgan_i574 = (rnode_335to337_bb3_cmp38_i_0_NO_SHIFT_REG | local_bb3_tobool214_i);

// This section implements an unregistered operation.
// 
wire local_bb3__42_i575_stall_local;
wire local_bb3__42_i575;

assign local_bb3__42_i575 = (local_bb3_tobool214_i & local_bb3_not_cmp38_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or2_i_i562_stall_local;
wire [31:0] local_bb3_or2_i_i562;

assign local_bb3_or2_i_i562 = ((local_bb3_shr1_i_i561 & 32'h1FFFFFF) | (local_bb3_or_i_i560 & 32'h7FFFFFF));

// Register node:
//  * latency = 36
//  * capacity = 36
 logic rnode_338to374_bb3_var__u37_0_valid_out_NO_SHIFT_REG;
 logic rnode_338to374_bb3_var__u37_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_338to374_bb3_var__u37_0_NO_SHIFT_REG;
 logic rnode_338to374_bb3_var__u37_0_reg_374_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_338to374_bb3_var__u37_0_reg_374_NO_SHIFT_REG;
 logic rnode_338to374_bb3_var__u37_0_valid_out_reg_374_NO_SHIFT_REG;
 logic rnode_338to374_bb3_var__u37_0_stall_in_reg_374_NO_SHIFT_REG;
 logic rnode_338to374_bb3_var__u37_0_stall_out_reg_374_NO_SHIFT_REG;

acl_data_fifo rnode_338to374_bb3_var__u37_0_reg_374_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to374_bb3_var__u37_0_reg_374_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to374_bb3_var__u37_0_stall_in_reg_374_NO_SHIFT_REG),
	.valid_out(rnode_338to374_bb3_var__u37_0_valid_out_reg_374_NO_SHIFT_REG),
	.stall_out(rnode_338to374_bb3_var__u37_0_stall_out_reg_374_NO_SHIFT_REG),
	.data_in(rnode_337to338_bb3_var__u37_0_NO_SHIFT_REG),
	.data_out(rnode_338to374_bb3_var__u37_0_reg_374_NO_SHIFT_REG)
);

defparam rnode_338to374_bb3_var__u37_0_reg_374_fifo.DEPTH = 36;
defparam rnode_338to374_bb3_var__u37_0_reg_374_fifo.DATA_WIDTH = 32;
defparam rnode_338to374_bb3_var__u37_0_reg_374_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to374_bb3_var__u37_0_reg_374_fifo.IMPL = "shift_reg";

assign rnode_338to374_bb3_var__u37_0_reg_374_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_337to338_bb3_var__u37_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_338to374_bb3_var__u37_0_NO_SHIFT_REG = rnode_338to374_bb3_var__u37_0_reg_374_NO_SHIFT_REG;
assign rnode_338to374_bb3_var__u37_0_stall_in_reg_374_NO_SHIFT_REG = 1'b0;
assign rnode_338to374_bb3_var__u37_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_373_374_0_inputs_ready;
 reg SFC_1_VALID_373_374_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_373_374_0_stall_in;
wire SFC_1_VALID_373_374_0_output_regs_ready;
 reg SFC_1_VALID_373_374_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_373_374_0_causedstall;

assign SFC_1_VALID_373_374_0_inputs_ready = 1'b1;
assign SFC_1_VALID_373_374_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_372_373_0_stall_in = 1'b0;
assign SFC_1_VALID_373_374_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_373_374_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_373_374_0_output_regs_ready)
		begin
			SFC_1_VALID_373_374_0_NO_SHIFT_REG <= SFC_1_VALID_372_373_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__43_i576_stall_local;
wire [31:0] local_bb3__43_i576;

assign local_bb3__43_i576 = (local_bb3__42_i575 ? 32'h0 : (local_bb3__pre_i573 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_shr3_i_i563_stall_local;
wire [31:0] local_bb3_shr3_i_i563;

assign local_bb3_shr3_i_i563 = ((local_bb3_or2_i_i562 & 32'h7FFFFFF) >> 32'h4);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_374to375_bb3_var__u37_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_374to375_bb3_var__u37_0_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_374to375_bb3_var__u37_1_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_374to375_bb3_var__u37_2_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_reg_375_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_374to375_bb3_var__u37_0_reg_375_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_valid_out_0_reg_375_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_stall_in_0_reg_375_NO_SHIFT_REG;
 logic rnode_374to375_bb3_var__u37_0_stall_out_reg_375_NO_SHIFT_REG;

acl_data_fifo rnode_374to375_bb3_var__u37_0_reg_375_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_374to375_bb3_var__u37_0_reg_375_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_374to375_bb3_var__u37_0_stall_in_0_reg_375_NO_SHIFT_REG),
	.valid_out(rnode_374to375_bb3_var__u37_0_valid_out_0_reg_375_NO_SHIFT_REG),
	.stall_out(rnode_374to375_bb3_var__u37_0_stall_out_reg_375_NO_SHIFT_REG),
	.data_in(rnode_338to374_bb3_var__u37_0_NO_SHIFT_REG),
	.data_out(rnode_374to375_bb3_var__u37_0_reg_375_NO_SHIFT_REG)
);

defparam rnode_374to375_bb3_var__u37_0_reg_375_fifo.DEPTH = 1;
defparam rnode_374to375_bb3_var__u37_0_reg_375_fifo.DATA_WIDTH = 32;
defparam rnode_374to375_bb3_var__u37_0_reg_375_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_374to375_bb3_var__u37_0_reg_375_fifo.IMPL = "shift_reg";

assign rnode_374to375_bb3_var__u37_0_reg_375_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_338to374_bb3_var__u37_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_374to375_bb3_var__u37_0_stall_in_0_reg_375_NO_SHIFT_REG = 1'b0;
assign rnode_374to375_bb3_var__u37_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_374to375_bb3_var__u37_0_NO_SHIFT_REG = rnode_374to375_bb3_var__u37_0_reg_375_NO_SHIFT_REG;
assign rnode_374to375_bb3_var__u37_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_374to375_bb3_var__u37_1_NO_SHIFT_REG = rnode_374to375_bb3_var__u37_0_reg_375_NO_SHIFT_REG;
assign rnode_374to375_bb3_var__u37_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_374to375_bb3_var__u37_2_NO_SHIFT_REG = rnode_374to375_bb3_var__u37_0_reg_375_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_1_VALID_374_375_0_inputs_ready;
 reg SFC_1_VALID_374_375_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_374_375_0_stall_in;
wire SFC_1_VALID_374_375_0_output_regs_ready;
 reg SFC_1_VALID_374_375_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_374_375_0_causedstall;

assign SFC_1_VALID_374_375_0_inputs_ready = 1'b1;
assign SFC_1_VALID_374_375_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_373_374_0_stall_in = 1'b0;
assign SFC_1_VALID_374_375_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_374_375_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_374_375_0_output_regs_ready)
		begin
			SFC_1_VALID_374_375_0_NO_SHIFT_REG <= SFC_1_VALID_373_374_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_or4_i_i564_stall_local;
wire [31:0] local_bb3_or4_i_i564;

assign local_bb3_or4_i_i564 = ((local_bb3_shr3_i_i563 & 32'h7FFFFF) | (local_bb3_or2_i_i562 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i220_stall_local;
wire [31:0] local_bb3_shr_i220;

assign local_bb3_shr_i220 = (rnode_374to375_bb3_var__u37_0_NO_SHIFT_REG >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and5_i226_stall_local;
wire [31:0] local_bb3_and5_i226;

assign local_bb3_and5_i226 = (rnode_374to375_bb3_var__u37_2_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements a registered operation.
// 
wire SFC_1_VALID_375_376_0_inputs_ready;
 reg SFC_1_VALID_375_376_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_375_376_0_stall_in;
wire SFC_1_VALID_375_376_0_output_regs_ready;
 reg SFC_1_VALID_375_376_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_375_376_0_causedstall;

assign SFC_1_VALID_375_376_0_inputs_ready = 1'b1;
assign SFC_1_VALID_375_376_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_374_375_0_stall_in = 1'b0;
assign SFC_1_VALID_375_376_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_375_376_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_375_376_0_output_regs_ready)
		begin
			SFC_1_VALID_375_376_0_NO_SHIFT_REG <= SFC_1_VALID_374_375_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_shr5_i_i565_stall_local;
wire [31:0] local_bb3_shr5_i_i565;

assign local_bb3_shr5_i_i565 = ((local_bb3_or4_i_i564 & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_and_i221_stall_local;
wire [31:0] local_bb3_and_i221;

assign local_bb3_and_i221 = ((local_bb3_shr_i220 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_i232_stall_local;
wire local_bb3_lnot14_i232;

assign local_bb3_lnot14_i232 = ((local_bb3_and5_i226 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i254_stall_local;
wire [31:0] local_bb3_or_i254;

assign local_bb3_or_i254 = ((local_bb3_and5_i226 & 32'h7FFFFF) | 32'h800000);

// This section implements a registered operation.
// 
wire SFC_1_VALID_376_377_0_inputs_ready;
 reg SFC_1_VALID_376_377_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_376_377_0_stall_in;
wire SFC_1_VALID_376_377_0_output_regs_ready;
 reg SFC_1_VALID_376_377_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_376_377_0_causedstall;

assign SFC_1_VALID_376_377_0_inputs_ready = 1'b1;
assign SFC_1_VALID_376_377_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_375_376_0_stall_in = 1'b0;
assign SFC_1_VALID_376_377_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_376_377_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_376_377_0_output_regs_ready)
		begin
			SFC_1_VALID_376_377_0_NO_SHIFT_REG <= SFC_1_VALID_375_376_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_or6_i_i566_stall_local;
wire [31:0] local_bb3_or6_i_i566;

assign local_bb3_or6_i_i566 = ((local_bb3_shr5_i_i565 & 32'h7FFFF) | (local_bb3_or4_i_i564 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_i228_stall_local;
wire local_bb3_lnot_i228;

assign local_bb3_lnot_i228 = ((local_bb3_and_i221 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i230_stall_local;
wire local_bb3_cmp_i230;

assign local_bb3_cmp_i230 = ((local_bb3_and_i221 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_conv_i_i256_stall_local;
wire [63:0] local_bb3_conv_i_i256;

assign local_bb3_conv_i_i256[63:32] = 32'h0;
assign local_bb3_conv_i_i256[31:0] = ((local_bb3_or_i254 & 32'hFFFFFF) | 32'h800000);

// This section implements a registered operation.
// 
wire SFC_1_VALID_377_378_0_inputs_ready;
 reg SFC_1_VALID_377_378_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_377_378_0_stall_in;
wire SFC_1_VALID_377_378_0_output_regs_ready;
 reg SFC_1_VALID_377_378_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_377_378_0_causedstall;

assign SFC_1_VALID_377_378_0_inputs_ready = 1'b1;
assign SFC_1_VALID_377_378_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_376_377_0_stall_in = 1'b0;
assign SFC_1_VALID_377_378_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_377_378_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_377_378_0_output_regs_ready)
		begin
			SFC_1_VALID_377_378_0_NO_SHIFT_REG <= SFC_1_VALID_376_377_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_shr7_i_i567_stall_local;
wire [31:0] local_bb3_shr7_i_i567;

assign local_bb3_shr7_i_i567 = ((local_bb3_or6_i_i566 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_or6_masked_i_i568_stall_local;
wire [31:0] local_bb3_or6_masked_i_i568;

assign local_bb3_or6_masked_i_i568 = ((local_bb3_or6_i_i566 & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_1_VALID_378_379_0_inputs_ready;
 reg SFC_1_VALID_378_379_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_378_379_0_stall_in;
wire SFC_1_VALID_378_379_0_output_regs_ready;
 reg SFC_1_VALID_378_379_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_378_379_0_causedstall;

assign SFC_1_VALID_378_379_0_inputs_ready = 1'b1;
assign SFC_1_VALID_378_379_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_377_378_0_stall_in = 1'b0;
assign SFC_1_VALID_378_379_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_378_379_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_378_379_0_output_regs_ready)
		begin
			SFC_1_VALID_378_379_0_NO_SHIFT_REG <= SFC_1_VALID_377_378_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_neg_i_i569_stall_local;
wire [31:0] local_bb3_neg_i_i569;

assign local_bb3_neg_i_i569 = ((local_bb3_or6_masked_i_i568 & 32'h7FFFFFF) | (local_bb3_shr7_i_i567 & 32'h7FF));

// This section implements a registered operation.
// 
wire SFC_1_VALID_379_380_0_inputs_ready;
 reg SFC_1_VALID_379_380_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_379_380_0_stall_in;
wire SFC_1_VALID_379_380_0_output_regs_ready;
 reg SFC_1_VALID_379_380_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_379_380_0_causedstall;

assign SFC_1_VALID_379_380_0_inputs_ready = 1'b1;
assign SFC_1_VALID_379_380_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_378_379_0_stall_in = 1'b0;
assign SFC_1_VALID_379_380_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_379_380_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_379_380_0_output_regs_ready)
		begin
			SFC_1_VALID_379_380_0_NO_SHIFT_REG <= SFC_1_VALID_378_379_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and_i_i570_stall_local;
wire [31:0] local_bb3_and_i_i570;

assign local_bb3_and_i_i570 = ((local_bb3_neg_i_i569 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_1_VALID_380_381_0_inputs_ready;
 reg SFC_1_VALID_380_381_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_380_381_0_stall_in;
wire SFC_1_VALID_380_381_0_output_regs_ready;
 reg SFC_1_VALID_380_381_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_380_381_0_causedstall;

assign SFC_1_VALID_380_381_0_inputs_ready = 1'b1;
assign SFC_1_VALID_380_381_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_379_380_0_stall_in = 1'b0;
assign SFC_1_VALID_380_381_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_380_381_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_380_381_0_output_regs_ready)
		begin
			SFC_1_VALID_380_381_0_NO_SHIFT_REG <= SFC_1_VALID_379_380_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__and_i_i570_valid_out;
wire local_bb3__and_i_i570_stall_in;
wire local_bb3__and_i_i570_inputs_ready;
wire local_bb3__and_i_i570_stall_local;
wire [31:0] local_bb3__and_i_i570;

thirtysix_six_comp local_bb3__and_i_i570_popcnt_instance (
	.data((local_bb3_and_i_i570 & 32'h7FFFFFF)),
	.sum(local_bb3__and_i_i570)
);


assign local_bb3__and_i_i570_inputs_ready = rnode_335to336_bb3_add193_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb3__and_i_i570_valid_out = 1'b1;
assign rnode_335to336_bb3_add193_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_381_382_0_inputs_ready;
 reg SFC_1_VALID_381_382_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_381_382_0_stall_in;
wire SFC_1_VALID_381_382_0_output_regs_ready;
 reg SFC_1_VALID_381_382_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_381_382_0_causedstall;

assign SFC_1_VALID_381_382_0_inputs_ready = 1'b1;
assign SFC_1_VALID_381_382_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_380_381_0_stall_in = 1'b0;
assign SFC_1_VALID_381_382_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_381_382_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_381_382_0_output_regs_ready)
		begin
			SFC_1_VALID_381_382_0_NO_SHIFT_REG <= SFC_1_VALID_380_381_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_336to337_bb3__and_i_i570_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3__and_i_i570_0_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3__and_i_i570_1_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3__and_i_i570_2_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_reg_337_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_336to337_bb3__and_i_i570_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_valid_out_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_stall_in_0_reg_337_NO_SHIFT_REG;
 logic rnode_336to337_bb3__and_i_i570_0_stall_out_reg_337_NO_SHIFT_REG;

acl_data_fifo rnode_336to337_bb3__and_i_i570_0_reg_337_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_336to337_bb3__and_i_i570_0_reg_337_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_336to337_bb3__and_i_i570_0_stall_in_0_reg_337_NO_SHIFT_REG),
	.valid_out(rnode_336to337_bb3__and_i_i570_0_valid_out_0_reg_337_NO_SHIFT_REG),
	.stall_out(rnode_336to337_bb3__and_i_i570_0_stall_out_reg_337_NO_SHIFT_REG),
	.data_in((local_bb3__and_i_i570 & 32'h3F)),
	.data_out(rnode_336to337_bb3__and_i_i570_0_reg_337_NO_SHIFT_REG)
);

defparam rnode_336to337_bb3__and_i_i570_0_reg_337_fifo.DEPTH = 1;
defparam rnode_336to337_bb3__and_i_i570_0_reg_337_fifo.DATA_WIDTH = 32;
defparam rnode_336to337_bb3__and_i_i570_0_reg_337_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_336to337_bb3__and_i_i570_0_reg_337_fifo.IMPL = "shift_reg";

assign rnode_336to337_bb3__and_i_i570_0_reg_337_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__and_i_i570_stall_in = 1'b0;
assign rnode_336to337_bb3__and_i_i570_0_stall_in_0_reg_337_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__and_i_i570_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3__and_i_i570_0_NO_SHIFT_REG = rnode_336to337_bb3__and_i_i570_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3__and_i_i570_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3__and_i_i570_1_NO_SHIFT_REG = rnode_336to337_bb3__and_i_i570_0_reg_337_NO_SHIFT_REG;
assign rnode_336to337_bb3__and_i_i570_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_336to337_bb3__and_i_i570_2_NO_SHIFT_REG = rnode_336to337_bb3__and_i_i570_0_reg_337_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_1_VALID_382_383_0_inputs_ready;
 reg SFC_1_VALID_382_383_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_382_383_0_stall_in;
wire SFC_1_VALID_382_383_0_output_regs_ready;
 reg SFC_1_VALID_382_383_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_382_383_0_causedstall;

assign SFC_1_VALID_382_383_0_inputs_ready = 1'b1;
assign SFC_1_VALID_382_383_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_381_382_0_stall_in = 1'b0;
assign SFC_1_VALID_382_383_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_382_383_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_382_383_0_output_regs_ready)
		begin
			SFC_1_VALID_382_383_0_NO_SHIFT_REG <= SFC_1_VALID_381_382_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and9_i_i571_stall_local;
wire [31:0] local_bb3_and9_i_i571;

assign local_bb3_and9_i_i571 = ((rnode_336to337_bb3__and_i_i570_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_and204_i_stall_local;
wire [31:0] local_bb3_and204_i;

assign local_bb3_and204_i = ((rnode_336to337_bb3__and_i_i570_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_and207_i_stall_local;
wire [31:0] local_bb3_and207_i;

assign local_bb3_and207_i = ((rnode_336to337_bb3__and_i_i570_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements a registered operation.
// 
wire SFC_1_VALID_383_384_0_inputs_ready;
 reg SFC_1_VALID_383_384_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_383_384_0_stall_in;
wire SFC_1_VALID_383_384_0_output_regs_ready;
 reg SFC_1_VALID_383_384_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_383_384_0_causedstall;

assign SFC_1_VALID_383_384_0_inputs_ready = 1'b1;
assign SFC_1_VALID_383_384_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_382_383_0_stall_in = 1'b0;
assign SFC_1_VALID_383_384_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_383_384_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_383_384_0_output_regs_ready)
		begin
			SFC_1_VALID_383_384_0_NO_SHIFT_REG <= SFC_1_VALID_382_383_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_sub240_i_stall_local;
wire [31:0] local_bb3_sub240_i;

assign local_bb3_sub240_i = (32'h0 - (local_bb3_and9_i_i571 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb3_shl205_i_stall_local;
wire [31:0] local_bb3_shl205_i;

assign local_bb3_shl205_i = ((rnode_336to337_bb3_and194_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb3_and204_i & 32'h18));

// This section implements a registered operation.
// 
wire SFC_1_VALID_384_385_0_inputs_ready;
 reg SFC_1_VALID_384_385_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_384_385_0_stall_in;
wire SFC_1_VALID_384_385_0_output_regs_ready;
 reg SFC_1_VALID_384_385_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_384_385_0_causedstall;

assign SFC_1_VALID_384_385_0_inputs_ready = 1'b1;
assign SFC_1_VALID_384_385_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_383_384_0_stall_in = 1'b0;
assign SFC_1_VALID_384_385_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_384_385_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_384_385_0_output_regs_ready)
		begin
			SFC_1_VALID_384_385_0_NO_SHIFT_REG <= SFC_1_VALID_383_384_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_cond245_i_stall_local;
wire [31:0] local_bb3_cond245_i;

assign local_bb3_cond245_i = (rnode_335to337_bb3_cmp38_i_2_NO_SHIFT_REG ? local_bb3_sub240_i : (local_bb3__43_i576 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and206_i572_stall_local;
wire [31:0] local_bb3_and206_i572;

assign local_bb3_and206_i572 = (local_bb3_shl205_i & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_1_VALID_385_386_0_inputs_ready;
 reg SFC_1_VALID_385_386_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_385_386_0_stall_in;
wire SFC_1_VALID_385_386_0_output_regs_ready;
 reg SFC_1_VALID_385_386_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_385_386_0_causedstall;

assign SFC_1_VALID_385_386_0_inputs_ready = 1'b1;
assign SFC_1_VALID_385_386_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_384_385_0_stall_in = 1'b0;
assign SFC_1_VALID_385_386_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_385_386_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_385_386_0_output_regs_ready)
		begin
			SFC_1_VALID_385_386_0_NO_SHIFT_REG <= SFC_1_VALID_384_385_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_add246_i_stall_local;
wire [31:0] local_bb3_add246_i;

assign local_bb3_add246_i = (local_bb3_cond245_i + (rnode_335to337_bb3_and17_i511_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_fold_i581_stall_local;
wire [31:0] local_bb3_fold_i581;

assign local_bb3_fold_i581 = (local_bb3_cond245_i + (rnode_335to337_bb3_shr16_i510_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb3_shl208_i_stall_local;
wire [31:0] local_bb3_shl208_i;

assign local_bb3_shl208_i = ((local_bb3_and206_i572 & 32'h7FFFFFF) << (local_bb3_and207_i & 32'h7));

// This section implements a registered operation.
// 
wire SFC_1_VALID_386_387_0_inputs_ready;
 reg SFC_1_VALID_386_387_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_386_387_0_stall_in;
wire SFC_1_VALID_386_387_0_output_regs_ready;
 reg SFC_1_VALID_386_387_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_386_387_0_causedstall;

assign SFC_1_VALID_386_387_0_inputs_ready = 1'b1;
assign SFC_1_VALID_386_387_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_385_386_0_stall_in = 1'b0;
assign SFC_1_VALID_386_387_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_386_387_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_386_387_0_output_regs_ready)
		begin
			SFC_1_VALID_386_387_0_NO_SHIFT_REG <= SFC_1_VALID_385_386_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and251_i_stall_local;
wire [31:0] local_bb3_and251_i;

assign local_bb3_and251_i = (local_bb3_fold_i581 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and270_i586_stall_local;
wire [31:0] local_bb3_and270_i586;

assign local_bb3_and270_i586 = (local_bb3_fold_i581 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and209_i_stall_local;
wire [31:0] local_bb3_and209_i;

assign local_bb3_and209_i = (local_bb3_shl208_i & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_1_VALID_387_388_0_inputs_ready;
 reg SFC_1_VALID_387_388_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_387_388_0_stall_in;
wire SFC_1_VALID_387_388_0_output_regs_ready;
 reg SFC_1_VALID_387_388_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_387_388_0_causedstall;

assign SFC_1_VALID_387_388_0_inputs_ready = 1'b1;
assign SFC_1_VALID_387_388_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_386_387_0_stall_in = 1'b0;
assign SFC_1_VALID_387_388_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_387_388_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_387_388_0_output_regs_ready)
		begin
			SFC_1_VALID_387_388_0_NO_SHIFT_REG <= SFC_1_VALID_386_387_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__44_i577_stall_local;
wire [31:0] local_bb3__44_i577;

assign local_bb3__44_i577 = (local_bb3__40_demorgan_i574 ? (local_bb3_and209_i & 32'h7FFFFFF) : (local_bb3_or220_i & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_1_VALID_388_389_0_inputs_ready;
 reg SFC_1_VALID_388_389_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_388_389_0_stall_in;
wire SFC_1_VALID_388_389_0_output_regs_ready;
 reg SFC_1_VALID_388_389_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_388_389_0_causedstall;

assign SFC_1_VALID_388_389_0_inputs_ready = 1'b1;
assign SFC_1_VALID_388_389_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_387_388_0_stall_in = 1'b0;
assign SFC_1_VALID_388_389_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_388_389_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_388_389_0_output_regs_ready)
		begin
			SFC_1_VALID_388_389_0_NO_SHIFT_REG <= SFC_1_VALID_387_388_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and251_i_valid_out;
wire local_bb3_and251_i_stall_in;
wire local_bb3_and270_i586_valid_out;
wire local_bb3_and270_i586_stall_in;
wire local_bb3_add246_i_valid_out;
wire local_bb3_add246_i_stall_in;
wire local_bb3__45_i578_valid_out;
wire local_bb3__45_i578_stall_in;
wire local_bb3_not_cmp38_i_valid_out_1;
wire local_bb3_not_cmp38_i_stall_in_1;
wire local_bb3__45_i578_inputs_ready;
wire local_bb3__45_i578_stall_local;
wire [31:0] local_bb3__45_i578;

assign local_bb3__45_i578_inputs_ready = (rnode_335to337_bb3_shr16_i510_0_valid_out_NO_SHIFT_REG & rnode_335to337_bb3_and17_i511_0_valid_out_NO_SHIFT_REG & rnode_335to337_bb3_cmp38_i_0_valid_out_2_NO_SHIFT_REG & rnode_335to337_bb3_cmp38_i_0_valid_out_0_NO_SHIFT_REG & rnode_336to337_bb3_and194_i_0_valid_out_2_NO_SHIFT_REG & rnode_335to337_bb3_cmp38_i_0_valid_out_1_NO_SHIFT_REG & rnode_336to337_bb3_and196_i_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3_and194_i_0_valid_out_1_NO_SHIFT_REG & rnode_336to337_bb3_and199_i_0_valid_out_NO_SHIFT_REG & rnode_336to337_bb3_and194_i_0_valid_out_0_NO_SHIFT_REG & rnode_336to337_bb3__and_i_i570_0_valid_out_1_NO_SHIFT_REG & rnode_336to337_bb3__and_i_i570_0_valid_out_2_NO_SHIFT_REG & rnode_336to337_bb3__and_i_i570_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3__45_i578 = (local_bb3__42_i575 ? (rnode_336to337_bb3_and194_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb3__44_i577 & 32'h7FFFFFF));
assign local_bb3_and251_i_valid_out = 1'b1;
assign local_bb3_and270_i586_valid_out = 1'b1;
assign local_bb3_add246_i_valid_out = 1'b1;
assign local_bb3__45_i578_valid_out = 1'b1;
assign local_bb3_not_cmp38_i_valid_out_1 = 1'b1;
assign rnode_335to337_bb3_shr16_i510_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_and17_i511_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_cmp38_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and194_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_335to337_bb3_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and196_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and194_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and199_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3_and194_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__and_i_i570_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__and_i_i570_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_336to337_bb3__and_i_i570_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_389_390_0_inputs_ready;
 reg SFC_1_VALID_389_390_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_389_390_0_stall_in;
wire SFC_1_VALID_389_390_0_output_regs_ready;
 reg SFC_1_VALID_389_390_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_389_390_0_causedstall;

assign SFC_1_VALID_389_390_0_inputs_ready = 1'b1;
assign SFC_1_VALID_389_390_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_388_389_0_stall_in = 1'b0;
assign SFC_1_VALID_389_390_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_389_390_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_389_390_0_output_regs_ready)
		begin
			SFC_1_VALID_389_390_0_NO_SHIFT_REG <= SFC_1_VALID_388_389_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_337to338_bb3_and251_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and251_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_and251_i_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and251_i_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_and251_i_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and251_i_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and251_i_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_and251_i_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_337to338_bb3_and251_i_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to338_bb3_and251_i_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to338_bb3_and251_i_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_337to338_bb3_and251_i_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_337to338_bb3_and251_i_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in((local_bb3_and251_i & 32'hFF)),
	.data_out(rnode_337to338_bb3_and251_i_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_337to338_bb3_and251_i_0_reg_338_fifo.DEPTH = 1;
defparam rnode_337to338_bb3_and251_i_0_reg_338_fifo.DATA_WIDTH = 32;
defparam rnode_337to338_bb3_and251_i_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to338_bb3_and251_i_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_337to338_bb3_and251_i_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and251_i_stall_in = 1'b0;
assign rnode_337to338_bb3_and251_i_0_NO_SHIFT_REG = rnode_337to338_bb3_and251_i_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3_and251_i_0_stall_in_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_and251_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_337to339_bb3_and270_i586_0_valid_out_NO_SHIFT_REG;
 logic rnode_337to339_bb3_and270_i586_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_337to339_bb3_and270_i586_0_NO_SHIFT_REG;
 logic rnode_337to339_bb3_and270_i586_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_337to339_bb3_and270_i586_0_reg_339_NO_SHIFT_REG;
 logic rnode_337to339_bb3_and270_i586_0_valid_out_reg_339_NO_SHIFT_REG;
 logic rnode_337to339_bb3_and270_i586_0_stall_in_reg_339_NO_SHIFT_REG;
 logic rnode_337to339_bb3_and270_i586_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_337to339_bb3_and270_i586_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to339_bb3_and270_i586_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to339_bb3_and270_i586_0_stall_in_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_337to339_bb3_and270_i586_0_valid_out_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_337to339_bb3_and270_i586_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in((local_bb3_and270_i586 & 32'hFF800000)),
	.data_out(rnode_337to339_bb3_and270_i586_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_337to339_bb3_and270_i586_0_reg_339_fifo.DEPTH = 2;
defparam rnode_337to339_bb3_and270_i586_0_reg_339_fifo.DATA_WIDTH = 32;
defparam rnode_337to339_bb3_and270_i586_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to339_bb3_and270_i586_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_337to339_bb3_and270_i586_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and270_i586_stall_in = 1'b0;
assign rnode_337to339_bb3_and270_i586_0_NO_SHIFT_REG = rnode_337to339_bb3_and270_i586_0_reg_339_NO_SHIFT_REG;
assign rnode_337to339_bb3_and270_i586_0_stall_in_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_337to339_bb3_and270_i586_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_337to338_bb3_add246_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3_add246_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_add246_i_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3_add246_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_337to338_bb3_add246_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_add246_i_1_NO_SHIFT_REG;
 logic rnode_337to338_bb3_add246_i_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3_add246_i_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_add246_i_0_valid_out_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_add246_i_0_stall_in_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_add246_i_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_337to338_bb3_add246_i_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to338_bb3_add246_i_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to338_bb3_add246_i_0_stall_in_0_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_337to338_bb3_add246_i_0_valid_out_0_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_337to338_bb3_add246_i_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(local_bb3_add246_i),
	.data_out(rnode_337to338_bb3_add246_i_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_337to338_bb3_add246_i_0_reg_338_fifo.DEPTH = 1;
defparam rnode_337to338_bb3_add246_i_0_reg_338_fifo.DATA_WIDTH = 32;
defparam rnode_337to338_bb3_add246_i_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to338_bb3_add246_i_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_337to338_bb3_add246_i_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add246_i_stall_in = 1'b0;
assign rnode_337to338_bb3_add246_i_0_stall_in_0_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_add246_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_337to338_bb3_add246_i_0_NO_SHIFT_REG = rnode_337to338_bb3_add246_i_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3_add246_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_337to338_bb3_add246_i_1_NO_SHIFT_REG = rnode_337to338_bb3_add246_i_0_reg_338_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_337to338_bb3__45_i578_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3__45_i578_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3__45_i578_1_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3__45_i578_2_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_337to338_bb3__45_i578_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_valid_out_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_stall_in_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3__45_i578_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_337to338_bb3__45_i578_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to338_bb3__45_i578_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to338_bb3__45_i578_0_stall_in_0_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_337to338_bb3__45_i578_0_valid_out_0_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_337to338_bb3__45_i578_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in((local_bb3__45_i578 & 32'hFFFFFFF)),
	.data_out(rnode_337to338_bb3__45_i578_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_337to338_bb3__45_i578_0_reg_338_fifo.DEPTH = 1;
defparam rnode_337to338_bb3__45_i578_0_reg_338_fifo.DATA_WIDTH = 32;
defparam rnode_337to338_bb3__45_i578_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to338_bb3__45_i578_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_337to338_bb3__45_i578_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__45_i578_stall_in = 1'b0;
assign rnode_337to338_bb3__45_i578_0_stall_in_0_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3__45_i578_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_337to338_bb3__45_i578_0_NO_SHIFT_REG = rnode_337to338_bb3__45_i578_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3__45_i578_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_337to338_bb3__45_i578_1_NO_SHIFT_REG = rnode_337to338_bb3__45_i578_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3__45_i578_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_337to338_bb3__45_i578_2_NO_SHIFT_REG = rnode_337to338_bb3__45_i578_0_reg_338_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_337to338_bb3_not_cmp38_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_337to338_bb3_not_cmp38_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_337to338_bb3_not_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_337to338_bb3_not_cmp38_i_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic rnode_337to338_bb3_not_cmp38_i_0_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_not_cmp38_i_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_not_cmp38_i_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_337to338_bb3_not_cmp38_i_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_337to338_bb3_not_cmp38_i_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_337to338_bb3_not_cmp38_i_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_337to338_bb3_not_cmp38_i_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_337to338_bb3_not_cmp38_i_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_337to338_bb3_not_cmp38_i_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(local_bb3_not_cmp38_i),
	.data_out(rnode_337to338_bb3_not_cmp38_i_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_337to338_bb3_not_cmp38_i_0_reg_338_fifo.DEPTH = 1;
defparam rnode_337to338_bb3_not_cmp38_i_0_reg_338_fifo.DATA_WIDTH = 1;
defparam rnode_337to338_bb3_not_cmp38_i_0_reg_338_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_337to338_bb3_not_cmp38_i_0_reg_338_fifo.IMPL = "shift_reg";

assign rnode_337to338_bb3_not_cmp38_i_0_reg_338_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_not_cmp38_i_stall_in_1 = 1'b0;
assign rnode_337to338_bb3_not_cmp38_i_0_NO_SHIFT_REG = rnode_337to338_bb3_not_cmp38_i_0_reg_338_NO_SHIFT_REG;
assign rnode_337to338_bb3_not_cmp38_i_0_stall_in_reg_338_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_not_cmp38_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_390_391_0_inputs_ready;
 reg SFC_1_VALID_390_391_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_390_391_0_stall_in;
wire SFC_1_VALID_390_391_0_output_regs_ready;
 reg SFC_1_VALID_390_391_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_390_391_0_causedstall;

assign SFC_1_VALID_390_391_0_inputs_ready = 1'b1;
assign SFC_1_VALID_390_391_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_389_390_0_stall_in = 1'b0;
assign SFC_1_VALID_390_391_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_390_391_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_390_391_0_output_regs_ready)
		begin
			SFC_1_VALID_390_391_0_NO_SHIFT_REG <= SFC_1_VALID_389_390_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_notrhs_i583_stall_local;
wire local_bb3_notrhs_i583;

assign local_bb3_notrhs_i583 = ((rnode_337to338_bb3_and251_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_shl274_i_stall_local;
wire [31:0] local_bb3_shl274_i;

assign local_bb3_shl274_i = ((rnode_337to339_bb3_and270_i586_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb3_and248_i_stall_local;
wire [31:0] local_bb3_and248_i;

assign local_bb3_and248_i = (rnode_337to338_bb3_add246_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp259_i_stall_local;
wire local_bb3_cmp259_i;

assign local_bb3_cmp259_i = ($signed(rnode_337to338_bb3_add246_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb3_and226_i_stall_local;
wire [31:0] local_bb3_and226_i;

assign local_bb3_and226_i = ((rnode_337to338_bb3__45_i578_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and271_i_stall_local;
wire [31:0] local_bb3_and271_i;

assign local_bb3_and271_i = ((rnode_337to338_bb3__45_i578_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb3_shr272_i_valid_out;
wire local_bb3_shr272_i_stall_in;
wire local_bb3_shr272_i_inputs_ready;
wire local_bb3_shr272_i_stall_local;
wire [31:0] local_bb3_shr272_i;

assign local_bb3_shr272_i_inputs_ready = rnode_337to338_bb3__45_i578_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_shr272_i = ((rnode_337to338_bb3__45_i578_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb3_shr272_i_valid_out = 1'b1;
assign rnode_337to338_bb3__45_i578_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_391_392_0_inputs_ready;
 reg SFC_1_VALID_391_392_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_391_392_0_stall_in;
wire SFC_1_VALID_391_392_0_output_regs_ready;
 reg SFC_1_VALID_391_392_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_391_392_0_causedstall;

assign SFC_1_VALID_391_392_0_inputs_ready = 1'b1;
assign SFC_1_VALID_391_392_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_390_391_0_stall_in = 1'b0;
assign SFC_1_VALID_391_392_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_391_392_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_391_392_0_output_regs_ready)
		begin
			SFC_1_VALID_391_392_0_NO_SHIFT_REG <= SFC_1_VALID_390_391_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_notlhs_i582_stall_local;
wire local_bb3_notlhs_i582;

assign local_bb3_notlhs_i582 = ((local_bb3_and248_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp227_i_stall_local;
wire local_bb3_cmp227_i;

assign local_bb3_cmp227_i = ((local_bb3_and226_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp297_i_stall_local;
wire local_bb3_cmp297_i;

assign local_bb3_cmp297_i = ((local_bb3_and271_i & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp297_i_valid_out;
wire local_bb3_cmp297_i_stall_in;
wire local_bb3_cmp300_i_valid_out;
wire local_bb3_cmp300_i_stall_in;
wire local_bb3_cmp300_i_inputs_ready;
wire local_bb3_cmp300_i_stall_local;
wire local_bb3_cmp300_i;

assign local_bb3_cmp300_i_inputs_ready = rnode_337to338_bb3__45_i578_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_cmp300_i = ((local_bb3_and271_i & 32'h7) == 32'h4);
assign local_bb3_cmp297_i_valid_out = 1'b1;
assign local_bb3_cmp300_i_valid_out = 1'b1;
assign rnode_337to338_bb3__45_i578_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb3_shr272_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_338to339_bb3_shr272_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_338to339_bb3_shr272_i_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3_shr272_i_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_338to339_bb3_shr272_i_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_shr272_i_0_valid_out_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_shr272_i_0_stall_in_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_shr272_i_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb3_shr272_i_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb3_shr272_i_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb3_shr272_i_0_stall_in_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb3_shr272_i_0_valid_out_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb3_shr272_i_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in((local_bb3_shr272_i & 32'h1FFFFFF)),
	.data_out(rnode_338to339_bb3_shr272_i_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb3_shr272_i_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb3_shr272_i_0_reg_339_fifo.DATA_WIDTH = 32;
defparam rnode_338to339_bb3_shr272_i_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb3_shr272_i_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_338to339_bb3_shr272_i_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr272_i_stall_in = 1'b0;
assign rnode_338to339_bb3_shr272_i_0_NO_SHIFT_REG = rnode_338to339_bb3_shr272_i_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3_shr272_i_0_stall_in_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_shr272_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_392_393_0_inputs_ready;
 reg SFC_1_VALID_392_393_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_392_393_0_stall_in;
wire SFC_1_VALID_392_393_0_output_regs_ready;
 reg SFC_1_VALID_392_393_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_392_393_0_causedstall;

assign SFC_1_VALID_392_393_0_inputs_ready = 1'b1;
assign SFC_1_VALID_392_393_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_391_392_0_stall_in = 1'b0;
assign SFC_1_VALID_392_393_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_392_393_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_392_393_0_output_regs_ready)
		begin
			SFC_1_VALID_392_393_0_NO_SHIFT_REG <= SFC_1_VALID_391_392_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_not__46_i584_stall_local;
wire local_bb3_not__46_i584;

assign local_bb3_not__46_i584 = (local_bb3_notrhs_i583 | local_bb3_notlhs_i582);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp227_not_i_stall_local;
wire local_bb3_cmp227_not_i;

assign local_bb3_cmp227_not_i = (local_bb3_cmp227_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb3_cmp297_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp297_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp297_i_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp297_i_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp297_i_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp297_i_0_valid_out_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp297_i_0_stall_in_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp297_i_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb3_cmp297_i_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb3_cmp297_i_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb3_cmp297_i_0_stall_in_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb3_cmp297_i_0_valid_out_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb3_cmp297_i_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in(local_bb3_cmp297_i),
	.data_out(rnode_338to339_bb3_cmp297_i_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb3_cmp297_i_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb3_cmp297_i_0_reg_339_fifo.DATA_WIDTH = 1;
defparam rnode_338to339_bb3_cmp297_i_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb3_cmp297_i_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_338to339_bb3_cmp297_i_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp297_i_stall_in = 1'b0;
assign rnode_338to339_bb3_cmp297_i_0_NO_SHIFT_REG = rnode_338to339_bb3_cmp297_i_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3_cmp297_i_0_stall_in_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_cmp297_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb3_cmp300_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp300_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp300_i_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp300_i_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp300_i_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp300_i_0_valid_out_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp300_i_0_stall_in_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_cmp300_i_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb3_cmp300_i_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb3_cmp300_i_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb3_cmp300_i_0_stall_in_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb3_cmp300_i_0_valid_out_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb3_cmp300_i_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in(local_bb3_cmp300_i),
	.data_out(rnode_338to339_bb3_cmp300_i_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb3_cmp300_i_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb3_cmp300_i_0_reg_339_fifo.DATA_WIDTH = 1;
defparam rnode_338to339_bb3_cmp300_i_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb3_cmp300_i_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_338to339_bb3_cmp300_i_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp300_i_stall_in = 1'b0;
assign rnode_338to339_bb3_cmp300_i_0_NO_SHIFT_REG = rnode_338to339_bb3_cmp300_i_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3_cmp300_i_0_stall_in_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_cmp300_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and273_i_stall_local;
wire [31:0] local_bb3_and273_i;

assign local_bb3_and273_i = ((rnode_338to339_bb3_shr272_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements a registered operation.
// 
wire SFC_1_VALID_393_394_0_inputs_ready;
 reg SFC_1_VALID_393_394_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_393_394_0_stall_in;
wire SFC_1_VALID_393_394_0_output_regs_ready;
 reg SFC_1_VALID_393_394_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_393_394_0_causedstall;

assign SFC_1_VALID_393_394_0_inputs_ready = 1'b1;
assign SFC_1_VALID_393_394_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_392_393_0_stall_in = 1'b0;
assign SFC_1_VALID_393_394_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_393_394_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_393_394_0_output_regs_ready)
		begin
			SFC_1_VALID_393_394_0_NO_SHIFT_REG <= SFC_1_VALID_392_393_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3__47_i585_stall_local;
wire local_bb3__47_i585;

assign local_bb3__47_i585 = (local_bb3_cmp227_i | local_bb3_not__46_i584);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge12_i579_stall_local;
wire local_bb3_brmerge12_i579;

assign local_bb3_brmerge12_i579 = (local_bb3_cmp227_not_i | rnode_337to338_bb3_not_cmp38_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot263__i_stall_local;
wire local_bb3_lnot263__i;

assign local_bb3_lnot263__i = (local_bb3_cmp259_i & local_bb3_cmp227_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp29749_i_stall_local;
wire [31:0] local_bb3_cmp29749_i;

assign local_bb3_cmp29749_i[31:1] = 31'h0;
assign local_bb3_cmp29749_i[0] = rnode_338to339_bb3_cmp297_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_conv301_i_stall_local;
wire [31:0] local_bb3_conv301_i;

assign local_bb3_conv301_i[31:1] = 31'h0;
assign local_bb3_conv301_i[0] = rnode_338to339_bb3_cmp300_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or275_i587_stall_local;
wire [31:0] local_bb3_or275_i587;

assign local_bb3_or275_i587 = ((local_bb3_and273_i & 32'h7FFFFF) | (local_bb3_shl274_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb3_resultSign_0_i580_stall_local;
wire [31:0] local_bb3_resultSign_0_i580;

assign local_bb3_resultSign_0_i580 = (local_bb3_brmerge12_i579 ? (rnode_337to338_bb3_and35_i520_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_resultSign_0_i580_valid_out;
wire local_bb3_resultSign_0_i580_stall_in;
wire local_bb3__47_i585_valid_out;
wire local_bb3__47_i585_stall_in;
wire local_bb3_or2672_i_valid_out;
wire local_bb3_or2672_i_stall_in;
wire local_bb3_or2672_i_inputs_ready;
wire local_bb3_or2672_i_stall_local;
wire local_bb3_or2672_i;

assign local_bb3_or2672_i_inputs_ready = (rnode_337to338_bb3_and35_i520_0_valid_out_NO_SHIFT_REG & rnode_337to338_bb3_not_cmp38_i_0_valid_out_NO_SHIFT_REG & rnode_337to338_bb3_add246_i_0_valid_out_0_NO_SHIFT_REG & rnode_337to338_bb3_and251_i_0_valid_out_NO_SHIFT_REG & rnode_337to338_bb3__45_i578_0_valid_out_0_NO_SHIFT_REG & rnode_337to338_bb3_add246_i_0_valid_out_1_NO_SHIFT_REG & rnode_337to338_bb3_var__u28_0_valid_out_NO_SHIFT_REG);
assign local_bb3_or2672_i = (rnode_337to338_bb3_var__u28_0_NO_SHIFT_REG | local_bb3_lnot263__i);
assign local_bb3_resultSign_0_i580_valid_out = 1'b1;
assign local_bb3__47_i585_valid_out = 1'b1;
assign local_bb3_or2672_i_valid_out = 1'b1;
assign rnode_337to338_bb3_and35_i520_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_not_cmp38_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_add246_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_and251_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3__45_i578_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_add246_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_337to338_bb3_var__u28_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb3_resultSign_0_i580_0_valid_out_NO_SHIFT_REG;
 logic rnode_338to339_bb3_resultSign_0_i580_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_338to339_bb3_resultSign_0_i580_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3_resultSign_0_i580_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_338to339_bb3_resultSign_0_i580_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_resultSign_0_i580_0_valid_out_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_resultSign_0_i580_0_stall_in_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_resultSign_0_i580_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb3_resultSign_0_i580_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb3_resultSign_0_i580_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb3_resultSign_0_i580_0_stall_in_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb3_resultSign_0_i580_0_valid_out_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb3_resultSign_0_i580_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in((local_bb3_resultSign_0_i580 & 32'h80000000)),
	.data_out(rnode_338to339_bb3_resultSign_0_i580_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb3_resultSign_0_i580_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb3_resultSign_0_i580_0_reg_339_fifo.DATA_WIDTH = 32;
defparam rnode_338to339_bb3_resultSign_0_i580_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb3_resultSign_0_i580_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_338to339_bb3_resultSign_0_i580_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_resultSign_0_i580_stall_in = 1'b0;
assign rnode_338to339_bb3_resultSign_0_i580_0_NO_SHIFT_REG = rnode_338to339_bb3_resultSign_0_i580_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3_resultSign_0_i580_0_stall_in_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_resultSign_0_i580_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb3__47_i585_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_valid_out_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_stall_in_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3__47_i585_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb3__47_i585_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb3__47_i585_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb3__47_i585_0_stall_in_0_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb3__47_i585_0_valid_out_0_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb3__47_i585_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in(local_bb3__47_i585),
	.data_out(rnode_338to339_bb3__47_i585_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb3__47_i585_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb3__47_i585_0_reg_339_fifo.DATA_WIDTH = 1;
defparam rnode_338to339_bb3__47_i585_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb3__47_i585_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_338to339_bb3__47_i585_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__47_i585_stall_in = 1'b0;
assign rnode_338to339_bb3__47_i585_0_stall_in_0_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__47_i585_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3__47_i585_0_NO_SHIFT_REG = rnode_338to339_bb3__47_i585_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3__47_i585_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3__47_i585_1_NO_SHIFT_REG = rnode_338to339_bb3__47_i585_0_reg_339_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb3_or2672_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_1_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_2_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_valid_out_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_stall_in_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb3_or2672_i_0_stall_out_reg_339_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb3_or2672_i_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb3_or2672_i_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb3_or2672_i_0_stall_in_0_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb3_or2672_i_0_valid_out_0_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb3_or2672_i_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in(local_bb3_or2672_i),
	.data_out(rnode_338to339_bb3_or2672_i_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb3_or2672_i_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb3_or2672_i_0_reg_339_fifo.DATA_WIDTH = 1;
defparam rnode_338to339_bb3_or2672_i_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb3_or2672_i_0_reg_339_fifo.IMPL = "shift_reg";

assign rnode_338to339_bb3_or2672_i_0_reg_339_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or2672_i_stall_in = 1'b0;
assign rnode_338to339_bb3_or2672_i_0_stall_in_0_reg_339_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_or2672_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3_or2672_i_0_NO_SHIFT_REG = rnode_338to339_bb3_or2672_i_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3_or2672_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3_or2672_i_1_NO_SHIFT_REG = rnode_338to339_bb3_or2672_i_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb3_or2672_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_338to339_bb3_or2672_i_2_NO_SHIFT_REG = rnode_338to339_bb3_or2672_i_0_reg_339_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or276_i_stall_local;
wire [31:0] local_bb3_or276_i;

assign local_bb3_or276_i = ((local_bb3_or275_i587 & 32'h7FFFFFFF) | (rnode_338to339_bb3_resultSign_0_i580_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u38_stall_local;
wire [31:0] local_bb3_var__u38;

assign local_bb3_var__u38[31:1] = 31'h0;
assign local_bb3_var__u38[0] = rnode_338to339_bb3__47_i585_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or2814_i_stall_local;
wire local_bb3_or2814_i;

assign local_bb3_or2814_i = (rnode_338to339_bb3__47_i585_0_NO_SHIFT_REG | rnode_338to339_bb3_or2672_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_or2885_i_stall_local;
wire local_bb3_or2885_i;

assign local_bb3_or2885_i = (rnode_338to339_bb3_or2672_i_1_NO_SHIFT_REG | rnode_338to339_bb3__26_i533_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u39_stall_local;
wire [31:0] local_bb3_var__u39;

assign local_bb3_var__u39[31:1] = 31'h0;
assign local_bb3_var__u39[0] = rnode_338to339_bb3_or2672_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext315_i_stall_local;
wire [31:0] local_bb3_lnot_ext315_i;

assign local_bb3_lnot_ext315_i = ((local_bb3_var__u38 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cond283_i_stall_local;
wire [31:0] local_bb3_cond283_i;

assign local_bb3_cond283_i = (local_bb3_or2814_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cond290_i_stall_local;
wire [31:0] local_bb3_cond290_i;

assign local_bb3_cond290_i = (local_bb3_or2885_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext311_i_stall_local;
wire [31:0] local_bb3_lnot_ext311_i;

assign local_bb3_lnot_ext311_i = ((local_bb3_var__u39 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and294_i_stall_local;
wire [31:0] local_bb3_and294_i;

assign local_bb3_and294_i = ((local_bb3_cond283_i | 32'h80000000) & local_bb3_or276_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or295_i588_stall_local;
wire [31:0] local_bb3_or295_i588;

assign local_bb3_or295_i588 = ((local_bb3_cond290_i & 32'h7F800000) | (local_bb3_cond293_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_0_i591_stall_local;
wire [31:0] local_bb3_reduction_0_i591;

assign local_bb3_reduction_0_i591 = ((local_bb3_lnot_ext311_i & 32'h1) & (local_bb3_lnot_ext_i590 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and303_i_stall_local;
wire [31:0] local_bb3_and303_i;

assign local_bb3_and303_i = ((local_bb3_conv301_i & 32'h1) & local_bb3_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or296_i_stall_local;
wire [31:0] local_bb3_or296_i;

assign local_bb3_or296_i = ((local_bb3_or295_i588 & 32'h7FC00000) | local_bb3_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb3_lor_ext_i589_stall_local;
wire [31:0] local_bb3_lor_ext_i589;

assign local_bb3_lor_ext_i589 = ((local_bb3_cmp29749_i & 32'h1) | (local_bb3_and303_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_1_i592_stall_local;
wire [31:0] local_bb3_reduction_1_i592;

assign local_bb3_reduction_1_i592 = ((local_bb3_lnot_ext315_i & 32'h1) & (local_bb3_lor_ext_i589 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_2_i593_stall_local;
wire [31:0] local_bb3_reduction_2_i593;

assign local_bb3_reduction_2_i593 = ((local_bb3_reduction_0_i591 & 32'h1) & (local_bb3_reduction_1_i592 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_add321_i_stall_local;
wire [31:0] local_bb3_add321_i;

assign local_bb3_add321_i = ((local_bb3_reduction_2_i593 & 32'h1) + local_bb3_or296_i);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i404_stall_local;
wire [31:0] local_bb3_shr_i404;

assign local_bb3_shr_i404 = (local_bb3_add321_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shr2_i406_stall_local;
wire [31:0] local_bb3_shr2_i406;

assign local_bb3_shr2_i406 = (local_bb3_add321_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and5_i410_stall_local;
wire [31:0] local_bb3_and5_i410;

assign local_bb3_and5_i410 = (local_bb3_add321_i & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and6_i411_stall_local;
wire [31:0] local_bb3_and6_i411;

assign local_bb3_and6_i411 = (local_bb3_add321_i & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i438_stall_local;
wire [31:0] local_bb3_or_i438;

assign local_bb3_or_i438 = ((local_bb3_and5_i410 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_or47_i439_stall_local;
wire [31:0] local_bb3_or47_i439;

assign local_bb3_or47_i439 = ((local_bb3_and6_i411 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_conv_i_i440_stall_local;
wire [63:0] local_bb3_conv_i_i440;

assign local_bb3_conv_i_i440[63:32] = 32'h0;
assign local_bb3_conv_i_i440[31:0] = ((local_bb3_or_i438 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i404_valid_out;
wire local_bb3_shr_i404_stall_in;
wire local_bb3_shr2_i406_valid_out;
wire local_bb3_shr2_i406_stall_in;
wire local_bb3_and5_i410_valid_out_1;
wire local_bb3_and5_i410_stall_in_1;
wire local_bb3_and6_i411_valid_out_1;
wire local_bb3_and6_i411_stall_in_1;
wire local_bb3_conv_i_i440_valid_out;
wire local_bb3_conv_i_i440_stall_in;
wire local_bb3_conv1_i_i441_valid_out;
wire local_bb3_conv1_i_i441_stall_in;
wire local_bb3_conv1_i_i441_inputs_ready;
wire local_bb3_conv1_i_i441_stall_local;
wire [63:0] local_bb3_conv1_i_i441;

assign local_bb3_conv1_i_i441_inputs_ready = (rnode_337to339_bb3_and270_i586_0_valid_out_NO_SHIFT_REG & rnode_338to339_bb3_resultSign_0_i580_0_valid_out_NO_SHIFT_REG & rnode_338to339_bb3_or2672_i_0_valid_out_1_NO_SHIFT_REG & rnode_338to339_bb3__26_i533_0_valid_out_0_NO_SHIFT_REG & rnode_338to339_bb3__26_i533_0_valid_out_1_NO_SHIFT_REG & rnode_338to339_bb3__47_i585_0_valid_out_0_NO_SHIFT_REG & rnode_338to339_bb3_or2672_i_0_valid_out_0_NO_SHIFT_REG & rnode_338to339_bb3__26_i533_0_valid_out_2_NO_SHIFT_REG & rnode_338to339_bb3_or2672_i_0_valid_out_2_NO_SHIFT_REG & rnode_338to339_bb3_shr272_i_0_valid_out_NO_SHIFT_REG & rnode_338to339_bb3__47_i585_0_valid_out_1_NO_SHIFT_REG & rnode_338to339_bb3_cmp297_i_0_valid_out_NO_SHIFT_REG & rnode_338to339_bb3_cmp300_i_0_valid_out_NO_SHIFT_REG);
assign local_bb3_conv1_i_i441[63:32] = 32'h0;
assign local_bb3_conv1_i_i441[31:0] = ((local_bb3_or47_i439 & 32'hFFFFFF) | 32'h800000);
assign local_bb3_shr_i404_valid_out = 1'b1;
assign local_bb3_shr2_i406_valid_out = 1'b1;
assign local_bb3_and5_i410_valid_out_1 = 1'b1;
assign local_bb3_and6_i411_valid_out_1 = 1'b1;
assign local_bb3_conv_i_i440_valid_out = 1'b1;
assign local_bb3_conv1_i_i441_valid_out = 1'b1;
assign rnode_337to339_bb3_and270_i586_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_resultSign_0_i580_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_or2672_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__26_i533_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__26_i533_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__47_i585_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_or2672_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__26_i533_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_or2672_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_shr272_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3__47_i585_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_cmp297_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_338to339_bb3_cmp300_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_339to340_bb3_shr_i404_0_valid_out_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr_i404_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_shr_i404_0_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr_i404_0_reg_340_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_shr_i404_0_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr_i404_0_valid_out_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr_i404_0_stall_in_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr_i404_0_stall_out_reg_340_NO_SHIFT_REG;

acl_data_fifo rnode_339to340_bb3_shr_i404_0_reg_340_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_339to340_bb3_shr_i404_0_reg_340_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_339to340_bb3_shr_i404_0_stall_in_reg_340_NO_SHIFT_REG),
	.valid_out(rnode_339to340_bb3_shr_i404_0_valid_out_reg_340_NO_SHIFT_REG),
	.stall_out(rnode_339to340_bb3_shr_i404_0_stall_out_reg_340_NO_SHIFT_REG),
	.data_in((local_bb3_shr_i404 & 32'h1FF)),
	.data_out(rnode_339to340_bb3_shr_i404_0_reg_340_NO_SHIFT_REG)
);

defparam rnode_339to340_bb3_shr_i404_0_reg_340_fifo.DEPTH = 1;
defparam rnode_339to340_bb3_shr_i404_0_reg_340_fifo.DATA_WIDTH = 32;
defparam rnode_339to340_bb3_shr_i404_0_reg_340_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_339to340_bb3_shr_i404_0_reg_340_fifo.IMPL = "shift_reg";

assign rnode_339to340_bb3_shr_i404_0_reg_340_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr_i404_stall_in = 1'b0;
assign rnode_339to340_bb3_shr_i404_0_NO_SHIFT_REG = rnode_339to340_bb3_shr_i404_0_reg_340_NO_SHIFT_REG;
assign rnode_339to340_bb3_shr_i404_0_stall_in_reg_340_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_shr_i404_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_339to340_bb3_shr2_i406_0_valid_out_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr2_i406_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_shr2_i406_0_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr2_i406_0_reg_340_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_shr2_i406_0_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr2_i406_0_valid_out_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr2_i406_0_stall_in_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_shr2_i406_0_stall_out_reg_340_NO_SHIFT_REG;

acl_data_fifo rnode_339to340_bb3_shr2_i406_0_reg_340_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_339to340_bb3_shr2_i406_0_reg_340_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_339to340_bb3_shr2_i406_0_stall_in_reg_340_NO_SHIFT_REG),
	.valid_out(rnode_339to340_bb3_shr2_i406_0_valid_out_reg_340_NO_SHIFT_REG),
	.stall_out(rnode_339to340_bb3_shr2_i406_0_stall_out_reg_340_NO_SHIFT_REG),
	.data_in((local_bb3_shr2_i406 & 32'h1FF)),
	.data_out(rnode_339to340_bb3_shr2_i406_0_reg_340_NO_SHIFT_REG)
);

defparam rnode_339to340_bb3_shr2_i406_0_reg_340_fifo.DEPTH = 1;
defparam rnode_339to340_bb3_shr2_i406_0_reg_340_fifo.DATA_WIDTH = 32;
defparam rnode_339to340_bb3_shr2_i406_0_reg_340_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_339to340_bb3_shr2_i406_0_reg_340_fifo.IMPL = "shift_reg";

assign rnode_339to340_bb3_shr2_i406_0_reg_340_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr2_i406_stall_in = 1'b0;
assign rnode_339to340_bb3_shr2_i406_0_NO_SHIFT_REG = rnode_339to340_bb3_shr2_i406_0_reg_340_NO_SHIFT_REG;
assign rnode_339to340_bb3_shr2_i406_0_stall_in_reg_340_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_shr2_i406_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_339to340_bb3_and5_i410_0_valid_out_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and5_i410_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_and5_i410_0_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and5_i410_0_reg_340_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_and5_i410_0_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and5_i410_0_valid_out_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and5_i410_0_stall_in_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and5_i410_0_stall_out_reg_340_NO_SHIFT_REG;

acl_data_fifo rnode_339to340_bb3_and5_i410_0_reg_340_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_339to340_bb3_and5_i410_0_reg_340_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_339to340_bb3_and5_i410_0_stall_in_reg_340_NO_SHIFT_REG),
	.valid_out(rnode_339to340_bb3_and5_i410_0_valid_out_reg_340_NO_SHIFT_REG),
	.stall_out(rnode_339to340_bb3_and5_i410_0_stall_out_reg_340_NO_SHIFT_REG),
	.data_in((local_bb3_and5_i410 & 32'h7FFFFF)),
	.data_out(rnode_339to340_bb3_and5_i410_0_reg_340_NO_SHIFT_REG)
);

defparam rnode_339to340_bb3_and5_i410_0_reg_340_fifo.DEPTH = 1;
defparam rnode_339to340_bb3_and5_i410_0_reg_340_fifo.DATA_WIDTH = 32;
defparam rnode_339to340_bb3_and5_i410_0_reg_340_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_339to340_bb3_and5_i410_0_reg_340_fifo.IMPL = "shift_reg";

assign rnode_339to340_bb3_and5_i410_0_reg_340_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and5_i410_stall_in_1 = 1'b0;
assign rnode_339to340_bb3_and5_i410_0_NO_SHIFT_REG = rnode_339to340_bb3_and5_i410_0_reg_340_NO_SHIFT_REG;
assign rnode_339to340_bb3_and5_i410_0_stall_in_reg_340_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_and5_i410_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_339to340_bb3_and6_i411_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_and6_i411_0_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_and6_i411_1_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_and6_i411_2_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_reg_340_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_339to340_bb3_and6_i411_0_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_valid_out_0_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_stall_in_0_reg_340_NO_SHIFT_REG;
 logic rnode_339to340_bb3_and6_i411_0_stall_out_reg_340_NO_SHIFT_REG;

acl_data_fifo rnode_339to340_bb3_and6_i411_0_reg_340_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_339to340_bb3_and6_i411_0_reg_340_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_339to340_bb3_and6_i411_0_stall_in_0_reg_340_NO_SHIFT_REG),
	.valid_out(rnode_339to340_bb3_and6_i411_0_valid_out_0_reg_340_NO_SHIFT_REG),
	.stall_out(rnode_339to340_bb3_and6_i411_0_stall_out_reg_340_NO_SHIFT_REG),
	.data_in((local_bb3_and6_i411 & 32'h7FFFFF)),
	.data_out(rnode_339to340_bb3_and6_i411_0_reg_340_NO_SHIFT_REG)
);

defparam rnode_339to340_bb3_and6_i411_0_reg_340_fifo.DEPTH = 1;
defparam rnode_339to340_bb3_and6_i411_0_reg_340_fifo.DATA_WIDTH = 32;
defparam rnode_339to340_bb3_and6_i411_0_reg_340_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_339to340_bb3_and6_i411_0_reg_340_fifo.IMPL = "shift_reg";

assign rnode_339to340_bb3_and6_i411_0_reg_340_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and6_i411_stall_in_1 = 1'b0;
assign rnode_339to340_bb3_and6_i411_0_stall_in_0_reg_340_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_and6_i411_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_339to340_bb3_and6_i411_0_NO_SHIFT_REG = rnode_339to340_bb3_and6_i411_0_reg_340_NO_SHIFT_REG;
assign rnode_339to340_bb3_and6_i411_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_339to340_bb3_and6_i411_1_NO_SHIFT_REG = rnode_339to340_bb3_and6_i411_0_reg_340_NO_SHIFT_REG;
assign rnode_339to340_bb3_and6_i411_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_339to340_bb3_and6_i411_2_NO_SHIFT_REG = rnode_339to340_bb3_and6_i411_0_reg_340_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb3_mul_i_i442_inputs_ready;
 reg local_bb3_mul_i_i442_valid_out_0_NO_SHIFT_REG;
wire local_bb3_mul_i_i442_stall_in_0;
 reg local_bb3_mul_i_i442_valid_out_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i442_stall_in_1;
wire local_bb3_mul_i_i442_output_regs_ready;
wire [63:0] local_bb3_mul_i_i442;
 reg local_bb3_mul_i_i442_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_mul_i_i442_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i442_causedstall;

acl_int_mult int_module_local_bb3_mul_i_i442 (
	.clock(clock),
	.dataa(((local_bb3_conv1_i_i441 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb3_conv_i_i440 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb3_mul_i_i442_output_regs_ready),
	.result(local_bb3_mul_i_i442)
);

defparam int_module_local_bb3_mul_i_i442.INPUT1_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i442.INPUT2_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i442.OUTPUT_WIDTH = 64;
defparam int_module_local_bb3_mul_i_i442.LATENCY = 3;
defparam int_module_local_bb3_mul_i_i442.SIGNED = 0;

assign local_bb3_mul_i_i442_inputs_ready = 1'b1;
assign local_bb3_mul_i_i442_output_regs_ready = 1'b1;
assign local_bb3_conv1_i_i441_stall_in = 1'b0;
assign local_bb3_conv_i_i440_stall_in = 1'b0;
assign local_bb3_mul_i_i442_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i442_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i442_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i442_output_regs_ready)
		begin
			local_bb3_mul_i_i442_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i442_valid_pipe_1_NO_SHIFT_REG <= local_bb3_mul_i_i442_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i442_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i442_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i442_output_regs_ready)
		begin
			local_bb3_mul_i_i442_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i442_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_mul_i_i442_stall_in_0))
			begin
				local_bb3_mul_i_i442_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_mul_i_i442_stall_in_1))
			begin
				local_bb3_mul_i_i442_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and_i405_stall_local;
wire [31:0] local_bb3_and_i405;

assign local_bb3_and_i405 = ((rnode_339to340_bb3_shr_i404_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and3_i407_stall_local;
wire [31:0] local_bb3_and3_i407;

assign local_bb3_and3_i407 = ((rnode_339to340_bb3_shr2_i406_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_i416_stall_local;
wire local_bb3_lnot14_i416;

assign local_bb3_lnot14_i416 = ((rnode_339to340_bb3_and5_i410_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_i417_stall_local;
wire local_bb3_lnot17_i417;

assign local_bb3_lnot17_i417 = ((rnode_339to340_bb3_and6_i411_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_conv3_i_i443_stall_local;
wire [31:0] local_bb3_conv3_i_i443;
wire [63:0] local_bb3_conv3_i_i443$ps;

assign local_bb3_conv3_i_i443$ps = (local_bb3_mul_i_i442 & 64'hFFFFFFFFFFFF);
assign local_bb3_conv3_i_i443 = local_bb3_conv3_i_i443$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_var__u40_stall_local;
wire [63:0] local_bb3_var__u40;

assign local_bb3_var__u40 = ((local_bb3_mul_i_i442 & 64'hFFFFFFFFFFFF) >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_i412_stall_local;
wire local_bb3_lnot_i412;

assign local_bb3_lnot_i412 = ((local_bb3_and_i405 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i414_stall_local;
wire local_bb3_cmp_i414;

assign local_bb3_cmp_i414 = ((local_bb3_and_i405 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u41_stall_local;
wire [31:0] local_bb3_var__u41;

assign local_bb3_var__u41 = ((rnode_339to340_bb3_and6_i411_2_NO_SHIFT_REG & 32'h7FFFFF) | (local_bb3_and_i405 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot8_i413_stall_local;
wire local_bb3_lnot8_i413;

assign local_bb3_lnot8_i413 = ((local_bb3_and3_i407 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_i415_stall_local;
wire local_bb3_cmp11_i415;

assign local_bb3_cmp11_i415 = ((local_bb3_and3_i407 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u42_stall_local;
wire [31:0] local_bb3_var__u42;

assign local_bb3_var__u42 = ((local_bb3_and3_i407 & 32'hFF) | (rnode_339to340_bb3_and6_i411_1_NO_SHIFT_REG & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_add_i449_stall_local;
wire [31:0] local_bb3_add_i449;

assign local_bb3_add_i449 = ((local_bb3_and3_i407 & 32'hFF) + (local_bb3_and_i405 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_not_i435_stall_local;
wire local_bb3_lnot14_not_i435;

assign local_bb3_lnot14_not_i435 = (local_bb3_lnot14_i416 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_not_i421_stall_local;
wire local_bb3_lnot17_not_i421;

assign local_bb3_lnot17_not_i421 = (local_bb3_lnot17_i417 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i16_i446_stall_local;
wire [31:0] local_bb3_shr_i16_i446;

assign local_bb3_shr_i16_i446 = (local_bb3_conv3_i_i443 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i18_i448_stall_local;
wire [31:0] local_bb3_shl1_i18_i448;

assign local_bb3_shl1_i18_i448 = (local_bb3_conv3_i_i443 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u43_stall_local;
wire [31:0] local_bb3_var__u43;

assign local_bb3_var__u43 = (local_bb3_conv3_i_i443 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i_i456_stall_local;
wire [31:0] local_bb3_shl1_i_i456;

assign local_bb3_shl1_i_i456 = (local_bb3_conv3_i_i443 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb3__tr_i444_stall_local;
wire [31:0] local_bb3__tr_i444;
wire [63:0] local_bb3__tr_i444$ps;

assign local_bb3__tr_i444$ps = (local_bb3_var__u40 & 64'hFFFFFF);
assign local_bb3__tr_i444 = local_bb3__tr_i444$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_var__u44_stall_local;
wire local_bb3_var__u44;

assign local_bb3_var__u44 = ((local_bb3_var__u41 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_0_i467_stall_local;
wire local_bb3_reduction_0_i467;

assign local_bb3_reduction_0_i467 = (local_bb3_lnot_i412 | local_bb3_lnot8_i413);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge8_demorgan_i418_stall_local;
wire local_bb3_brmerge8_demorgan_i418;

assign local_bb3_brmerge8_demorgan_i418 = (local_bb3_cmp11_i415 & local_bb3_lnot17_i417);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_not_i422_stall_local;
wire local_bb3_cmp11_not_i422;

assign local_bb3_cmp11_not_i422 = (local_bb3_cmp11_i415 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u45_stall_local;
wire local_bb3_var__u45;

assign local_bb3_var__u45 = (local_bb3_cmp_i414 | local_bb3_cmp11_i415);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u46_stall_local;
wire local_bb3_var__u46;

assign local_bb3_var__u46 = ((local_bb3_var__u42 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__28_i436_stall_local;
wire local_bb3__28_i436;

assign local_bb3__28_i436 = (local_bb3_cmp_i414 & local_bb3_lnot14_not_i435);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i_i454_stall_local;
wire [31:0] local_bb3_shr_i_i454;

assign local_bb3_shr_i_i454 = ((local_bb3_var__u43 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i15_i445_stall_local;
wire [31:0] local_bb3_shl_i15_i445;

assign local_bb3_shl_i15_i445 = ((local_bb3__tr_i444 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb3_and48_i450_stall_local;
wire [31:0] local_bb3_and48_i450;

assign local_bb3_and48_i450 = ((local_bb3__tr_i444 & 32'hFFFFFF) & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge10_demorgan_i419_stall_local;
wire local_bb3_brmerge10_demorgan_i419;

assign local_bb3_brmerge10_demorgan_i419 = (local_bb3_brmerge8_demorgan_i418 & local_bb3_lnot_i412);

// This section implements an unregistered operation.
// 
wire local_bb3__mux9_mux_i420_stall_local;
wire local_bb3__mux9_mux_i420;

assign local_bb3__mux9_mux_i420 = (local_bb3_brmerge8_demorgan_i418 ^ local_bb3_cmp11_i415);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge3_i423_stall_local;
wire local_bb3_brmerge3_i423;

assign local_bb3_brmerge3_i423 = (local_bb3_var__u46 | local_bb3_cmp11_not_i422);

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_i425_stall_local;
wire local_bb3__mux_mux_i425;

assign local_bb3__mux_mux_i425 = (local_bb3_var__u46 | local_bb3_cmp11_i415);

// This section implements an unregistered operation.
// 
wire local_bb3__not_i427_stall_local;
wire local_bb3__not_i427;

assign local_bb3__not_i427 = (local_bb3_var__u46 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i17_i447_stall_local;
wire [31:0] local_bb3_or_i17_i447;

assign local_bb3_or_i17_i447 = ((local_bb3_shl_i15_i445 & 32'hFFFF00) | (local_bb3_shr_i16_i446 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool49_i451_stall_local;
wire local_bb3_tobool49_i451;

assign local_bb3_tobool49_i451 = ((local_bb3_and48_i450 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__26_demorgan_i433_stall_local;
wire local_bb3__26_demorgan_i433;

assign local_bb3__26_demorgan_i433 = (local_bb3_cmp_i414 | local_bb3_brmerge10_demorgan_i419);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge5_i424_stall_local;
wire local_bb3_brmerge5_i424;

assign local_bb3_brmerge5_i424 = (local_bb3_brmerge3_i423 | local_bb3_lnot17_not_i421);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_3_i428_stall_local;
wire local_bb3_reduction_3_i428;

assign local_bb3_reduction_3_i428 = (local_bb3_cmp11_i415 & local_bb3__not_i427);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i_i453_stall_local;
wire [31:0] local_bb3_shl_i_i453;

assign local_bb3_shl_i_i453 = ((local_bb3_or_i17_i447 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_mux_i426_stall_local;
wire local_bb3__mux_mux_mux_i426;

assign local_bb3__mux_mux_mux_i426 = (local_bb3_brmerge5_i424 & local_bb3__mux_mux_i425);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_5_i429_stall_local;
wire local_bb3_reduction_5_i429;

assign local_bb3_reduction_5_i429 = (local_bb3_lnot14_i416 & local_bb3_reduction_3_i428);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i_i455_stall_local;
wire [31:0] local_bb3_or_i_i455;

assign local_bb3_or_i_i455 = ((local_bb3_shl_i_i453 & 32'h1FFFFFE) | (local_bb3_shr_i_i454 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_6_i430_stall_local;
wire local_bb3_reduction_6_i430;

assign local_bb3_reduction_6_i430 = (local_bb3_var__u44 & local_bb3_reduction_5_i429);

// This section implements an unregistered operation.
// 
wire local_bb3__24_i431_stall_local;
wire local_bb3__24_i431;

assign local_bb3__24_i431 = (local_bb3_cmp_i414 ? local_bb3_reduction_6_i430 : local_bb3_brmerge10_demorgan_i419);

// This section implements an unregistered operation.
// 
wire local_bb3__25_i432_stall_local;
wire local_bb3__25_i432;

assign local_bb3__25_i432 = (local_bb3__24_i431 ? local_bb3_lnot14_i416 : local_bb3__mux_mux_mux_i426);

// This section implements an unregistered operation.
// 
wire local_bb3__27_i434_stall_local;
wire local_bb3__27_i434;

assign local_bb3__27_i434 = (local_bb3__26_demorgan_i433 ? local_bb3__25_i432 : local_bb3__mux9_mux_i420);

// This section implements an unregistered operation.
// 
wire local_bb3_add_i449_valid_out;
wire local_bb3_add_i449_stall_in;
wire local_bb3_reduction_0_i467_valid_out;
wire local_bb3_reduction_0_i467_stall_in;
wire local_bb3_var__u45_valid_out;
wire local_bb3_var__u45_stall_in;
wire local_bb3__29_i437_valid_out;
wire local_bb3__29_i437_stall_in;
wire local_bb3__29_i437_inputs_ready;
wire local_bb3__29_i437_stall_local;
wire local_bb3__29_i437;

assign local_bb3__29_i437_inputs_ready = (rnode_339to340_bb3_shr_i404_0_valid_out_NO_SHIFT_REG & rnode_339to340_bb3_and6_i411_0_valid_out_2_NO_SHIFT_REG & rnode_339to340_bb3_shr2_i406_0_valid_out_NO_SHIFT_REG & rnode_339to340_bb3_and6_i411_0_valid_out_1_NO_SHIFT_REG & rnode_339to340_bb3_and6_i411_0_valid_out_0_NO_SHIFT_REG & rnode_339to340_bb3_and5_i410_0_valid_out_NO_SHIFT_REG);
assign local_bb3__29_i437 = (local_bb3__28_i436 | local_bb3__27_i434);
assign local_bb3_add_i449_valid_out = 1'b1;
assign local_bb3_reduction_0_i467_valid_out = 1'b1;
assign local_bb3_var__u45_valid_out = 1'b1;
assign local_bb3__29_i437_valid_out = 1'b1;
assign rnode_339to340_bb3_shr_i404_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_and6_i411_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_shr2_i406_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_and6_i411_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_and6_i411_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_339to340_bb3_and5_i410_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_340to342_bb3_add_i449_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_340to342_bb3_add_i449_0_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_340to342_bb3_add_i449_1_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_340to342_bb3_add_i449_2_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to342_bb3_add_i449_0_reg_342_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_valid_out_0_reg_342_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_stall_in_0_reg_342_NO_SHIFT_REG;
 logic rnode_340to342_bb3_add_i449_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_340to342_bb3_add_i449_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to342_bb3_add_i449_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to342_bb3_add_i449_0_stall_in_0_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_340to342_bb3_add_i449_0_valid_out_0_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_340to342_bb3_add_i449_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in((local_bb3_add_i449 & 32'h1FF)),
	.data_out(rnode_340to342_bb3_add_i449_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_340to342_bb3_add_i449_0_reg_342_fifo.DEPTH = 2;
defparam rnode_340to342_bb3_add_i449_0_reg_342_fifo.DATA_WIDTH = 32;
defparam rnode_340to342_bb3_add_i449_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to342_bb3_add_i449_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_340to342_bb3_add_i449_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add_i449_stall_in = 1'b0;
assign rnode_340to342_bb3_add_i449_0_stall_in_0_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_340to342_bb3_add_i449_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_340to342_bb3_add_i449_0_NO_SHIFT_REG = rnode_340to342_bb3_add_i449_0_reg_342_NO_SHIFT_REG;
assign rnode_340to342_bb3_add_i449_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_340to342_bb3_add_i449_1_NO_SHIFT_REG = rnode_340to342_bb3_add_i449_0_reg_342_NO_SHIFT_REG;
assign rnode_340to342_bb3_add_i449_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_340to342_bb3_add_i449_2_NO_SHIFT_REG = rnode_340to342_bb3_add_i449_0_reg_342_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb3_reduction_0_i467_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb3_reduction_0_i467_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb3_reduction_0_i467_0_NO_SHIFT_REG;
 logic rnode_340to341_bb3_reduction_0_i467_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb3_reduction_0_i467_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb3_reduction_0_i467_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb3_reduction_0_i467_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb3_reduction_0_i467_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb3_reduction_0_i467_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb3_reduction_0_i467_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb3_reduction_0_i467_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb3_reduction_0_i467_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb3_reduction_0_i467_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb3_reduction_0_i467),
	.data_out(rnode_340to341_bb3_reduction_0_i467_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb3_reduction_0_i467_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb3_reduction_0_i467_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb3_reduction_0_i467_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb3_reduction_0_i467_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb3_reduction_0_i467_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_reduction_0_i467_stall_in = 1'b0;
assign rnode_340to341_bb3_reduction_0_i467_0_NO_SHIFT_REG = rnode_340to341_bb3_reduction_0_i467_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb3_reduction_0_i467_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb3_reduction_0_i467_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_340to342_bb3_var__u45_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to342_bb3_var__u45_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to342_bb3_var__u45_0_NO_SHIFT_REG;
 logic rnode_340to342_bb3_var__u45_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to342_bb3_var__u45_0_reg_342_NO_SHIFT_REG;
 logic rnode_340to342_bb3_var__u45_0_valid_out_reg_342_NO_SHIFT_REG;
 logic rnode_340to342_bb3_var__u45_0_stall_in_reg_342_NO_SHIFT_REG;
 logic rnode_340to342_bb3_var__u45_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_340to342_bb3_var__u45_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to342_bb3_var__u45_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to342_bb3_var__u45_0_stall_in_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_340to342_bb3_var__u45_0_valid_out_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_340to342_bb3_var__u45_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in(local_bb3_var__u45),
	.data_out(rnode_340to342_bb3_var__u45_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_340to342_bb3_var__u45_0_reg_342_fifo.DEPTH = 2;
defparam rnode_340to342_bb3_var__u45_0_reg_342_fifo.DATA_WIDTH = 1;
defparam rnode_340to342_bb3_var__u45_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to342_bb3_var__u45_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_340to342_bb3_var__u45_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u45_stall_in = 1'b0;
assign rnode_340to342_bb3_var__u45_0_NO_SHIFT_REG = rnode_340to342_bb3_var__u45_0_reg_342_NO_SHIFT_REG;
assign rnode_340to342_bb3_var__u45_0_stall_in_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_340to342_bb3_var__u45_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb3__29_i437_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb3__29_i437_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb3__29_i437_0_NO_SHIFT_REG;
 logic rnode_340to341_bb3__29_i437_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb3__29_i437_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb3__29_i437_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb3__29_i437_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb3__29_i437_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb3__29_i437_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb3__29_i437_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb3__29_i437_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb3__29_i437_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb3__29_i437_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb3__29_i437),
	.data_out(rnode_340to341_bb3__29_i437_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb3__29_i437_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb3__29_i437_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb3__29_i437_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb3__29_i437_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb3__29_i437_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__29_i437_stall_in = 1'b0;
assign rnode_340to341_bb3__29_i437_0_NO_SHIFT_REG = rnode_340to341_bb3__29_i437_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb3__29_i437_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb3__29_i437_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_inc_i452_stall_local;
wire [31:0] local_bb3_inc_i452;

assign local_bb3_inc_i452 = ((rnode_340to342_bb3_add_i449_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp50_not_i457_stall_local;
wire local_bb3_cmp50_not_i457;

assign local_bb3_cmp50_not_i457 = ((rnode_340to342_bb3_add_i449_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_341to343_bb3_reduction_0_i467_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to343_bb3_reduction_0_i467_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to343_bb3_reduction_0_i467_0_NO_SHIFT_REG;
 logic rnode_341to343_bb3_reduction_0_i467_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to343_bb3_reduction_0_i467_0_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb3_reduction_0_i467_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb3_reduction_0_i467_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb3_reduction_0_i467_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_341to343_bb3_reduction_0_i467_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to343_bb3_reduction_0_i467_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to343_bb3_reduction_0_i467_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_341to343_bb3_reduction_0_i467_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_341to343_bb3_reduction_0_i467_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb3_reduction_0_i467_0_NO_SHIFT_REG),
	.data_out(rnode_341to343_bb3_reduction_0_i467_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_341to343_bb3_reduction_0_i467_0_reg_343_fifo.DEPTH = 2;
defparam rnode_341to343_bb3_reduction_0_i467_0_reg_343_fifo.DATA_WIDTH = 1;
defparam rnode_341to343_bb3_reduction_0_i467_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to343_bb3_reduction_0_i467_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_341to343_bb3_reduction_0_i467_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb3_reduction_0_i467_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to343_bb3_reduction_0_i467_0_NO_SHIFT_REG = rnode_341to343_bb3_reduction_0_i467_0_reg_343_NO_SHIFT_REG;
assign rnode_341to343_bb3_reduction_0_i467_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_341to343_bb3_reduction_0_i467_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_341to344_bb3__29_i437_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to344_bb3__29_i437_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to344_bb3__29_i437_0_NO_SHIFT_REG;
 logic rnode_341to344_bb3__29_i437_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to344_bb3__29_i437_0_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb3__29_i437_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb3__29_i437_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb3__29_i437_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_341to344_bb3__29_i437_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to344_bb3__29_i437_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to344_bb3__29_i437_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_341to344_bb3__29_i437_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_341to344_bb3__29_i437_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb3__29_i437_0_NO_SHIFT_REG),
	.data_out(rnode_341to344_bb3__29_i437_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_341to344_bb3__29_i437_0_reg_344_fifo.DEPTH = 3;
defparam rnode_341to344_bb3__29_i437_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_341to344_bb3__29_i437_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to344_bb3__29_i437_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_341to344_bb3__29_i437_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb3__29_i437_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb3__29_i437_0_NO_SHIFT_REG = rnode_341to344_bb3__29_i437_0_reg_344_NO_SHIFT_REG;
assign rnode_341to344_bb3__29_i437_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb3__29_i437_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__31_i458_stall_local;
wire local_bb3__31_i458;

assign local_bb3__31_i458 = (local_bb3_tobool49_i451 & local_bb3_cmp50_not_i457);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb3_reduction_0_i467_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to344_bb3_reduction_0_i467_0_stall_in_NO_SHIFT_REG;
 logic rnode_343to344_bb3_reduction_0_i467_0_NO_SHIFT_REG;
 logic rnode_343to344_bb3_reduction_0_i467_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to344_bb3_reduction_0_i467_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3_reduction_0_i467_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3_reduction_0_i467_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3_reduction_0_i467_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb3_reduction_0_i467_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb3_reduction_0_i467_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb3_reduction_0_i467_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb3_reduction_0_i467_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb3_reduction_0_i467_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(rnode_341to343_bb3_reduction_0_i467_0_NO_SHIFT_REG),
	.data_out(rnode_343to344_bb3_reduction_0_i467_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb3_reduction_0_i467_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb3_reduction_0_i467_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_343to344_bb3_reduction_0_i467_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb3_reduction_0_i467_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb3_reduction_0_i467_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to343_bb3_reduction_0_i467_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb3_reduction_0_i467_0_NO_SHIFT_REG = rnode_343to344_bb3_reduction_0_i467_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb3_reduction_0_i467_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb3_reduction_0_i467_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb3__29_i437_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb3__29_i437_0_stall_in_NO_SHIFT_REG;
 logic rnode_344to345_bb3__29_i437_0_NO_SHIFT_REG;
 logic rnode_344to345_bb3__29_i437_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_344to345_bb3__29_i437_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3__29_i437_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3__29_i437_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3__29_i437_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb3__29_i437_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb3__29_i437_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb3__29_i437_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb3__29_i437_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb3__29_i437_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(rnode_341to344_bb3__29_i437_0_NO_SHIFT_REG),
	.data_out(rnode_344to345_bb3__29_i437_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb3__29_i437_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb3__29_i437_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_344to345_bb3__29_i437_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb3__29_i437_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb3__29_i437_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to344_bb3__29_i437_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb3__29_i437_0_NO_SHIFT_REG = rnode_344to345_bb3__29_i437_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb3__29_i437_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb3__29_i437_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__32_i459_stall_local;
wire [31:0] local_bb3__32_i459;

assign local_bb3__32_i459 = (local_bb3__31_i458 ? (local_bb3_shl1_i_i456 & 32'hFFFFFE00) : (local_bb3_shl1_i18_i448 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__34_i461_stall_local;
wire [31:0] local_bb3__34_i461;

assign local_bb3__34_i461 = (local_bb3__31_i458 ? (local_bb3_or_i_i455 & 32'h1FFFFFF) : (local_bb3_or_i17_i447 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__36_i463_stall_local;
wire [31:0] local_bb3__36_i463;

assign local_bb3__36_i463 = (local_bb3__31_i458 ? (rnode_340to342_bb3_add_i449_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb3__33_i460_stall_local;
wire [31:0] local_bb3__33_i460;

assign local_bb3__33_i460 = (local_bb3_tobool49_i451 ? (local_bb3__32_i459 & 32'hFFFFFF00) : (local_bb3_shl1_i18_i448 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__35_i462_stall_local;
wire [31:0] local_bb3__35_i462;

assign local_bb3__35_i462 = (local_bb3_tobool49_i451 ? (local_bb3__34_i461 & 32'h1FFFFFF) : (local_bb3_or_i17_i447 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__37_i464_stall_local;
wire [31:0] local_bb3__37_i464;

assign local_bb3__37_i464 = (local_bb3_tobool49_i451 ? (local_bb3__36_i463 & 32'h1FF) : (local_bb3_inc_i452 & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb3_and75_i470_stall_local;
wire [31:0] local_bb3_and75_i470;

assign local_bb3_and75_i470 = ((local_bb3__35_i462 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and83_i476_stall_local;
wire [31:0] local_bb3_and83_i476;

assign local_bb3_and83_i476 = ((local_bb3__35_i462 & 32'h1FFFFFF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp53_i465_stall_local;
wire local_bb3_cmp53_i465;

assign local_bb3_cmp53_i465 = ((local_bb3__37_i464 & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp68_i469_stall_local;
wire local_bb3_cmp68_i469;

assign local_bb3_cmp68_i469 = ((local_bb3__37_i464 & 32'h3FF) < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb3_sub_i471_stall_local;
wire [31:0] local_bb3_sub_i471;

assign local_bb3_sub_i471 = ((local_bb3__37_i464 & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp71_not_i486_stall_local;
wire local_bb3_cmp71_not_i486;

assign local_bb3_cmp71_not_i486 = ((local_bb3__37_i464 & 32'h3FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb3_or581_i466_stall_local;
wire local_bb3_or581_i466;

assign local_bb3_or581_i466 = (rnode_340to342_bb3_var__u45_0_NO_SHIFT_REG | local_bb3_cmp53_i465);

// This section implements an unregistered operation.
// 
wire local_bb3_and74_i472_stall_local;
wire [31:0] local_bb3_and74_i472;

assign local_bb3_and74_i472 = ((local_bb3_sub_i471 & 32'hFF800000) + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb3__33_i460_valid_out;
wire local_bb3__33_i460_stall_in;
wire local_bb3_cmp68_i469_valid_out;
wire local_bb3_cmp68_i469_stall_in;
wire local_bb3_cmp71_not_i486_valid_out;
wire local_bb3_cmp71_not_i486_stall_in;
wire local_bb3_or581_i466_valid_out;
wire local_bb3_or581_i466_stall_in;
wire local_bb3_and75_i470_valid_out;
wire local_bb3_and75_i470_stall_in;
wire local_bb3_and83_i476_valid_out;
wire local_bb3_and83_i476_stall_in;
wire local_bb3_shl_i473_valid_out;
wire local_bb3_shl_i473_stall_in;
wire local_bb3_shl_i473_inputs_ready;
wire local_bb3_shl_i473_stall_local;
wire [31:0] local_bb3_shl_i473;

assign local_bb3_shl_i473_inputs_ready = (local_bb3_mul_i_i442_valid_out_0_NO_SHIFT_REG & rnode_340to342_bb3_add_i449_0_valid_out_1_NO_SHIFT_REG & rnode_340to342_bb3_add_i449_0_valid_out_0_NO_SHIFT_REG & rnode_340to342_bb3_add_i449_0_valid_out_2_NO_SHIFT_REG & local_bb3_mul_i_i442_valid_out_1_NO_SHIFT_REG & rnode_340to342_bb3_var__u45_0_valid_out_NO_SHIFT_REG);
assign local_bb3_shl_i473 = ((local_bb3_and74_i472 & 32'hFF800000) & 32'h7F800000);
assign local_bb3__33_i460_valid_out = 1'b1;
assign local_bb3_cmp68_i469_valid_out = 1'b1;
assign local_bb3_cmp71_not_i486_valid_out = 1'b1;
assign local_bb3_or581_i466_valid_out = 1'b1;
assign local_bb3_and75_i470_valid_out = 1'b1;
assign local_bb3_and83_i476_valid_out = 1'b1;
assign local_bb3_shl_i473_valid_out = 1'b1;
assign local_bb3_mul_i_i442_stall_in_0 = 1'b0;
assign rnode_340to342_bb3_add_i449_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_340to342_bb3_add_i449_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_340to342_bb3_add_i449_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign local_bb3_mul_i_i442_stall_in_1 = 1'b0;
assign rnode_340to342_bb3_var__u45_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb3__33_i460_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_342to343_bb3__33_i460_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3__33_i460_0_NO_SHIFT_REG;
 logic rnode_342to343_bb3__33_i460_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_342to343_bb3__33_i460_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3__33_i460_1_NO_SHIFT_REG;
 logic rnode_342to343_bb3__33_i460_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3__33_i460_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3__33_i460_0_valid_out_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3__33_i460_0_stall_in_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3__33_i460_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb3__33_i460_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb3__33_i460_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb3__33_i460_0_stall_in_0_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb3__33_i460_0_valid_out_0_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb3__33_i460_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb3__33_i460 & 32'hFFFFFF00)),
	.data_out(rnode_342to343_bb3__33_i460_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb3__33_i460_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb3__33_i460_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb3__33_i460_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb3__33_i460_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb3__33_i460_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__33_i460_stall_in = 1'b0;
assign rnode_342to343_bb3__33_i460_0_stall_in_0_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb3__33_i460_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb3__33_i460_0_NO_SHIFT_REG = rnode_342to343_bb3__33_i460_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb3__33_i460_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb3__33_i460_1_NO_SHIFT_REG = rnode_342to343_bb3__33_i460_0_reg_343_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_342to344_bb3_cmp68_i469_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp68_i469_0_stall_in_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp68_i469_0_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp68_i469_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp68_i469_0_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp68_i469_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp68_i469_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp68_i469_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_342to344_bb3_cmp68_i469_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to344_bb3_cmp68_i469_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to344_bb3_cmp68_i469_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_342to344_bb3_cmp68_i469_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_342to344_bb3_cmp68_i469_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(local_bb3_cmp68_i469),
	.data_out(rnode_342to344_bb3_cmp68_i469_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_342to344_bb3_cmp68_i469_0_reg_344_fifo.DEPTH = 2;
defparam rnode_342to344_bb3_cmp68_i469_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_342to344_bb3_cmp68_i469_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to344_bb3_cmp68_i469_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_342to344_bb3_cmp68_i469_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp68_i469_stall_in = 1'b0;
assign rnode_342to344_bb3_cmp68_i469_0_NO_SHIFT_REG = rnode_342to344_bb3_cmp68_i469_0_reg_344_NO_SHIFT_REG;
assign rnode_342to344_bb3_cmp68_i469_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_342to344_bb3_cmp68_i469_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_342to344_bb3_cmp71_not_i486_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp71_not_i486_0_stall_in_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp71_not_i486_0_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp71_not_i486_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp71_not_i486_0_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp71_not_i486_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp71_not_i486_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_cmp71_not_i486_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_342to344_bb3_cmp71_not_i486_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to344_bb3_cmp71_not_i486_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to344_bb3_cmp71_not_i486_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_342to344_bb3_cmp71_not_i486_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_342to344_bb3_cmp71_not_i486_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(local_bb3_cmp71_not_i486),
	.data_out(rnode_342to344_bb3_cmp71_not_i486_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_342to344_bb3_cmp71_not_i486_0_reg_344_fifo.DEPTH = 2;
defparam rnode_342to344_bb3_cmp71_not_i486_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_342to344_bb3_cmp71_not_i486_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to344_bb3_cmp71_not_i486_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_342to344_bb3_cmp71_not_i486_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp71_not_i486_stall_in = 1'b0;
assign rnode_342to344_bb3_cmp71_not_i486_0_NO_SHIFT_REG = rnode_342to344_bb3_cmp71_not_i486_0_reg_344_NO_SHIFT_REG;
assign rnode_342to344_bb3_cmp71_not_i486_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_342to344_bb3_cmp71_not_i486_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_342to344_bb3_or581_i466_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_1_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_valid_out_0_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_stall_in_0_reg_344_NO_SHIFT_REG;
 logic rnode_342to344_bb3_or581_i466_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_342to344_bb3_or581_i466_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to344_bb3_or581_i466_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to344_bb3_or581_i466_0_stall_in_0_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_342to344_bb3_or581_i466_0_valid_out_0_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_342to344_bb3_or581_i466_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(local_bb3_or581_i466),
	.data_out(rnode_342to344_bb3_or581_i466_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_342to344_bb3_or581_i466_0_reg_344_fifo.DEPTH = 2;
defparam rnode_342to344_bb3_or581_i466_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_342to344_bb3_or581_i466_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to344_bb3_or581_i466_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_342to344_bb3_or581_i466_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or581_i466_stall_in = 1'b0;
assign rnode_342to344_bb3_or581_i466_0_stall_in_0_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_342to344_bb3_or581_i466_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_342to344_bb3_or581_i466_0_NO_SHIFT_REG = rnode_342to344_bb3_or581_i466_0_reg_344_NO_SHIFT_REG;
assign rnode_342to344_bb3_or581_i466_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_342to344_bb3_or581_i466_1_NO_SHIFT_REG = rnode_342to344_bb3_or581_i466_0_reg_344_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb3_and75_i470_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and75_i470_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3_and75_i470_0_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and75_i470_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3_and75_i470_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and75_i470_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and75_i470_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and75_i470_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb3_and75_i470_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb3_and75_i470_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb3_and75_i470_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb3_and75_i470_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb3_and75_i470_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb3_and75_i470 & 32'h7FFFFF)),
	.data_out(rnode_342to343_bb3_and75_i470_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb3_and75_i470_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb3_and75_i470_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb3_and75_i470_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb3_and75_i470_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb3_and75_i470_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and75_i470_stall_in = 1'b0;
assign rnode_342to343_bb3_and75_i470_0_NO_SHIFT_REG = rnode_342to343_bb3_and75_i470_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb3_and75_i470_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb3_and75_i470_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb3_and83_i476_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and83_i476_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3_and83_i476_0_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and83_i476_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3_and83_i476_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and83_i476_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and83_i476_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_and83_i476_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb3_and83_i476_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb3_and83_i476_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb3_and83_i476_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb3_and83_i476_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb3_and83_i476_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb3_and83_i476 & 32'h1)),
	.data_out(rnode_342to343_bb3_and83_i476_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb3_and83_i476_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb3_and83_i476_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb3_and83_i476_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb3_and83_i476_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb3_and83_i476_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and83_i476_stall_in = 1'b0;
assign rnode_342to343_bb3_and83_i476_0_NO_SHIFT_REG = rnode_342to343_bb3_and83_i476_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb3_and83_i476_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb3_and83_i476_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb3_shl_i473_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb3_shl_i473_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3_shl_i473_0_NO_SHIFT_REG;
 logic rnode_342to343_bb3_shl_i473_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb3_shl_i473_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_shl_i473_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_shl_i473_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb3_shl_i473_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb3_shl_i473_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb3_shl_i473_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb3_shl_i473_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb3_shl_i473_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb3_shl_i473_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb3_shl_i473 & 32'h7F800000)),
	.data_out(rnode_342to343_bb3_shl_i473_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb3_shl_i473_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb3_shl_i473_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb3_shl_i473_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb3_shl_i473_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb3_shl_i473_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shl_i473_stall_in = 1'b0;
assign rnode_342to343_bb3_shl_i473_0_NO_SHIFT_REG = rnode_342to343_bb3_shl_i473_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb3_shl_i473_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb3_shl_i473_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp77_i475_stall_local;
wire local_bb3_cmp77_i475;

assign local_bb3_cmp77_i475 = ((rnode_342to343_bb3__33_i460_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u47_stall_local;
wire local_bb3_var__u47;

assign local_bb3_var__u47 = ($signed((rnode_342to343_bb3__33_i460_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u48_stall_local;
wire [31:0] local_bb3_var__u48;

assign local_bb3_var__u48[31:1] = 31'h0;
assign local_bb3_var__u48[0] = rnode_342to344_bb3_cmp68_i469_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_2_i468_stall_local;
wire local_bb3_reduction_2_i468;

assign local_bb3_reduction_2_i468 = (rnode_343to344_bb3_reduction_0_i467_0_NO_SHIFT_REG | rnode_342to344_bb3_or581_i466_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb3_or581_i466_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb3_or581_i466_0_stall_in_NO_SHIFT_REG;
 logic rnode_344to345_bb3_or581_i466_0_NO_SHIFT_REG;
 logic rnode_344to345_bb3_or581_i466_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_344to345_bb3_or581_i466_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3_or581_i466_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3_or581_i466_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3_or581_i466_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb3_or581_i466_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb3_or581_i466_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb3_or581_i466_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb3_or581_i466_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb3_or581_i466_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(rnode_342to344_bb3_or581_i466_1_NO_SHIFT_REG),
	.data_out(rnode_344to345_bb3_or581_i466_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb3_or581_i466_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb3_or581_i466_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_344to345_bb3_or581_i466_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb3_or581_i466_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb3_or581_i466_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_342to344_bb3_or581_i466_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb3_or581_i466_0_NO_SHIFT_REG = rnode_344to345_bb3_or581_i466_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb3_or581_i466_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb3_or581_i466_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_tobool84_i477_stall_local;
wire local_bb3_tobool84_i477;

assign local_bb3_tobool84_i477 = ((rnode_342to343_bb3_and83_i476_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or76_i474_valid_out;
wire local_bb3_or76_i474_stall_in;
wire local_bb3_or76_i474_inputs_ready;
wire local_bb3_or76_i474_stall_local;
wire [31:0] local_bb3_or76_i474;

assign local_bb3_or76_i474_inputs_ready = (rnode_342to343_bb3_shl_i473_0_valid_out_NO_SHIFT_REG & rnode_342to343_bb3_and75_i470_0_valid_out_NO_SHIFT_REG);
assign local_bb3_or76_i474 = ((rnode_342to343_bb3_shl_i473_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_342to343_bb3_and75_i470_0_NO_SHIFT_REG & 32'h7FFFFF));
assign local_bb3_or76_i474_valid_out = 1'b1;
assign rnode_342to343_bb3_shl_i473_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb3_and75_i470_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_conv101_i489_stall_local;
wire [31:0] local_bb3_conv101_i489;

assign local_bb3_conv101_i489[31:1] = 31'h0;
assign local_bb3_conv101_i489[0] = local_bb3_reduction_2_i468;

// This section implements an unregistered operation.
// 
wire local_bb3_cond111_i494_stall_local;
wire [31:0] local_bb3_cond111_i494;

assign local_bb3_cond111_i494 = (rnode_344to345_bb3_or581_i466_0_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__39_i478_stall_local;
wire local_bb3__39_i478;

assign local_bb3__39_i478 = (local_bb3_tobool84_i477 & local_bb3_var__u47);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb3_or76_i474_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to344_bb3_or76_i474_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb3_or76_i474_0_NO_SHIFT_REG;
 logic rnode_343to344_bb3_or76_i474_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb3_or76_i474_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3_or76_i474_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3_or76_i474_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3_or76_i474_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb3_or76_i474_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb3_or76_i474_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb3_or76_i474_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb3_or76_i474_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb3_or76_i474_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in((local_bb3_or76_i474 & 32'h7FFFFFFF)),
	.data_out(rnode_343to344_bb3_or76_i474_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb3_or76_i474_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb3_or76_i474_0_reg_344_fifo.DATA_WIDTH = 32;
defparam rnode_343to344_bb3_or76_i474_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb3_or76_i474_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb3_or76_i474_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or76_i474_stall_in = 1'b0;
assign rnode_343to344_bb3_or76_i474_0_NO_SHIFT_REG = rnode_343to344_bb3_or76_i474_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb3_or76_i474_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb3_or76_i474_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__40_i479_valid_out;
wire local_bb3__40_i479_stall_in;
wire local_bb3__40_i479_inputs_ready;
wire local_bb3__40_i479_stall_local;
wire local_bb3__40_i479;

assign local_bb3__40_i479_inputs_ready = (rnode_342to343_bb3__33_i460_0_valid_out_0_NO_SHIFT_REG & rnode_342to343_bb3__33_i460_0_valid_out_1_NO_SHIFT_REG & rnode_342to343_bb3_and83_i476_0_valid_out_NO_SHIFT_REG);
assign local_bb3__40_i479 = (local_bb3_cmp77_i475 | local_bb3__39_i478);
assign local_bb3__40_i479_valid_out = 1'b1;
assign rnode_342to343_bb3__33_i460_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb3__33_i460_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb3_and83_i476_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb3__40_i479_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to344_bb3__40_i479_0_stall_in_NO_SHIFT_REG;
 logic rnode_343to344_bb3__40_i479_0_NO_SHIFT_REG;
 logic rnode_343to344_bb3__40_i479_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to344_bb3__40_i479_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3__40_i479_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3__40_i479_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb3__40_i479_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb3__40_i479_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb3__40_i479_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb3__40_i479_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb3__40_i479_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb3__40_i479_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(local_bb3__40_i479),
	.data_out(rnode_343to344_bb3__40_i479_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb3__40_i479_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb3__40_i479_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_343to344_bb3__40_i479_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb3__40_i479_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb3__40_i479_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__40_i479_stall_in = 1'b0;
assign rnode_343to344_bb3__40_i479_0_NO_SHIFT_REG = rnode_343to344_bb3__40_i479_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb3__40_i479_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb3__40_i479_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cond_i480_stall_local;
wire [31:0] local_bb3_cond_i480;

assign local_bb3_cond_i480[31:1] = 31'h0;
assign local_bb3_cond_i480[0] = rnode_343to344_bb3__40_i479_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_add87_i481_stall_local;
wire [31:0] local_bb3_add87_i481;

assign local_bb3_add87_i481 = ((local_bb3_cond_i480 & 32'h1) + (rnode_343to344_bb3_or76_i474_0_NO_SHIFT_REG & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_and90_i484_stall_local;
wire [31:0] local_bb3_and90_i484;

assign local_bb3_and90_i484 = (local_bb3_add87_i481 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp91_i485_stall_local;
wire local_bb3_cmp91_i485;

assign local_bb3_cmp91_i485 = ((local_bb3_and90_i484 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge14_i487_stall_local;
wire local_bb3_brmerge14_i487;

assign local_bb3_brmerge14_i487 = (local_bb3_cmp91_i485 | rnode_342to344_bb3_cmp71_not_i486_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_conv99_i488_stall_local;
wire [31:0] local_bb3_conv99_i488;

assign local_bb3_conv99_i488 = (local_bb3_brmerge14_i487 ? (local_bb3_var__u48 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or102_i490_stall_local;
wire [31:0] local_bb3_or102_i490;

assign local_bb3_or102_i490 = ((local_bb3_conv99_i488 & 32'h1) | (local_bb3_conv101_i489 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_sext_stall_local;
wire [31:0] local_bb3_sext;

assign local_bb3_sext = ((local_bb3_or102_i490 & 32'h1) + 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and108_i493_valid_out;
wire local_bb3_and108_i493_stall_in;
wire local_bb3_and108_i493_inputs_ready;
wire local_bb3_and108_i493_stall_local;
wire [31:0] local_bb3_and108_i493;

assign local_bb3_and108_i493_inputs_ready = (rnode_342to344_bb3_or581_i466_0_valid_out_0_NO_SHIFT_REG & rnode_343to344_bb3_reduction_0_i467_0_valid_out_NO_SHIFT_REG & rnode_342to344_bb3_cmp68_i469_0_valid_out_NO_SHIFT_REG & rnode_342to344_bb3_cmp71_not_i486_0_valid_out_NO_SHIFT_REG & rnode_343to344_bb3__40_i479_0_valid_out_NO_SHIFT_REG & rnode_343to344_bb3_or76_i474_0_valid_out_NO_SHIFT_REG);
assign local_bb3_and108_i493 = (local_bb3_sext & local_bb3_add87_i481);
assign local_bb3_and108_i493_valid_out = 1'b1;
assign rnode_342to344_bb3_or581_i466_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb3_reduction_0_i467_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_342to344_bb3_cmp68_i469_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_342to344_bb3_cmp71_not_i486_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb3__40_i479_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb3_or76_i474_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb3_and108_i493_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb3_and108_i493_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb3_and108_i493_0_NO_SHIFT_REG;
 logic rnode_344to345_bb3_and108_i493_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb3_and108_i493_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3_and108_i493_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3_and108_i493_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb3_and108_i493_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb3_and108_i493_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb3_and108_i493_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb3_and108_i493_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb3_and108_i493_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb3_and108_i493_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(local_bb3_and108_i493),
	.data_out(rnode_344to345_bb3_and108_i493_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb3_and108_i493_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb3_and108_i493_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_344to345_bb3_and108_i493_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb3_and108_i493_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb3_and108_i493_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and108_i493_stall_in = 1'b0;
assign rnode_344to345_bb3_and108_i493_0_NO_SHIFT_REG = rnode_344to345_bb3_and108_i493_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb3_and108_i493_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb3_and108_i493_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_or112_i495_stall_local;
wire [31:0] local_bb3_or112_i495;

assign local_bb3_or112_i495 = (rnode_344to345_bb3_and108_i493_0_NO_SHIFT_REG | (local_bb3_cond111_i494 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb3_or112_i495_op_stall_local;
wire [31:0] local_bb3_or112_i495_op;

assign local_bb3_or112_i495_op = (local_bb3_or112_i495 | 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u49_stall_local;
wire [31:0] local_bb3_var__u49;

assign local_bb3_var__u49 = (local_bb3_or112_i495_op | 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_cast_after_negation_valid_out;
wire local_bb3_cast_after_negation_stall_in;
wire local_bb3_cast_after_negation_inputs_ready;
wire local_bb3_cast_after_negation_stall_local;
wire [31:0] local_bb3_cast_after_negation;

assign local_bb3_cast_after_negation_inputs_ready = (rnode_344to345_bb3__29_i437_0_valid_out_NO_SHIFT_REG & rnode_344to345_bb3_or581_i466_0_valid_out_NO_SHIFT_REG & rnode_344to345_bb3_and108_i493_0_valid_out_NO_SHIFT_REG);
assign local_bb3_cast_after_negation = (rnode_344to345_bb3__29_i437_0_NO_SHIFT_REG ? 32'hFFC00000 : local_bb3_var__u49);
assign local_bb3_cast_after_negation_valid_out = 1'b1;
assign rnode_344to345_bb3__29_i437_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb3_or581_i466_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb3_and108_i493_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb3_div_inputs_ready;
 reg local_bb3_div_valid_out_NO_SHIFT_REG;
wire local_bb3_div_stall_in;
wire local_bb3_div_output_regs_ready;
wire [31:0] local_bb3_div;
 reg local_bb3_div_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb3_div_valid_pipe_12_NO_SHIFT_REG;
wire local_bb3_div_causedstall;

acl_fp_div_s5 fp_module_local_bb3_div (
	.clock(clock),
	.dataa(local_bb3_cast_after_negation),
	.datab(input_wii_mul50),
	.enable(local_bb3_div_output_regs_ready),
	.result(local_bb3_div)
);


assign local_bb3_div_inputs_ready = 1'b1;
assign local_bb3_div_output_regs_ready = 1'b1;
assign local_bb3_cast_after_negation_stall_in = 1'b0;
assign local_bb3_div_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_div_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb3_div_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_div_output_regs_ready)
		begin
			local_bb3_div_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_div_valid_pipe_1_NO_SHIFT_REG <= local_bb3_div_valid_pipe_0_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_2_NO_SHIFT_REG <= local_bb3_div_valid_pipe_1_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_3_NO_SHIFT_REG <= local_bb3_div_valid_pipe_2_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_4_NO_SHIFT_REG <= local_bb3_div_valid_pipe_3_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_5_NO_SHIFT_REG <= local_bb3_div_valid_pipe_4_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_6_NO_SHIFT_REG <= local_bb3_div_valid_pipe_5_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_7_NO_SHIFT_REG <= local_bb3_div_valid_pipe_6_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_8_NO_SHIFT_REG <= local_bb3_div_valid_pipe_7_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_9_NO_SHIFT_REG <= local_bb3_div_valid_pipe_8_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_10_NO_SHIFT_REG <= local_bb3_div_valid_pipe_9_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_11_NO_SHIFT_REG <= local_bb3_div_valid_pipe_10_NO_SHIFT_REG;
			local_bb3_div_valid_pipe_12_NO_SHIFT_REG <= local_bb3_div_valid_pipe_11_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_div_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_div_output_regs_ready)
		begin
			local_bb3_div_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_div_stall_in))
			begin
				local_bb3_div_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_call_i_div_inputs_ready;
 reg local_bb3_call_i_div_valid_out_0_NO_SHIFT_REG;
wire local_bb3_call_i_div_stall_in_0;
 reg local_bb3_call_i_div_valid_out_1_NO_SHIFT_REG;
wire local_bb3_call_i_div_stall_in_1;
wire local_bb3_call_i_div_output_regs_ready;
wire [31:0] local_bb3_call_i_div;
 reg local_bb3_call_i_div_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_12_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_13_NO_SHIFT_REG;
 reg local_bb3_call_i_div_valid_pipe_14_NO_SHIFT_REG;
wire local_bb3_call_i_div_causedstall;

acl_fp_exp_s5 fp_module_local_bb3_call_i_div (
	.clock(clock),
	.dataa(local_bb3_div),
	.enable(local_bb3_call_i_div_output_regs_ready),
	.result(local_bb3_call_i_div)
);


assign local_bb3_call_i_div_inputs_ready = 1'b1;
assign local_bb3_call_i_div_output_regs_ready = 1'b1;
assign local_bb3_div_stall_in = 1'b0;
assign local_bb3_call_i_div_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_call_i_div_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_13_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_pipe_14_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_call_i_div_output_regs_ready)
		begin
			local_bb3_call_i_div_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_call_i_div_valid_pipe_1_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_0_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_2_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_1_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_3_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_2_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_4_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_3_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_5_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_4_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_6_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_5_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_7_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_6_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_8_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_7_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_9_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_8_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_10_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_9_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_11_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_10_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_12_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_11_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_13_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_12_NO_SHIFT_REG;
			local_bb3_call_i_div_valid_pipe_14_NO_SHIFT_REG <= local_bb3_call_i_div_valid_pipe_13_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_call_i_div_output_regs_ready)
		begin
			local_bb3_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_call_i_div_stall_in_0))
			begin
				local_bb3_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_call_i_div_stall_in_1))
			begin
				local_bb3_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_astype_i_i_stall_local;
wire [31:0] local_bb3_astype_i_i;

assign local_bb3_astype_i_i = local_bb3_call_i_div;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u50_stall_local;
wire [31:0] local_bb3_var__u50;

assign local_bb3_var__u50 = local_bb3_call_i_div;

// This section implements an unregistered operation.
// 
wire local_bb3_and_i_i_stall_local;
wire [31:0] local_bb3_and_i_i;

assign local_bb3_and_i_i = (local_bb3_astype_i_i & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i_i_stall_local;
wire local_bb3_cmp_i_i;

assign local_bb3_cmp_i_i = ((local_bb3_and_i_i & 32'h7F800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u51_stall_local;
wire [31:0] local_bb3_var__u51;

assign local_bb3_var__u51 = (local_bb3_cmp_i_i ? 32'h0 : local_bb3_var__u50);

// This section implements an unregistered operation.
// 
wire local_bb3_shr2_i222_stall_local;
wire [31:0] local_bb3_shr2_i222;

assign local_bb3_shr2_i222 = (local_bb3_var__u51 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_xor_i224_stall_local;
wire [31:0] local_bb3_xor_i224;

assign local_bb3_xor_i224 = (local_bb3_var__u51 ^ rnode_374to375_bb3_var__u37_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_and6_i227_stall_local;
wire [31:0] local_bb3_and6_i227;

assign local_bb3_and6_i227 = (local_bb3_var__u51 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and3_i223_stall_local;
wire [31:0] local_bb3_and3_i223;

assign local_bb3_and3_i223 = ((local_bb3_shr2_i222 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_i233_stall_local;
wire local_bb3_lnot17_i233;

assign local_bb3_lnot17_i233 = ((local_bb3_and6_i227 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u52_stall_local;
wire [31:0] local_bb3_var__u52;

assign local_bb3_var__u52 = ((local_bb3_and6_i227 & 32'h7FFFFF) | (local_bb3_and_i221 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_or47_i255_stall_local;
wire [31:0] local_bb3_or47_i255;

assign local_bb3_or47_i255 = ((local_bb3_and6_i227 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot8_i229_stall_local;
wire local_bb3_lnot8_i229;

assign local_bb3_lnot8_i229 = ((local_bb3_and3_i223 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_i231_stall_local;
wire local_bb3_cmp11_i231;

assign local_bb3_cmp11_i231 = ((local_bb3_and3_i223 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u53_stall_local;
wire [31:0] local_bb3_var__u53;

assign local_bb3_var__u53 = ((local_bb3_and3_i223 & 32'hFF) | (local_bb3_and6_i227 & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_add_i265_stall_local;
wire [31:0] local_bb3_add_i265;

assign local_bb3_add_i265 = ((local_bb3_and3_i223 & 32'hFF) + (local_bb3_and_i221 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_not_i237_stall_local;
wire local_bb3_lnot17_not_i237;

assign local_bb3_lnot17_not_i237 = (local_bb3_lnot17_i233 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u54_stall_local;
wire local_bb3_var__u54;

assign local_bb3_var__u54 = ((local_bb3_var__u52 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_conv1_i_i257_stall_local;
wire [63:0] local_bb3_conv1_i_i257;

assign local_bb3_conv1_i_i257[63:32] = 32'h0;
assign local_bb3_conv1_i_i257[31:0] = ((local_bb3_or47_i255 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_0_i283_stall_local;
wire local_bb3_reduction_0_i283;

assign local_bb3_reduction_0_i283 = (local_bb3_lnot_i228 | local_bb3_lnot8_i229);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge8_demorgan_i234_stall_local;
wire local_bb3_brmerge8_demorgan_i234;

assign local_bb3_brmerge8_demorgan_i234 = (local_bb3_cmp11_i231 & local_bb3_lnot17_i233);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_not_i238_stall_local;
wire local_bb3_cmp11_not_i238;

assign local_bb3_cmp11_not_i238 = (local_bb3_cmp11_i231 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u55_stall_local;
wire local_bb3_var__u55;

assign local_bb3_var__u55 = ((local_bb3_var__u53 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge10_demorgan_i235_stall_local;
wire local_bb3_brmerge10_demorgan_i235;

assign local_bb3_brmerge10_demorgan_i235 = (local_bb3_brmerge8_demorgan_i234 & local_bb3_lnot_i228);

// This section implements an unregistered operation.
// 
wire local_bb3__mux9_mux_i236_stall_local;
wire local_bb3__mux9_mux_i236;

assign local_bb3__mux9_mux_i236 = (local_bb3_brmerge8_demorgan_i234 ^ local_bb3_cmp11_i231);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge3_i239_stall_local;
wire local_bb3_brmerge3_i239;

assign local_bb3_brmerge3_i239 = (local_bb3_var__u55 | local_bb3_cmp11_not_i238);

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_i241_stall_local;
wire local_bb3__mux_mux_i241;

assign local_bb3__mux_mux_i241 = (local_bb3_var__u55 | local_bb3_cmp11_i231);

// This section implements an unregistered operation.
// 
wire local_bb3__not_i243_stall_local;
wire local_bb3__not_i243;

assign local_bb3__not_i243 = (local_bb3_var__u55 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge5_i240_stall_local;
wire local_bb3_brmerge5_i240;

assign local_bb3_brmerge5_i240 = (local_bb3_brmerge3_i239 | local_bb3_lnot17_not_i237);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_3_i244_stall_local;
wire local_bb3_reduction_3_i244;

assign local_bb3_reduction_3_i244 = (local_bb3_cmp11_i231 & local_bb3__not_i243);

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_mux_i242_stall_local;
wire local_bb3__mux_mux_mux_i242;

assign local_bb3__mux_mux_mux_i242 = (local_bb3_brmerge5_i240 & local_bb3__mux_mux_i241);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_5_i245_stall_local;
wire local_bb3_reduction_5_i245;

assign local_bb3_reduction_5_i245 = (local_bb3_lnot14_i232 & local_bb3_reduction_3_i244);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i230_valid_out;
wire local_bb3_cmp_i230_stall_in;
wire local_bb3_add_i265_valid_out;
wire local_bb3_add_i265_stall_in;
wire local_bb3_brmerge10_demorgan_i235_valid_out;
wire local_bb3_brmerge10_demorgan_i235_stall_in;
wire local_bb3_reduction_0_i283_valid_out;
wire local_bb3_reduction_0_i283_stall_in;
wire local_bb3_lnot14_i232_valid_out_1;
wire local_bb3_lnot14_i232_stall_in_1;
wire local_bb3_conv_i_i256_valid_out;
wire local_bb3_conv_i_i256_stall_in;
wire local_bb3_reduction_6_i246_valid_out;
wire local_bb3_reduction_6_i246_stall_in;
wire local_bb3_xor_i224_valid_out;
wire local_bb3_xor_i224_stall_in;
wire local_bb3_cmp11_i231_valid_out_5;
wire local_bb3_cmp11_i231_stall_in_5;
wire local_bb3_conv1_i_i257_valid_out;
wire local_bb3_conv1_i_i257_stall_in;
wire local_bb3__mux9_mux_i236_valid_out;
wire local_bb3__mux9_mux_i236_stall_in;
wire local_bb3__mux_mux_mux_i242_valid_out;
wire local_bb3__mux_mux_mux_i242_stall_in;
wire local_bb3_reduction_6_i246_inputs_ready;
wire local_bb3_reduction_6_i246_stall_local;
wire local_bb3_reduction_6_i246;

assign local_bb3_reduction_6_i246_inputs_ready = (rnode_374to375_bb3_var__u37_0_valid_out_0_NO_SHIFT_REG & rnode_374to375_bb3_var__u37_0_valid_out_2_NO_SHIFT_REG & rnode_374to375_bb3_var__u37_0_valid_out_1_NO_SHIFT_REG & local_bb3_call_i_div_valid_out_1_NO_SHIFT_REG & local_bb3_call_i_div_valid_out_0_NO_SHIFT_REG);
assign local_bb3_reduction_6_i246 = (local_bb3_var__u54 & local_bb3_reduction_5_i245);
assign local_bb3_cmp_i230_valid_out = 1'b1;
assign local_bb3_add_i265_valid_out = 1'b1;
assign local_bb3_brmerge10_demorgan_i235_valid_out = 1'b1;
assign local_bb3_reduction_0_i283_valid_out = 1'b1;
assign local_bb3_lnot14_i232_valid_out_1 = 1'b1;
assign local_bb3_conv_i_i256_valid_out = 1'b1;
assign local_bb3_reduction_6_i246_valid_out = 1'b1;
assign local_bb3_xor_i224_valid_out = 1'b1;
assign local_bb3_cmp11_i231_valid_out_5 = 1'b1;
assign local_bb3_conv1_i_i257_valid_out = 1'b1;
assign local_bb3__mux9_mux_i236_valid_out = 1'b1;
assign local_bb3__mux_mux_mux_i242_valid_out = 1'b1;
assign rnode_374to375_bb3_var__u37_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_374to375_bb3_var__u37_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_374to375_bb3_var__u37_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign local_bb3_call_i_div_stall_in_1 = 1'b0;
assign local_bb3_call_i_div_stall_in_0 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_cmp_i230_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_2_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_3_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_valid_out_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_stall_in_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp_i230_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_cmp_i230_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_cmp_i230_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_cmp_i230_0_stall_in_0_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_cmp_i230_0_valid_out_0_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_cmp_i230_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3_cmp_i230),
	.data_out(rnode_375to376_bb3_cmp_i230_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_cmp_i230_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_cmp_i230_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3_cmp_i230_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_cmp_i230_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_cmp_i230_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp_i230_stall_in = 1'b0;
assign rnode_375to376_bb3_cmp_i230_0_stall_in_0_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_cmp_i230_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_cmp_i230_0_NO_SHIFT_REG = rnode_375to376_bb3_cmp_i230_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_cmp_i230_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_cmp_i230_1_NO_SHIFT_REG = rnode_375to376_bb3_cmp_i230_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_cmp_i230_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_cmp_i230_2_NO_SHIFT_REG = rnode_375to376_bb3_cmp_i230_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_cmp_i230_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_cmp_i230_3_NO_SHIFT_REG = rnode_375to376_bb3_cmp_i230_0_reg_376_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_add_i265_0_valid_out_NO_SHIFT_REG;
 logic rnode_375to376_bb3_add_i265_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_375to376_bb3_add_i265_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_add_i265_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_375to376_bb3_add_i265_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_add_i265_0_valid_out_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_add_i265_0_stall_in_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_add_i265_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_add_i265_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_add_i265_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_add_i265_0_stall_in_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_add_i265_0_valid_out_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_add_i265_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in((local_bb3_add_i265 & 32'h1FF)),
	.data_out(rnode_375to376_bb3_add_i265_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_add_i265_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_add_i265_0_reg_376_fifo.DATA_WIDTH = 32;
defparam rnode_375to376_bb3_add_i265_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_add_i265_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_add_i265_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add_i265_stall_in = 1'b0;
assign rnode_375to376_bb3_add_i265_0_NO_SHIFT_REG = rnode_375to376_bb3_add_i265_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_add_i265_0_stall_in_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_add_i265_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_in_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_in_0_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_0_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3_brmerge10_demorgan_i235),
	.data_out(rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_brmerge10_demorgan_i235_stall_in = 1'b0;
assign rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_in_0_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_brmerge10_demorgan_i235_0_NO_SHIFT_REG = rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_brmerge10_demorgan_i235_1_NO_SHIFT_REG = rnode_375to376_bb3_brmerge10_demorgan_i235_0_reg_376_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_0_i283_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_0_i283_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_0_i283_0_valid_out_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_0_i283_0_stall_in_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_0_i283_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_reduction_0_i283_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_reduction_0_i283_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_reduction_0_i283_0_stall_in_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_reduction_0_i283_0_valid_out_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_reduction_0_i283_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3_reduction_0_i283),
	.data_out(rnode_375to376_bb3_reduction_0_i283_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_reduction_0_i283_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_reduction_0_i283_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3_reduction_0_i283_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_reduction_0_i283_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_reduction_0_i283_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_reduction_0_i283_stall_in = 1'b0;
assign rnode_375to376_bb3_reduction_0_i283_0_NO_SHIFT_REG = rnode_375to376_bb3_reduction_0_i283_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_reduction_0_i283_0_stall_in_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_lnot14_i232_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_1_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_valid_out_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_stall_in_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_lnot14_i232_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_lnot14_i232_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_lnot14_i232_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_lnot14_i232_0_stall_in_0_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_lnot14_i232_0_valid_out_0_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_lnot14_i232_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3_lnot14_i232),
	.data_out(rnode_375to376_bb3_lnot14_i232_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_lnot14_i232_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_lnot14_i232_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3_lnot14_i232_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_lnot14_i232_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_lnot14_i232_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_lnot14_i232_stall_in_1 = 1'b0;
assign rnode_375to376_bb3_lnot14_i232_0_stall_in_0_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_lnot14_i232_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_lnot14_i232_0_NO_SHIFT_REG = rnode_375to376_bb3_lnot14_i232_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_lnot14_i232_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_lnot14_i232_1_NO_SHIFT_REG = rnode_375to376_bb3_lnot14_i232_0_reg_376_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_reduction_6_i246_0_valid_out_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_6_i246_0_stall_in_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_6_i246_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_6_i246_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_6_i246_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_6_i246_0_valid_out_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_6_i246_0_stall_in_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_reduction_6_i246_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_reduction_6_i246_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_reduction_6_i246_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_reduction_6_i246_0_stall_in_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_reduction_6_i246_0_valid_out_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_reduction_6_i246_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3_reduction_6_i246),
	.data_out(rnode_375to376_bb3_reduction_6_i246_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_reduction_6_i246_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_reduction_6_i246_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3_reduction_6_i246_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_reduction_6_i246_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_reduction_6_i246_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_reduction_6_i246_stall_in = 1'b0;
assign rnode_375to376_bb3_reduction_6_i246_0_NO_SHIFT_REG = rnode_375to376_bb3_reduction_6_i246_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_reduction_6_i246_0_stall_in_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_reduction_6_i246_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_375to376_bb3_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_375to376_bb3_xor_i224_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_xor_i224_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_375to376_bb3_xor_i224_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_xor_i224_0_valid_out_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_xor_i224_0_stall_in_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_xor_i224_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_xor_i224_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_xor_i224_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_xor_i224_0_stall_in_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_xor_i224_0_valid_out_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_xor_i224_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3_xor_i224),
	.data_out(rnode_375to376_bb3_xor_i224_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_xor_i224_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_xor_i224_0_reg_376_fifo.DATA_WIDTH = 32;
defparam rnode_375to376_bb3_xor_i224_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_xor_i224_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_xor_i224_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_xor_i224_stall_in = 1'b0;
assign rnode_375to376_bb3_xor_i224_0_NO_SHIFT_REG = rnode_375to376_bb3_xor_i224_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_xor_i224_0_stall_in_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3_cmp11_i231_0_valid_out_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp11_i231_0_stall_in_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp11_i231_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp11_i231_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp11_i231_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp11_i231_0_valid_out_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp11_i231_0_stall_in_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3_cmp11_i231_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3_cmp11_i231_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3_cmp11_i231_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3_cmp11_i231_0_stall_in_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3_cmp11_i231_0_valid_out_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3_cmp11_i231_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3_cmp11_i231),
	.data_out(rnode_375to376_bb3_cmp11_i231_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3_cmp11_i231_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3_cmp11_i231_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3_cmp11_i231_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3_cmp11_i231_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3_cmp11_i231_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp11_i231_stall_in_5 = 1'b0;
assign rnode_375to376_bb3_cmp11_i231_0_NO_SHIFT_REG = rnode_375to376_bb3_cmp11_i231_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3_cmp11_i231_0_stall_in_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_cmp11_i231_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb3_mul_i_i258_inputs_ready;
 reg local_bb3_mul_i_i258_valid_out_0_NO_SHIFT_REG;
wire local_bb3_mul_i_i258_stall_in_0;
 reg local_bb3_mul_i_i258_valid_out_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i258_stall_in_1;
wire local_bb3_mul_i_i258_output_regs_ready;
wire [63:0] local_bb3_mul_i_i258;
 reg local_bb3_mul_i_i258_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_mul_i_i258_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i258_causedstall;

acl_int_mult int_module_local_bb3_mul_i_i258 (
	.clock(clock),
	.dataa(((local_bb3_conv1_i_i257 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb3_conv_i_i256 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb3_mul_i_i258_output_regs_ready),
	.result(local_bb3_mul_i_i258)
);

defparam int_module_local_bb3_mul_i_i258.INPUT1_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i258.INPUT2_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i258.OUTPUT_WIDTH = 64;
defparam int_module_local_bb3_mul_i_i258.LATENCY = 3;
defparam int_module_local_bb3_mul_i_i258.SIGNED = 0;

assign local_bb3_mul_i_i258_inputs_ready = 1'b1;
assign local_bb3_mul_i_i258_output_regs_ready = 1'b1;
assign local_bb3_conv1_i_i257_stall_in = 1'b0;
assign local_bb3_conv_i_i256_stall_in = 1'b0;
assign local_bb3_mul_i_i258_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i258_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i258_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i258_output_regs_ready)
		begin
			local_bb3_mul_i_i258_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i258_valid_pipe_1_NO_SHIFT_REG <= local_bb3_mul_i_i258_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i258_output_regs_ready)
		begin
			local_bb3_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_mul_i_i258_stall_in_0))
			begin
				local_bb3_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_mul_i_i258_stall_in_1))
			begin
				local_bb3_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3__mux9_mux_i236_0_valid_out_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux9_mux_i236_0_stall_in_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux9_mux_i236_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux9_mux_i236_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux9_mux_i236_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux9_mux_i236_0_valid_out_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux9_mux_i236_0_stall_in_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux9_mux_i236_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3__mux9_mux_i236_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3__mux9_mux_i236_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3__mux9_mux_i236_0_stall_in_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3__mux9_mux_i236_0_valid_out_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3__mux9_mux_i236_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3__mux9_mux_i236),
	.data_out(rnode_375to376_bb3__mux9_mux_i236_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3__mux9_mux_i236_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3__mux9_mux_i236_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3__mux9_mux_i236_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3__mux9_mux_i236_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3__mux9_mux_i236_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__mux9_mux_i236_stall_in = 1'b0;
assign rnode_375to376_bb3__mux9_mux_i236_0_NO_SHIFT_REG = rnode_375to376_bb3__mux9_mux_i236_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3__mux9_mux_i236_0_stall_in_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3__mux9_mux_i236_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_valid_out_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_stall_in_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_inputs_ready_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_valid_out_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_stall_in_reg_376_NO_SHIFT_REG;
 logic rnode_375to376_bb3__mux_mux_mux_i242_0_stall_out_reg_376_NO_SHIFT_REG;

acl_data_fifo rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_375to376_bb3__mux_mux_mux_i242_0_stall_in_reg_376_NO_SHIFT_REG),
	.valid_out(rnode_375to376_bb3__mux_mux_mux_i242_0_valid_out_reg_376_NO_SHIFT_REG),
	.stall_out(rnode_375to376_bb3__mux_mux_mux_i242_0_stall_out_reg_376_NO_SHIFT_REG),
	.data_in(local_bb3__mux_mux_mux_i242),
	.data_out(rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_NO_SHIFT_REG)
);

defparam rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_fifo.DEPTH = 1;
defparam rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_fifo.DATA_WIDTH = 1;
defparam rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_fifo.IMPL = "shift_reg";

assign rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__mux_mux_mux_i242_stall_in = 1'b0;
assign rnode_375to376_bb3__mux_mux_mux_i242_0_NO_SHIFT_REG = rnode_375to376_bb3__mux_mux_mux_i242_0_reg_376_NO_SHIFT_REG;
assign rnode_375to376_bb3__mux_mux_mux_i242_0_stall_in_reg_376_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3__mux_mux_mux_i242_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_376to377_bb3_add_i265_0_valid_out_NO_SHIFT_REG;
 logic rnode_376to377_bb3_add_i265_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_376to377_bb3_add_i265_0_NO_SHIFT_REG;
 logic rnode_376to377_bb3_add_i265_0_reg_377_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_376to377_bb3_add_i265_0_reg_377_NO_SHIFT_REG;
 logic rnode_376to377_bb3_add_i265_0_valid_out_reg_377_NO_SHIFT_REG;
 logic rnode_376to377_bb3_add_i265_0_stall_in_reg_377_NO_SHIFT_REG;
 logic rnode_376to377_bb3_add_i265_0_stall_out_reg_377_NO_SHIFT_REG;

acl_data_fifo rnode_376to377_bb3_add_i265_0_reg_377_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_376to377_bb3_add_i265_0_reg_377_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_376to377_bb3_add_i265_0_stall_in_reg_377_NO_SHIFT_REG),
	.valid_out(rnode_376to377_bb3_add_i265_0_valid_out_reg_377_NO_SHIFT_REG),
	.stall_out(rnode_376to377_bb3_add_i265_0_stall_out_reg_377_NO_SHIFT_REG),
	.data_in((rnode_375to376_bb3_add_i265_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_376to377_bb3_add_i265_0_reg_377_NO_SHIFT_REG)
);

defparam rnode_376to377_bb3_add_i265_0_reg_377_fifo.DEPTH = 1;
defparam rnode_376to377_bb3_add_i265_0_reg_377_fifo.DATA_WIDTH = 32;
defparam rnode_376to377_bb3_add_i265_0_reg_377_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_376to377_bb3_add_i265_0_reg_377_fifo.IMPL = "shift_reg";

assign rnode_376to377_bb3_add_i265_0_reg_377_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_add_i265_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_376to377_bb3_add_i265_0_NO_SHIFT_REG = rnode_376to377_bb3_add_i265_0_reg_377_NO_SHIFT_REG;
assign rnode_376to377_bb3_add_i265_0_stall_in_reg_377_NO_SHIFT_REG = 1'b0;
assign rnode_376to377_bb3_add_i265_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__26_demorgan_i249_stall_local;
wire local_bb3__26_demorgan_i249;

assign local_bb3__26_demorgan_i249 = (rnode_375to376_bb3_cmp_i230_1_NO_SHIFT_REG | rnode_375to376_bb3_brmerge10_demorgan_i235_1_NO_SHIFT_REG);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_376to379_bb3_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_376to379_bb3_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_376to379_bb3_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_376to379_bb3_reduction_0_i283_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic rnode_376to379_bb3_reduction_0_i283_0_reg_379_NO_SHIFT_REG;
 logic rnode_376to379_bb3_reduction_0_i283_0_valid_out_reg_379_NO_SHIFT_REG;
 logic rnode_376to379_bb3_reduction_0_i283_0_stall_in_reg_379_NO_SHIFT_REG;
 logic rnode_376to379_bb3_reduction_0_i283_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_376to379_bb3_reduction_0_i283_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_376to379_bb3_reduction_0_i283_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_376to379_bb3_reduction_0_i283_0_stall_in_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_376to379_bb3_reduction_0_i283_0_valid_out_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_376to379_bb3_reduction_0_i283_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in(rnode_375to376_bb3_reduction_0_i283_0_NO_SHIFT_REG),
	.data_out(rnode_376to379_bb3_reduction_0_i283_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_376to379_bb3_reduction_0_i283_0_reg_379_fifo.DEPTH = 3;
defparam rnode_376to379_bb3_reduction_0_i283_0_reg_379_fifo.DATA_WIDTH = 1;
defparam rnode_376to379_bb3_reduction_0_i283_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_376to379_bb3_reduction_0_i283_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_376to379_bb3_reduction_0_i283_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_376to379_bb3_reduction_0_i283_0_NO_SHIFT_REG = rnode_376to379_bb3_reduction_0_i283_0_reg_379_NO_SHIFT_REG;
assign rnode_376to379_bb3_reduction_0_i283_0_stall_in_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_376to379_bb3_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_not_i251_stall_local;
wire local_bb3_lnot14_not_i251;

assign local_bb3_lnot14_not_i251 = (rnode_375to376_bb3_lnot14_i232_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3__24_i247_stall_local;
wire local_bb3__24_i247;

assign local_bb3__24_i247 = (rnode_375to376_bb3_cmp_i230_0_NO_SHIFT_REG ? rnode_375to376_bb3_reduction_6_i246_0_NO_SHIFT_REG : rnode_375to376_bb3_brmerge10_demorgan_i235_0_NO_SHIFT_REG);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_376to379_bb3_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_376to379_bb3_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_376to379_bb3_xor_i224_0_NO_SHIFT_REG;
 logic rnode_376to379_bb3_xor_i224_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_376to379_bb3_xor_i224_0_reg_379_NO_SHIFT_REG;
 logic rnode_376to379_bb3_xor_i224_0_valid_out_reg_379_NO_SHIFT_REG;
 logic rnode_376to379_bb3_xor_i224_0_stall_in_reg_379_NO_SHIFT_REG;
 logic rnode_376to379_bb3_xor_i224_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_376to379_bb3_xor_i224_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_376to379_bb3_xor_i224_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_376to379_bb3_xor_i224_0_stall_in_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_376to379_bb3_xor_i224_0_valid_out_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_376to379_bb3_xor_i224_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in(rnode_375to376_bb3_xor_i224_0_NO_SHIFT_REG),
	.data_out(rnode_376to379_bb3_xor_i224_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_376to379_bb3_xor_i224_0_reg_379_fifo.DEPTH = 3;
defparam rnode_376to379_bb3_xor_i224_0_reg_379_fifo.DATA_WIDTH = 32;
defparam rnode_376to379_bb3_xor_i224_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_376to379_bb3_xor_i224_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_376to379_bb3_xor_i224_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_375to376_bb3_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_376to379_bb3_xor_i224_0_NO_SHIFT_REG = rnode_376to379_bb3_xor_i224_0_reg_379_NO_SHIFT_REG;
assign rnode_376to379_bb3_xor_i224_0_stall_in_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_376to379_bb3_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u56_valid_out;
wire local_bb3_var__u56_stall_in;
wire local_bb3_var__u56_inputs_ready;
wire local_bb3_var__u56_stall_local;
wire local_bb3_var__u56;

assign local_bb3_var__u56_inputs_ready = (rnode_375to376_bb3_cmp_i230_0_valid_out_3_NO_SHIFT_REG & rnode_375to376_bb3_cmp11_i231_0_valid_out_NO_SHIFT_REG);
assign local_bb3_var__u56 = (rnode_375to376_bb3_cmp_i230_3_NO_SHIFT_REG | rnode_375to376_bb3_cmp11_i231_0_NO_SHIFT_REG);
assign local_bb3_var__u56_valid_out = 1'b1;
assign rnode_375to376_bb3_cmp_i230_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_cmp11_i231_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_conv3_i_i259_stall_local;
wire [31:0] local_bb3_conv3_i_i259;
wire [63:0] local_bb3_conv3_i_i259$ps;

assign local_bb3_conv3_i_i259$ps = (local_bb3_mul_i_i258 & 64'hFFFFFFFFFFFF);
assign local_bb3_conv3_i_i259 = local_bb3_conv3_i_i259$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_var__u57_stall_local;
wire [63:0] local_bb3_var__u57;

assign local_bb3_var__u57 = ((local_bb3_mul_i_i258 & 64'hFFFFFFFFFFFF) >> 64'h18);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_377to378_bb3_add_i265_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_377to378_bb3_add_i265_0_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_377to378_bb3_add_i265_1_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_377to378_bb3_add_i265_2_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_reg_378_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_377to378_bb3_add_i265_0_reg_378_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_valid_out_0_reg_378_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_stall_in_0_reg_378_NO_SHIFT_REG;
 logic rnode_377to378_bb3_add_i265_0_stall_out_reg_378_NO_SHIFT_REG;

acl_data_fifo rnode_377to378_bb3_add_i265_0_reg_378_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_377to378_bb3_add_i265_0_reg_378_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_377to378_bb3_add_i265_0_stall_in_0_reg_378_NO_SHIFT_REG),
	.valid_out(rnode_377to378_bb3_add_i265_0_valid_out_0_reg_378_NO_SHIFT_REG),
	.stall_out(rnode_377to378_bb3_add_i265_0_stall_out_reg_378_NO_SHIFT_REG),
	.data_in((rnode_376to377_bb3_add_i265_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_377to378_bb3_add_i265_0_reg_378_NO_SHIFT_REG)
);

defparam rnode_377to378_bb3_add_i265_0_reg_378_fifo.DEPTH = 1;
defparam rnode_377to378_bb3_add_i265_0_reg_378_fifo.DATA_WIDTH = 32;
defparam rnode_377to378_bb3_add_i265_0_reg_378_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_377to378_bb3_add_i265_0_reg_378_fifo.IMPL = "shift_reg";

assign rnode_377to378_bb3_add_i265_0_reg_378_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_376to377_bb3_add_i265_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_377to378_bb3_add_i265_0_stall_in_0_reg_378_NO_SHIFT_REG = 1'b0;
assign rnode_377to378_bb3_add_i265_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_377to378_bb3_add_i265_0_NO_SHIFT_REG = rnode_377to378_bb3_add_i265_0_reg_378_NO_SHIFT_REG;
assign rnode_377to378_bb3_add_i265_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_377to378_bb3_add_i265_1_NO_SHIFT_REG = rnode_377to378_bb3_add_i265_0_reg_378_NO_SHIFT_REG;
assign rnode_377to378_bb3_add_i265_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_377to378_bb3_add_i265_2_NO_SHIFT_REG = rnode_377to378_bb3_add_i265_0_reg_378_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_379to380_bb3_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_379to380_bb3_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_379to380_bb3_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_379to380_bb3_reduction_0_i283_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic rnode_379to380_bb3_reduction_0_i283_0_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_reduction_0_i283_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_reduction_0_i283_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_reduction_0_i283_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_379to380_bb3_reduction_0_i283_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_379to380_bb3_reduction_0_i283_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_379to380_bb3_reduction_0_i283_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_379to380_bb3_reduction_0_i283_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_379to380_bb3_reduction_0_i283_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(rnode_376to379_bb3_reduction_0_i283_0_NO_SHIFT_REG),
	.data_out(rnode_379to380_bb3_reduction_0_i283_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_379to380_bb3_reduction_0_i283_0_reg_380_fifo.DEPTH = 1;
defparam rnode_379to380_bb3_reduction_0_i283_0_reg_380_fifo.DATA_WIDTH = 1;
defparam rnode_379to380_bb3_reduction_0_i283_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_379to380_bb3_reduction_0_i283_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_379to380_bb3_reduction_0_i283_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_376to379_bb3_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_reduction_0_i283_0_NO_SHIFT_REG = rnode_379to380_bb3_reduction_0_i283_0_reg_380_NO_SHIFT_REG;
assign rnode_379to380_bb3_reduction_0_i283_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__28_i252_stall_local;
wire local_bb3__28_i252;

assign local_bb3__28_i252 = (rnode_375to376_bb3_cmp_i230_2_NO_SHIFT_REG & local_bb3_lnot14_not_i251);

// This section implements an unregistered operation.
// 
wire local_bb3__25_i248_stall_local;
wire local_bb3__25_i248;

assign local_bb3__25_i248 = (local_bb3__24_i247 ? rnode_375to376_bb3_lnot14_i232_0_NO_SHIFT_REG : rnode_375to376_bb3__mux_mux_mux_i242_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_379to380_bb3_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_379to380_bb3_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_379to380_bb3_xor_i224_0_NO_SHIFT_REG;
 logic rnode_379to380_bb3_xor_i224_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_379to380_bb3_xor_i224_0_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_xor_i224_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_xor_i224_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_xor_i224_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_379to380_bb3_xor_i224_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_379to380_bb3_xor_i224_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_379to380_bb3_xor_i224_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_379to380_bb3_xor_i224_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_379to380_bb3_xor_i224_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(rnode_376to379_bb3_xor_i224_0_NO_SHIFT_REG),
	.data_out(rnode_379to380_bb3_xor_i224_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_379to380_bb3_xor_i224_0_reg_380_fifo.DEPTH = 1;
defparam rnode_379to380_bb3_xor_i224_0_reg_380_fifo.DATA_WIDTH = 32;
defparam rnode_379to380_bb3_xor_i224_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_379to380_bb3_xor_i224_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_379to380_bb3_xor_i224_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_376to379_bb3_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_xor_i224_0_NO_SHIFT_REG = rnode_379to380_bb3_xor_i224_0_reg_380_NO_SHIFT_REG;
assign rnode_379to380_bb3_xor_i224_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_376to378_bb3_var__u56_0_valid_out_NO_SHIFT_REG;
 logic rnode_376to378_bb3_var__u56_0_stall_in_NO_SHIFT_REG;
 logic rnode_376to378_bb3_var__u56_0_NO_SHIFT_REG;
 logic rnode_376to378_bb3_var__u56_0_reg_378_inputs_ready_NO_SHIFT_REG;
 logic rnode_376to378_bb3_var__u56_0_reg_378_NO_SHIFT_REG;
 logic rnode_376to378_bb3_var__u56_0_valid_out_reg_378_NO_SHIFT_REG;
 logic rnode_376to378_bb3_var__u56_0_stall_in_reg_378_NO_SHIFT_REG;
 logic rnode_376to378_bb3_var__u56_0_stall_out_reg_378_NO_SHIFT_REG;

acl_data_fifo rnode_376to378_bb3_var__u56_0_reg_378_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_376to378_bb3_var__u56_0_reg_378_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_376to378_bb3_var__u56_0_stall_in_reg_378_NO_SHIFT_REG),
	.valid_out(rnode_376to378_bb3_var__u56_0_valid_out_reg_378_NO_SHIFT_REG),
	.stall_out(rnode_376to378_bb3_var__u56_0_stall_out_reg_378_NO_SHIFT_REG),
	.data_in(local_bb3_var__u56),
	.data_out(rnode_376to378_bb3_var__u56_0_reg_378_NO_SHIFT_REG)
);

defparam rnode_376to378_bb3_var__u56_0_reg_378_fifo.DEPTH = 2;
defparam rnode_376to378_bb3_var__u56_0_reg_378_fifo.DATA_WIDTH = 1;
defparam rnode_376to378_bb3_var__u56_0_reg_378_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_376to378_bb3_var__u56_0_reg_378_fifo.IMPL = "shift_reg";

assign rnode_376to378_bb3_var__u56_0_reg_378_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u56_stall_in = 1'b0;
assign rnode_376to378_bb3_var__u56_0_NO_SHIFT_REG = rnode_376to378_bb3_var__u56_0_reg_378_NO_SHIFT_REG;
assign rnode_376to378_bb3_var__u56_0_stall_in_reg_378_NO_SHIFT_REG = 1'b0;
assign rnode_376to378_bb3_var__u56_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i16_i262_stall_local;
wire [31:0] local_bb3_shr_i16_i262;

assign local_bb3_shr_i16_i262 = (local_bb3_conv3_i_i259 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i18_i264_stall_local;
wire [31:0] local_bb3_shl1_i18_i264;

assign local_bb3_shl1_i18_i264 = (local_bb3_conv3_i_i259 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u58_stall_local;
wire [31:0] local_bb3_var__u58;

assign local_bb3_var__u58 = (local_bb3_conv3_i_i259 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i_i272_stall_local;
wire [31:0] local_bb3_shl1_i_i272;

assign local_bb3_shl1_i_i272 = (local_bb3_conv3_i_i259 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb3__tr_i260_stall_local;
wire [31:0] local_bb3__tr_i260;
wire [63:0] local_bb3__tr_i260$ps;

assign local_bb3__tr_i260$ps = (local_bb3_var__u57 & 64'hFFFFFF);
assign local_bb3__tr_i260 = local_bb3__tr_i260$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_inc_i268_stall_local;
wire [31:0] local_bb3_inc_i268;

assign local_bb3_inc_i268 = ((rnode_377to378_bb3_add_i265_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp50_not_i273_stall_local;
wire local_bb3_cmp50_not_i273;

assign local_bb3_cmp50_not_i273 = ((rnode_377to378_bb3_add_i265_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb3__27_i250_stall_local;
wire local_bb3__27_i250;

assign local_bb3__27_i250 = (local_bb3__26_demorgan_i249 ? local_bb3__25_i248 : rnode_375to376_bb3__mux9_mux_i236_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_and4_i225_stall_local;
wire [31:0] local_bb3_and4_i225;

assign local_bb3_and4_i225 = (rnode_379to380_bb3_xor_i224_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i_i270_stall_local;
wire [31:0] local_bb3_shr_i_i270;

assign local_bb3_shr_i_i270 = ((local_bb3_var__u58 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i15_i261_stall_local;
wire [31:0] local_bb3_shl_i15_i261;

assign local_bb3_shl_i15_i261 = ((local_bb3__tr_i260 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb3_and48_i266_stall_local;
wire [31:0] local_bb3_and48_i266;

assign local_bb3_and48_i266 = ((local_bb3__tr_i260 & 32'hFFFFFF) & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3__29_i253_valid_out;
wire local_bb3__29_i253_stall_in;
wire local_bb3__29_i253_inputs_ready;
wire local_bb3__29_i253_stall_local;
wire local_bb3__29_i253;

assign local_bb3__29_i253_inputs_ready = (rnode_375to376_bb3_lnot14_i232_0_valid_out_0_NO_SHIFT_REG & rnode_375to376_bb3__mux_mux_mux_i242_0_valid_out_NO_SHIFT_REG & rnode_375to376_bb3__mux9_mux_i236_0_valid_out_NO_SHIFT_REG & rnode_375to376_bb3_cmp_i230_0_valid_out_0_NO_SHIFT_REG & rnode_375to376_bb3_reduction_6_i246_0_valid_out_NO_SHIFT_REG & rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_0_NO_SHIFT_REG & rnode_375to376_bb3_cmp_i230_0_valid_out_1_NO_SHIFT_REG & rnode_375to376_bb3_brmerge10_demorgan_i235_0_valid_out_1_NO_SHIFT_REG & rnode_375to376_bb3_lnot14_i232_0_valid_out_1_NO_SHIFT_REG & rnode_375to376_bb3_cmp_i230_0_valid_out_2_NO_SHIFT_REG);
assign local_bb3__29_i253 = (local_bb3__28_i252 | local_bb3__27_i250);
assign local_bb3__29_i253_valid_out = 1'b1;
assign rnode_375to376_bb3_lnot14_i232_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3__mux_mux_mux_i242_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3__mux9_mux_i236_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_cmp_i230_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_reduction_6_i246_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_cmp_i230_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_brmerge10_demorgan_i235_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_lnot14_i232_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_375to376_bb3_cmp_i230_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_or_i17_i263_stall_local;
wire [31:0] local_bb3_or_i17_i263;

assign local_bb3_or_i17_i263 = ((local_bb3_shl_i15_i261 & 32'hFFFF00) | (local_bb3_shr_i16_i262 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool49_i267_stall_local;
wire local_bb3_tobool49_i267;

assign local_bb3_tobool49_i267 = ((local_bb3_and48_i266 & 32'h800000) == 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_376to377_bb3__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_376to377_bb3__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_376to377_bb3__29_i253_0_NO_SHIFT_REG;
 logic rnode_376to377_bb3__29_i253_0_reg_377_inputs_ready_NO_SHIFT_REG;
 logic rnode_376to377_bb3__29_i253_0_reg_377_NO_SHIFT_REG;
 logic rnode_376to377_bb3__29_i253_0_valid_out_reg_377_NO_SHIFT_REG;
 logic rnode_376to377_bb3__29_i253_0_stall_in_reg_377_NO_SHIFT_REG;
 logic rnode_376to377_bb3__29_i253_0_stall_out_reg_377_NO_SHIFT_REG;

acl_data_fifo rnode_376to377_bb3__29_i253_0_reg_377_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_376to377_bb3__29_i253_0_reg_377_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_376to377_bb3__29_i253_0_stall_in_reg_377_NO_SHIFT_REG),
	.valid_out(rnode_376to377_bb3__29_i253_0_valid_out_reg_377_NO_SHIFT_REG),
	.stall_out(rnode_376to377_bb3__29_i253_0_stall_out_reg_377_NO_SHIFT_REG),
	.data_in(local_bb3__29_i253),
	.data_out(rnode_376to377_bb3__29_i253_0_reg_377_NO_SHIFT_REG)
);

defparam rnode_376to377_bb3__29_i253_0_reg_377_fifo.DEPTH = 1;
defparam rnode_376to377_bb3__29_i253_0_reg_377_fifo.DATA_WIDTH = 1;
defparam rnode_376to377_bb3__29_i253_0_reg_377_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_376to377_bb3__29_i253_0_reg_377_fifo.IMPL = "shift_reg";

assign rnode_376to377_bb3__29_i253_0_reg_377_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__29_i253_stall_in = 1'b0;
assign rnode_376to377_bb3__29_i253_0_NO_SHIFT_REG = rnode_376to377_bb3__29_i253_0_reg_377_NO_SHIFT_REG;
assign rnode_376to377_bb3__29_i253_0_stall_in_reg_377_NO_SHIFT_REG = 1'b0;
assign rnode_376to377_bb3__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i_i269_stall_local;
wire [31:0] local_bb3_shl_i_i269;

assign local_bb3_shl_i_i269 = ((local_bb3_or_i17_i263 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__31_i274_stall_local;
wire local_bb3__31_i274;

assign local_bb3__31_i274 = (local_bb3_tobool49_i267 & local_bb3_cmp50_not_i273);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_377to379_bb3__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_377to379_bb3__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_377to379_bb3__29_i253_0_NO_SHIFT_REG;
 logic rnode_377to379_bb3__29_i253_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic rnode_377to379_bb3__29_i253_0_reg_379_NO_SHIFT_REG;
 logic rnode_377to379_bb3__29_i253_0_valid_out_reg_379_NO_SHIFT_REG;
 logic rnode_377to379_bb3__29_i253_0_stall_in_reg_379_NO_SHIFT_REG;
 logic rnode_377to379_bb3__29_i253_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_377to379_bb3__29_i253_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_377to379_bb3__29_i253_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_377to379_bb3__29_i253_0_stall_in_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_377to379_bb3__29_i253_0_valid_out_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_377to379_bb3__29_i253_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in(rnode_376to377_bb3__29_i253_0_NO_SHIFT_REG),
	.data_out(rnode_377to379_bb3__29_i253_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_377to379_bb3__29_i253_0_reg_379_fifo.DEPTH = 2;
defparam rnode_377to379_bb3__29_i253_0_reg_379_fifo.DATA_WIDTH = 1;
defparam rnode_377to379_bb3__29_i253_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_377to379_bb3__29_i253_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_377to379_bb3__29_i253_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_376to377_bb3__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_377to379_bb3__29_i253_0_NO_SHIFT_REG = rnode_377to379_bb3__29_i253_0_reg_379_NO_SHIFT_REG;
assign rnode_377to379_bb3__29_i253_0_stall_in_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_377to379_bb3__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_or_i_i271_stall_local;
wire [31:0] local_bb3_or_i_i271;

assign local_bb3_or_i_i271 = ((local_bb3_shl_i_i269 & 32'h1FFFFFE) | (local_bb3_shr_i_i270 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__32_i275_stall_local;
wire [31:0] local_bb3__32_i275;

assign local_bb3__32_i275 = (local_bb3__31_i274 ? (local_bb3_shl1_i_i272 & 32'hFFFFFE00) : (local_bb3_shl1_i18_i264 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__36_i279_stall_local;
wire [31:0] local_bb3__36_i279;

assign local_bb3__36_i279 = (local_bb3__31_i274 ? (rnode_377to378_bb3_add_i265_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_379to380_bb3__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_379to380_bb3__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_379to380_bb3__29_i253_0_NO_SHIFT_REG;
 logic rnode_379to380_bb3__29_i253_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic rnode_379to380_bb3__29_i253_0_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3__29_i253_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3__29_i253_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3__29_i253_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_379to380_bb3__29_i253_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_379to380_bb3__29_i253_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_379to380_bb3__29_i253_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_379to380_bb3__29_i253_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_379to380_bb3__29_i253_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(rnode_377to379_bb3__29_i253_0_NO_SHIFT_REG),
	.data_out(rnode_379to380_bb3__29_i253_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_379to380_bb3__29_i253_0_reg_380_fifo.DEPTH = 1;
defparam rnode_379to380_bb3__29_i253_0_reg_380_fifo.DATA_WIDTH = 1;
defparam rnode_379to380_bb3__29_i253_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_379to380_bb3__29_i253_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_379to380_bb3__29_i253_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_377to379_bb3__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3__29_i253_0_NO_SHIFT_REG = rnode_379to380_bb3__29_i253_0_reg_380_NO_SHIFT_REG;
assign rnode_379to380_bb3__29_i253_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__34_i277_stall_local;
wire [31:0] local_bb3__34_i277;

assign local_bb3__34_i277 = (local_bb3__31_i274 ? (local_bb3_or_i_i271 & 32'h1FFFFFF) : (local_bb3_or_i17_i263 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__33_i276_stall_local;
wire [31:0] local_bb3__33_i276;

assign local_bb3__33_i276 = (local_bb3_tobool49_i267 ? (local_bb3__32_i275 & 32'hFFFFFF00) : (local_bb3_shl1_i18_i264 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__37_i280_stall_local;
wire [31:0] local_bb3__37_i280;

assign local_bb3__37_i280 = (local_bb3_tobool49_i267 ? (local_bb3__36_i279 & 32'h1FF) : (local_bb3_inc_i268 & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb3__35_i278_stall_local;
wire [31:0] local_bb3__35_i278;

assign local_bb3__35_i278 = (local_bb3_tobool49_i267 ? (local_bb3__34_i277 & 32'h1FFFFFF) : (local_bb3_or_i17_i263 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp53_i281_stall_local;
wire local_bb3_cmp53_i281;

assign local_bb3_cmp53_i281 = ((local_bb3__37_i280 & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp68_i285_stall_local;
wire local_bb3_cmp68_i285;

assign local_bb3_cmp68_i285 = ((local_bb3__37_i280 & 32'h3FF) < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb3_sub_i287_stall_local;
wire [31:0] local_bb3_sub_i287;

assign local_bb3_sub_i287 = ((local_bb3__37_i280 & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp71_not_i302_stall_local;
wire local_bb3_cmp71_not_i302;

assign local_bb3_cmp71_not_i302 = ((local_bb3__37_i280 & 32'h3FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb3_and75_i286_stall_local;
wire [31:0] local_bb3_and75_i286;

assign local_bb3_and75_i286 = ((local_bb3__35_i278 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and83_i292_stall_local;
wire [31:0] local_bb3_and83_i292;

assign local_bb3_and83_i292 = ((local_bb3__35_i278 & 32'h1FFFFFF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or581_i282_stall_local;
wire local_bb3_or581_i282;

assign local_bb3_or581_i282 = (rnode_376to378_bb3_var__u56_0_NO_SHIFT_REG | local_bb3_cmp53_i281);

// This section implements an unregistered operation.
// 
wire local_bb3_and74_i288_stall_local;
wire [31:0] local_bb3_and74_i288;

assign local_bb3_and74_i288 = ((local_bb3_sub_i287 & 32'hFF800000) + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb3__33_i276_valid_out;
wire local_bb3__33_i276_stall_in;
wire local_bb3_cmp68_i285_valid_out;
wire local_bb3_cmp68_i285_stall_in;
wire local_bb3_cmp71_not_i302_valid_out;
wire local_bb3_cmp71_not_i302_stall_in;
wire local_bb3_and75_i286_valid_out;
wire local_bb3_and75_i286_stall_in;
wire local_bb3_and83_i292_valid_out;
wire local_bb3_and83_i292_stall_in;
wire local_bb3_or581_i282_valid_out;
wire local_bb3_or581_i282_stall_in;
wire local_bb3_shl_i289_valid_out;
wire local_bb3_shl_i289_stall_in;
wire local_bb3_shl_i289_inputs_ready;
wire local_bb3_shl_i289_stall_local;
wire [31:0] local_bb3_shl_i289;

assign local_bb3_shl_i289_inputs_ready = (local_bb3_mul_i_i258_valid_out_0_NO_SHIFT_REG & local_bb3_mul_i_i258_valid_out_1_NO_SHIFT_REG & rnode_377to378_bb3_add_i265_0_valid_out_1_NO_SHIFT_REG & rnode_377to378_bb3_add_i265_0_valid_out_0_NO_SHIFT_REG & rnode_377to378_bb3_add_i265_0_valid_out_2_NO_SHIFT_REG & rnode_376to378_bb3_var__u56_0_valid_out_NO_SHIFT_REG);
assign local_bb3_shl_i289 = ((local_bb3_and74_i288 & 32'hFF800000) & 32'h7F800000);
assign local_bb3__33_i276_valid_out = 1'b1;
assign local_bb3_cmp68_i285_valid_out = 1'b1;
assign local_bb3_cmp71_not_i302_valid_out = 1'b1;
assign local_bb3_and75_i286_valid_out = 1'b1;
assign local_bb3_and83_i292_valid_out = 1'b1;
assign local_bb3_or581_i282_valid_out = 1'b1;
assign local_bb3_shl_i289_valid_out = 1'b1;
assign local_bb3_mul_i_i258_stall_in_0 = 1'b0;
assign local_bb3_mul_i_i258_stall_in_1 = 1'b0;
assign rnode_377to378_bb3_add_i265_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_377to378_bb3_add_i265_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_377to378_bb3_add_i265_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_376to378_bb3_var__u56_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_378to379_bb3__33_i276_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_378to379_bb3__33_i276_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3__33_i276_0_NO_SHIFT_REG;
 logic rnode_378to379_bb3__33_i276_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_378to379_bb3__33_i276_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3__33_i276_1_NO_SHIFT_REG;
 logic rnode_378to379_bb3__33_i276_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3__33_i276_0_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3__33_i276_0_valid_out_0_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3__33_i276_0_stall_in_0_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3__33_i276_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_378to379_bb3__33_i276_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_378to379_bb3__33_i276_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_378to379_bb3__33_i276_0_stall_in_0_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_378to379_bb3__33_i276_0_valid_out_0_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_378to379_bb3__33_i276_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in((local_bb3__33_i276 & 32'hFFFFFF00)),
	.data_out(rnode_378to379_bb3__33_i276_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_378to379_bb3__33_i276_0_reg_379_fifo.DEPTH = 1;
defparam rnode_378to379_bb3__33_i276_0_reg_379_fifo.DATA_WIDTH = 32;
defparam rnode_378to379_bb3__33_i276_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_378to379_bb3__33_i276_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_378to379_bb3__33_i276_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__33_i276_stall_in = 1'b0;
assign rnode_378to379_bb3__33_i276_0_stall_in_0_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_378to379_bb3__33_i276_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_378to379_bb3__33_i276_0_NO_SHIFT_REG = rnode_378to379_bb3__33_i276_0_reg_379_NO_SHIFT_REG;
assign rnode_378to379_bb3__33_i276_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_378to379_bb3__33_i276_1_NO_SHIFT_REG = rnode_378to379_bb3__33_i276_0_reg_379_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_378to380_bb3_cmp68_i285_0_valid_out_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp68_i285_0_stall_in_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp68_i285_0_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp68_i285_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp68_i285_0_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp68_i285_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp68_i285_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp68_i285_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_378to380_bb3_cmp68_i285_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_378to380_bb3_cmp68_i285_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_378to380_bb3_cmp68_i285_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_378to380_bb3_cmp68_i285_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_378to380_bb3_cmp68_i285_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(local_bb3_cmp68_i285),
	.data_out(rnode_378to380_bb3_cmp68_i285_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_378to380_bb3_cmp68_i285_0_reg_380_fifo.DEPTH = 2;
defparam rnode_378to380_bb3_cmp68_i285_0_reg_380_fifo.DATA_WIDTH = 1;
defparam rnode_378to380_bb3_cmp68_i285_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_378to380_bb3_cmp68_i285_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_378to380_bb3_cmp68_i285_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp68_i285_stall_in = 1'b0;
assign rnode_378to380_bb3_cmp68_i285_0_NO_SHIFT_REG = rnode_378to380_bb3_cmp68_i285_0_reg_380_NO_SHIFT_REG;
assign rnode_378to380_bb3_cmp68_i285_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_378to380_bb3_cmp68_i285_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_378to380_bb3_cmp71_not_i302_0_valid_out_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp71_not_i302_0_stall_in_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp71_not_i302_0_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp71_not_i302_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp71_not_i302_0_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp71_not_i302_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp71_not_i302_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_cmp71_not_i302_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_378to380_bb3_cmp71_not_i302_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_378to380_bb3_cmp71_not_i302_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_378to380_bb3_cmp71_not_i302_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_378to380_bb3_cmp71_not_i302_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_378to380_bb3_cmp71_not_i302_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(local_bb3_cmp71_not_i302),
	.data_out(rnode_378to380_bb3_cmp71_not_i302_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_378to380_bb3_cmp71_not_i302_0_reg_380_fifo.DEPTH = 2;
defparam rnode_378to380_bb3_cmp71_not_i302_0_reg_380_fifo.DATA_WIDTH = 1;
defparam rnode_378to380_bb3_cmp71_not_i302_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_378to380_bb3_cmp71_not_i302_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_378to380_bb3_cmp71_not_i302_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp71_not_i302_stall_in = 1'b0;
assign rnode_378to380_bb3_cmp71_not_i302_0_NO_SHIFT_REG = rnode_378to380_bb3_cmp71_not_i302_0_reg_380_NO_SHIFT_REG;
assign rnode_378to380_bb3_cmp71_not_i302_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_378to380_bb3_cmp71_not_i302_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_378to379_bb3_and75_i286_0_valid_out_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and75_i286_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3_and75_i286_0_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and75_i286_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3_and75_i286_0_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and75_i286_0_valid_out_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and75_i286_0_stall_in_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and75_i286_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_378to379_bb3_and75_i286_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_378to379_bb3_and75_i286_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_378to379_bb3_and75_i286_0_stall_in_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_378to379_bb3_and75_i286_0_valid_out_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_378to379_bb3_and75_i286_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in((local_bb3_and75_i286 & 32'h7FFFFF)),
	.data_out(rnode_378to379_bb3_and75_i286_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_378to379_bb3_and75_i286_0_reg_379_fifo.DEPTH = 1;
defparam rnode_378to379_bb3_and75_i286_0_reg_379_fifo.DATA_WIDTH = 32;
defparam rnode_378to379_bb3_and75_i286_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_378to379_bb3_and75_i286_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_378to379_bb3_and75_i286_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and75_i286_stall_in = 1'b0;
assign rnode_378to379_bb3_and75_i286_0_NO_SHIFT_REG = rnode_378to379_bb3_and75_i286_0_reg_379_NO_SHIFT_REG;
assign rnode_378to379_bb3_and75_i286_0_stall_in_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_378to379_bb3_and75_i286_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_378to379_bb3_and83_i292_0_valid_out_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and83_i292_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3_and83_i292_0_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and83_i292_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3_and83_i292_0_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and83_i292_0_valid_out_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and83_i292_0_stall_in_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_and83_i292_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_378to379_bb3_and83_i292_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_378to379_bb3_and83_i292_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_378to379_bb3_and83_i292_0_stall_in_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_378to379_bb3_and83_i292_0_valid_out_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_378to379_bb3_and83_i292_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in((local_bb3_and83_i292 & 32'h1)),
	.data_out(rnode_378to379_bb3_and83_i292_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_378to379_bb3_and83_i292_0_reg_379_fifo.DEPTH = 1;
defparam rnode_378to379_bb3_and83_i292_0_reg_379_fifo.DATA_WIDTH = 32;
defparam rnode_378to379_bb3_and83_i292_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_378to379_bb3_and83_i292_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_378to379_bb3_and83_i292_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and83_i292_stall_in = 1'b0;
assign rnode_378to379_bb3_and83_i292_0_NO_SHIFT_REG = rnode_378to379_bb3_and83_i292_0_reg_379_NO_SHIFT_REG;
assign rnode_378to379_bb3_and83_i292_0_stall_in_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_378to379_bb3_and83_i292_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_378to380_bb3_or581_i282_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_1_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_valid_out_0_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_stall_in_0_reg_380_NO_SHIFT_REG;
 logic rnode_378to380_bb3_or581_i282_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_378to380_bb3_or581_i282_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_378to380_bb3_or581_i282_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_378to380_bb3_or581_i282_0_stall_in_0_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_378to380_bb3_or581_i282_0_valid_out_0_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_378to380_bb3_or581_i282_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(local_bb3_or581_i282),
	.data_out(rnode_378to380_bb3_or581_i282_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_378to380_bb3_or581_i282_0_reg_380_fifo.DEPTH = 2;
defparam rnode_378to380_bb3_or581_i282_0_reg_380_fifo.DATA_WIDTH = 1;
defparam rnode_378to380_bb3_or581_i282_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_378to380_bb3_or581_i282_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_378to380_bb3_or581_i282_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or581_i282_stall_in = 1'b0;
assign rnode_378to380_bb3_or581_i282_0_stall_in_0_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_378to380_bb3_or581_i282_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_378to380_bb3_or581_i282_0_NO_SHIFT_REG = rnode_378to380_bb3_or581_i282_0_reg_380_NO_SHIFT_REG;
assign rnode_378to380_bb3_or581_i282_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_378to380_bb3_or581_i282_1_NO_SHIFT_REG = rnode_378to380_bb3_or581_i282_0_reg_380_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_378to379_bb3_shl_i289_0_valid_out_NO_SHIFT_REG;
 logic rnode_378to379_bb3_shl_i289_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3_shl_i289_0_NO_SHIFT_REG;
 logic rnode_378to379_bb3_shl_i289_0_reg_379_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_378to379_bb3_shl_i289_0_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_shl_i289_0_valid_out_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_shl_i289_0_stall_in_reg_379_NO_SHIFT_REG;
 logic rnode_378to379_bb3_shl_i289_0_stall_out_reg_379_NO_SHIFT_REG;

acl_data_fifo rnode_378to379_bb3_shl_i289_0_reg_379_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_378to379_bb3_shl_i289_0_reg_379_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_378to379_bb3_shl_i289_0_stall_in_reg_379_NO_SHIFT_REG),
	.valid_out(rnode_378to379_bb3_shl_i289_0_valid_out_reg_379_NO_SHIFT_REG),
	.stall_out(rnode_378to379_bb3_shl_i289_0_stall_out_reg_379_NO_SHIFT_REG),
	.data_in((local_bb3_shl_i289 & 32'h7F800000)),
	.data_out(rnode_378to379_bb3_shl_i289_0_reg_379_NO_SHIFT_REG)
);

defparam rnode_378to379_bb3_shl_i289_0_reg_379_fifo.DEPTH = 1;
defparam rnode_378to379_bb3_shl_i289_0_reg_379_fifo.DATA_WIDTH = 32;
defparam rnode_378to379_bb3_shl_i289_0_reg_379_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_378to379_bb3_shl_i289_0_reg_379_fifo.IMPL = "shift_reg";

assign rnode_378to379_bb3_shl_i289_0_reg_379_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shl_i289_stall_in = 1'b0;
assign rnode_378to379_bb3_shl_i289_0_NO_SHIFT_REG = rnode_378to379_bb3_shl_i289_0_reg_379_NO_SHIFT_REG;
assign rnode_378to379_bb3_shl_i289_0_stall_in_reg_379_NO_SHIFT_REG = 1'b0;
assign rnode_378to379_bb3_shl_i289_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp77_i291_stall_local;
wire local_bb3_cmp77_i291;

assign local_bb3_cmp77_i291 = ((rnode_378to379_bb3__33_i276_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u59_stall_local;
wire local_bb3_var__u59;

assign local_bb3_var__u59 = ($signed((rnode_378to379_bb3__33_i276_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u60_stall_local;
wire [31:0] local_bb3_var__u60;

assign local_bb3_var__u60[31:1] = 31'h0;
assign local_bb3_var__u60[0] = rnode_378to380_bb3_cmp68_i285_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_tobool84_i293_stall_local;
wire local_bb3_tobool84_i293;

assign local_bb3_tobool84_i293 = ((rnode_378to379_bb3_and83_i292_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_2_i284_stall_local;
wire local_bb3_reduction_2_i284;

assign local_bb3_reduction_2_i284 = (rnode_379to380_bb3_reduction_0_i283_0_NO_SHIFT_REG | rnode_378to380_bb3_or581_i282_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_cond111_i310_stall_local;
wire [31:0] local_bb3_cond111_i310;

assign local_bb3_cond111_i310 = (rnode_378to380_bb3_or581_i282_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or76_i290_valid_out;
wire local_bb3_or76_i290_stall_in;
wire local_bb3_or76_i290_inputs_ready;
wire local_bb3_or76_i290_stall_local;
wire [31:0] local_bb3_or76_i290;

assign local_bb3_or76_i290_inputs_ready = (rnode_378to379_bb3_shl_i289_0_valid_out_NO_SHIFT_REG & rnode_378to379_bb3_and75_i286_0_valid_out_NO_SHIFT_REG);
assign local_bb3_or76_i290 = ((rnode_378to379_bb3_shl_i289_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_378to379_bb3_and75_i286_0_NO_SHIFT_REG & 32'h7FFFFF));
assign local_bb3_or76_i290_valid_out = 1'b1;
assign rnode_378to379_bb3_shl_i289_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_378to379_bb3_and75_i286_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__39_i294_stall_local;
wire local_bb3__39_i294;

assign local_bb3__39_i294 = (local_bb3_tobool84_i293 & local_bb3_var__u59);

// This section implements an unregistered operation.
// 
wire local_bb3_conv101_i305_stall_local;
wire [31:0] local_bb3_conv101_i305;

assign local_bb3_conv101_i305[31:1] = 31'h0;
assign local_bb3_conv101_i305[0] = local_bb3_reduction_2_i284;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_379to380_bb3_or76_i290_0_valid_out_NO_SHIFT_REG;
 logic rnode_379to380_bb3_or76_i290_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_379to380_bb3_or76_i290_0_NO_SHIFT_REG;
 logic rnode_379to380_bb3_or76_i290_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_379to380_bb3_or76_i290_0_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_or76_i290_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_or76_i290_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3_or76_i290_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_379to380_bb3_or76_i290_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_379to380_bb3_or76_i290_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_379to380_bb3_or76_i290_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_379to380_bb3_or76_i290_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_379to380_bb3_or76_i290_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in((local_bb3_or76_i290 & 32'h7FFFFFFF)),
	.data_out(rnode_379to380_bb3_or76_i290_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_379to380_bb3_or76_i290_0_reg_380_fifo.DEPTH = 1;
defparam rnode_379to380_bb3_or76_i290_0_reg_380_fifo.DATA_WIDTH = 32;
defparam rnode_379to380_bb3_or76_i290_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_379to380_bb3_or76_i290_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_379to380_bb3_or76_i290_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or76_i290_stall_in = 1'b0;
assign rnode_379to380_bb3_or76_i290_0_NO_SHIFT_REG = rnode_379to380_bb3_or76_i290_0_reg_380_NO_SHIFT_REG;
assign rnode_379to380_bb3_or76_i290_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_or76_i290_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__40_i295_valid_out;
wire local_bb3__40_i295_stall_in;
wire local_bb3__40_i295_inputs_ready;
wire local_bb3__40_i295_stall_local;
wire local_bb3__40_i295;

assign local_bb3__40_i295_inputs_ready = (rnode_378to379_bb3__33_i276_0_valid_out_0_NO_SHIFT_REG & rnode_378to379_bb3__33_i276_0_valid_out_1_NO_SHIFT_REG & rnode_378to379_bb3_and83_i292_0_valid_out_NO_SHIFT_REG);
assign local_bb3__40_i295 = (local_bb3_cmp77_i291 | local_bb3__39_i294);
assign local_bb3__40_i295_valid_out = 1'b1;
assign rnode_378to379_bb3__33_i276_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_378to379_bb3__33_i276_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_378to379_bb3_and83_i292_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_379to380_bb3__40_i295_0_valid_out_NO_SHIFT_REG;
 logic rnode_379to380_bb3__40_i295_0_stall_in_NO_SHIFT_REG;
 logic rnode_379to380_bb3__40_i295_0_NO_SHIFT_REG;
 logic rnode_379to380_bb3__40_i295_0_reg_380_inputs_ready_NO_SHIFT_REG;
 logic rnode_379to380_bb3__40_i295_0_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3__40_i295_0_valid_out_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3__40_i295_0_stall_in_reg_380_NO_SHIFT_REG;
 logic rnode_379to380_bb3__40_i295_0_stall_out_reg_380_NO_SHIFT_REG;

acl_data_fifo rnode_379to380_bb3__40_i295_0_reg_380_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_379to380_bb3__40_i295_0_reg_380_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_379to380_bb3__40_i295_0_stall_in_reg_380_NO_SHIFT_REG),
	.valid_out(rnode_379to380_bb3__40_i295_0_valid_out_reg_380_NO_SHIFT_REG),
	.stall_out(rnode_379to380_bb3__40_i295_0_stall_out_reg_380_NO_SHIFT_REG),
	.data_in(local_bb3__40_i295),
	.data_out(rnode_379to380_bb3__40_i295_0_reg_380_NO_SHIFT_REG)
);

defparam rnode_379to380_bb3__40_i295_0_reg_380_fifo.DEPTH = 1;
defparam rnode_379to380_bb3__40_i295_0_reg_380_fifo.DATA_WIDTH = 1;
defparam rnode_379to380_bb3__40_i295_0_reg_380_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_379to380_bb3__40_i295_0_reg_380_fifo.IMPL = "shift_reg";

assign rnode_379to380_bb3__40_i295_0_reg_380_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__40_i295_stall_in = 1'b0;
assign rnode_379to380_bb3__40_i295_0_NO_SHIFT_REG = rnode_379to380_bb3__40_i295_0_reg_380_NO_SHIFT_REG;
assign rnode_379to380_bb3__40_i295_0_stall_in_reg_380_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3__40_i295_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cond_i296_stall_local;
wire [31:0] local_bb3_cond_i296;

assign local_bb3_cond_i296[31:1] = 31'h0;
assign local_bb3_cond_i296[0] = rnode_379to380_bb3__40_i295_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_add87_i297_stall_local;
wire [31:0] local_bb3_add87_i297;

assign local_bb3_add87_i297 = ((local_bb3_cond_i296 & 32'h1) + (rnode_379to380_bb3_or76_i290_0_NO_SHIFT_REG & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_and88_i298_stall_local;
wire [31:0] local_bb3_and88_i298;

assign local_bb3_and88_i298 = (local_bb3_add87_i297 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and90_i300_stall_local;
wire [31:0] local_bb3_and90_i300;

assign local_bb3_and90_i300 = (local_bb3_add87_i297 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_or89_i299_stall_local;
wire [31:0] local_bb3_or89_i299;

assign local_bb3_or89_i299 = ((local_bb3_and88_i298 & 32'h7FFFFFFF) | (local_bb3_and4_i225 & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp91_i301_stall_local;
wire local_bb3_cmp91_i301;

assign local_bb3_cmp91_i301 = ((local_bb3_and90_i300 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge14_i303_stall_local;
wire local_bb3_brmerge14_i303;

assign local_bb3_brmerge14_i303 = (local_bb3_cmp91_i301 | rnode_378to380_bb3_cmp71_not_i302_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_conv99_i304_stall_local;
wire [31:0] local_bb3_conv99_i304;

assign local_bb3_conv99_i304 = (local_bb3_brmerge14_i303 ? (local_bb3_var__u60 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or102_i306_stall_local;
wire [31:0] local_bb3_or102_i306;

assign local_bb3_or102_i306 = ((local_bb3_conv99_i304 & 32'h1) | (local_bb3_conv101_i305 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool103_i307_stall_local;
wire local_bb3_tobool103_i307;

assign local_bb3_tobool103_i307 = ((local_bb3_or102_i306 & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cond107_i308_stall_local;
wire [31:0] local_bb3_cond107_i308;

assign local_bb3_cond107_i308 = (local_bb3_tobool103_i307 ? (local_bb3_and4_i225 & 32'h80000000) : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and108_i309_stall_local;
wire [31:0] local_bb3_and108_i309;

assign local_bb3_and108_i309 = (local_bb3_cond107_i308 & local_bb3_or89_i299);

// This section implements an unregistered operation.
// 
wire local_bb3_or112_i311_stall_local;
wire [31:0] local_bb3_or112_i311;

assign local_bb3_or112_i311 = (local_bb3_and108_i309 | (local_bb3_cond111_i310 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u61_stall_local;
wire [31:0] local_bb3_var__u61;

assign local_bb3_var__u61 = local_bb3_or112_i311;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u62_stall_local;
wire [31:0] local_bb3_var__u62;

assign local_bb3_var__u62 = (rnode_379to380_bb3__29_i253_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb3_var__u61);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u63_stall_local;
wire [31:0] local_bb3_var__u63;

assign local_bb3_var__u63 = local_bb3_var__u62;

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i193_stall_local;
wire [31:0] local_bb3_shr_i193;

assign local_bb3_shr_i193 = (local_bb3_var__u63 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_xor_i195_stall_local;
wire [31:0] local_bb3_xor_i195;

assign local_bb3_xor_i195 = (local_bb3_var__u25 ^ local_bb3_var__u63);

// This section implements an unregistered operation.
// 
wire local_bb3_and5_i_stall_local;
wire [31:0] local_bb3_and5_i;

assign local_bb3_and5_i = (local_bb3_var__u63 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i205_stall_local;
wire [31:0] local_bb3_or_i205;

assign local_bb3_or_i205 = ((local_bb3_and5_i & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_shr2_i_valid_out;
wire local_bb3_shr2_i_stall_in;
wire local_bb3_xor_i195_valid_out;
wire local_bb3_xor_i195_stall_in;
wire local_bb3_and6_i_valid_out_1;
wire local_bb3_and6_i_stall_in_1;
wire local_bb3_conv1_i_i_valid_out;
wire local_bb3_conv1_i_i_stall_in;
wire local_bb3_var__u62_valid_out_1;
wire local_bb3_var__u62_stall_in_1;
wire local_bb3_shr_i193_valid_out;
wire local_bb3_shr_i193_stall_in;
wire local_bb3_and5_i_valid_out_1;
wire local_bb3_and5_i_stall_in_1;
wire local_bb3_conv_i_i_valid_out;
wire local_bb3_conv_i_i_stall_in;
wire local_bb3_conv_i_i_inputs_ready;
wire local_bb3_conv_i_i_stall_local;
wire [63:0] local_bb3_conv_i_i;

assign local_bb3_conv_i_i_inputs_ready = (rnode_379to380_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG & rnode_379to380_bb3_xor_i224_0_valid_out_NO_SHIFT_REG & rnode_378to380_bb3_or581_i282_0_valid_out_1_NO_SHIFT_REG & rnode_379to380_bb3__29_i253_0_valid_out_NO_SHIFT_REG & rnode_378to380_bb3_or581_i282_0_valid_out_0_NO_SHIFT_REG & rnode_379to380_bb3_reduction_0_i283_0_valid_out_NO_SHIFT_REG & rnode_378to380_bb3_cmp68_i285_0_valid_out_NO_SHIFT_REG & rnode_378to380_bb3_cmp71_not_i302_0_valid_out_NO_SHIFT_REG & rnode_379to380_bb3__40_i295_0_valid_out_NO_SHIFT_REG & rnode_379to380_bb3_or76_i290_0_valid_out_NO_SHIFT_REG);
assign local_bb3_conv_i_i[63:32] = 32'h0;
assign local_bb3_conv_i_i[31:0] = ((local_bb3_or_i205 & 32'hFFFFFF) | 32'h800000);
assign local_bb3_shr2_i_valid_out = 1'b1;
assign local_bb3_xor_i195_valid_out = 1'b1;
assign local_bb3_and6_i_valid_out_1 = 1'b1;
assign local_bb3_conv1_i_i_valid_out = 1'b1;
assign local_bb3_var__u62_valid_out_1 = 1'b1;
assign local_bb3_shr_i193_valid_out = 1'b1;
assign local_bb3_and5_i_valid_out_1 = 1'b1;
assign local_bb3_conv_i_i_valid_out = 1'b1;
assign rnode_379to380_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_378to380_bb3_or581_i282_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_378to380_bb3_or581_i282_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_378to380_bb3_cmp68_i285_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_378to380_bb3_cmp71_not_i302_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3__40_i295_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_379to380_bb3_or76_i290_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_380to381_bb3_shr2_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr2_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_shr2_i_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr2_i_0_reg_381_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_shr2_i_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr2_i_0_valid_out_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr2_i_0_stall_in_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr2_i_0_stall_out_reg_381_NO_SHIFT_REG;

acl_data_fifo rnode_380to381_bb3_shr2_i_0_reg_381_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_380to381_bb3_shr2_i_0_reg_381_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_380to381_bb3_shr2_i_0_stall_in_reg_381_NO_SHIFT_REG),
	.valid_out(rnode_380to381_bb3_shr2_i_0_valid_out_reg_381_NO_SHIFT_REG),
	.stall_out(rnode_380to381_bb3_shr2_i_0_stall_out_reg_381_NO_SHIFT_REG),
	.data_in((local_bb3_shr2_i & 32'h1FF)),
	.data_out(rnode_380to381_bb3_shr2_i_0_reg_381_NO_SHIFT_REG)
);

defparam rnode_380to381_bb3_shr2_i_0_reg_381_fifo.DEPTH = 1;
defparam rnode_380to381_bb3_shr2_i_0_reg_381_fifo.DATA_WIDTH = 32;
defparam rnode_380to381_bb3_shr2_i_0_reg_381_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_380to381_bb3_shr2_i_0_reg_381_fifo.IMPL = "shift_reg";

assign rnode_380to381_bb3_shr2_i_0_reg_381_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr2_i_stall_in = 1'b0;
assign rnode_380to381_bb3_shr2_i_0_NO_SHIFT_REG = rnode_380to381_bb3_shr2_i_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_shr2_i_0_stall_in_reg_381_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_shr2_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_380to381_bb3_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_380to381_bb3_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_xor_i195_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_xor_i195_0_reg_381_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_xor_i195_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_xor_i195_0_valid_out_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_xor_i195_0_stall_in_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_xor_i195_0_stall_out_reg_381_NO_SHIFT_REG;

acl_data_fifo rnode_380to381_bb3_xor_i195_0_reg_381_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_380to381_bb3_xor_i195_0_reg_381_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_380to381_bb3_xor_i195_0_stall_in_reg_381_NO_SHIFT_REG),
	.valid_out(rnode_380to381_bb3_xor_i195_0_valid_out_reg_381_NO_SHIFT_REG),
	.stall_out(rnode_380to381_bb3_xor_i195_0_stall_out_reg_381_NO_SHIFT_REG),
	.data_in(local_bb3_xor_i195),
	.data_out(rnode_380to381_bb3_xor_i195_0_reg_381_NO_SHIFT_REG)
);

defparam rnode_380to381_bb3_xor_i195_0_reg_381_fifo.DEPTH = 1;
defparam rnode_380to381_bb3_xor_i195_0_reg_381_fifo.DATA_WIDTH = 32;
defparam rnode_380to381_bb3_xor_i195_0_reg_381_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_380to381_bb3_xor_i195_0_reg_381_fifo.IMPL = "shift_reg";

assign rnode_380to381_bb3_xor_i195_0_reg_381_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_xor_i195_stall_in = 1'b0;
assign rnode_380to381_bb3_xor_i195_0_NO_SHIFT_REG = rnode_380to381_bb3_xor_i195_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_xor_i195_0_stall_in_reg_381_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_380to381_bb3_and6_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_and6_i_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_and6_i_1_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_and6_i_2_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_reg_381_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_and6_i_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_valid_out_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_stall_in_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and6_i_0_stall_out_reg_381_NO_SHIFT_REG;

acl_data_fifo rnode_380to381_bb3_and6_i_0_reg_381_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_380to381_bb3_and6_i_0_reg_381_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_380to381_bb3_and6_i_0_stall_in_0_reg_381_NO_SHIFT_REG),
	.valid_out(rnode_380to381_bb3_and6_i_0_valid_out_0_reg_381_NO_SHIFT_REG),
	.stall_out(rnode_380to381_bb3_and6_i_0_stall_out_reg_381_NO_SHIFT_REG),
	.data_in((local_bb3_and6_i & 32'h7FFFFF)),
	.data_out(rnode_380to381_bb3_and6_i_0_reg_381_NO_SHIFT_REG)
);

defparam rnode_380to381_bb3_and6_i_0_reg_381_fifo.DEPTH = 1;
defparam rnode_380to381_bb3_and6_i_0_reg_381_fifo.DATA_WIDTH = 32;
defparam rnode_380to381_bb3_and6_i_0_reg_381_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_380to381_bb3_and6_i_0_reg_381_fifo.IMPL = "shift_reg";

assign rnode_380to381_bb3_and6_i_0_reg_381_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and6_i_stall_in_1 = 1'b0;
assign rnode_380to381_bb3_and6_i_0_stall_in_0_reg_381_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_and6_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_380to381_bb3_and6_i_0_NO_SHIFT_REG = rnode_380to381_bb3_and6_i_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_and6_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_380to381_bb3_and6_i_1_NO_SHIFT_REG = rnode_380to381_bb3_and6_i_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_and6_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_380to381_bb3_and6_i_2_NO_SHIFT_REG = rnode_380to381_bb3_and6_i_0_reg_381_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_380to381_bb3_var__u62_0_valid_out_NO_SHIFT_REG;
 logic rnode_380to381_bb3_var__u62_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_var__u62_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_var__u62_0_reg_381_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_var__u62_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_var__u62_0_valid_out_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_var__u62_0_stall_in_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_var__u62_0_stall_out_reg_381_NO_SHIFT_REG;

acl_data_fifo rnode_380to381_bb3_var__u62_0_reg_381_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_380to381_bb3_var__u62_0_reg_381_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_380to381_bb3_var__u62_0_stall_in_reg_381_NO_SHIFT_REG),
	.valid_out(rnode_380to381_bb3_var__u62_0_valid_out_reg_381_NO_SHIFT_REG),
	.stall_out(rnode_380to381_bb3_var__u62_0_stall_out_reg_381_NO_SHIFT_REG),
	.data_in(local_bb3_var__u62),
	.data_out(rnode_380to381_bb3_var__u62_0_reg_381_NO_SHIFT_REG)
);

defparam rnode_380to381_bb3_var__u62_0_reg_381_fifo.DEPTH = 1;
defparam rnode_380to381_bb3_var__u62_0_reg_381_fifo.DATA_WIDTH = 32;
defparam rnode_380to381_bb3_var__u62_0_reg_381_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_380to381_bb3_var__u62_0_reg_381_fifo.IMPL = "shift_reg";

assign rnode_380to381_bb3_var__u62_0_reg_381_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u62_stall_in_1 = 1'b0;
assign rnode_380to381_bb3_var__u62_0_NO_SHIFT_REG = rnode_380to381_bb3_var__u62_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_var__u62_0_stall_in_reg_381_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_var__u62_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_380to381_bb3_shr_i193_0_valid_out_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr_i193_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_shr_i193_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr_i193_0_reg_381_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_shr_i193_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr_i193_0_valid_out_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr_i193_0_stall_in_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_shr_i193_0_stall_out_reg_381_NO_SHIFT_REG;

acl_data_fifo rnode_380to381_bb3_shr_i193_0_reg_381_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_380to381_bb3_shr_i193_0_reg_381_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_380to381_bb3_shr_i193_0_stall_in_reg_381_NO_SHIFT_REG),
	.valid_out(rnode_380to381_bb3_shr_i193_0_valid_out_reg_381_NO_SHIFT_REG),
	.stall_out(rnode_380to381_bb3_shr_i193_0_stall_out_reg_381_NO_SHIFT_REG),
	.data_in((local_bb3_shr_i193 & 32'h1FF)),
	.data_out(rnode_380to381_bb3_shr_i193_0_reg_381_NO_SHIFT_REG)
);

defparam rnode_380to381_bb3_shr_i193_0_reg_381_fifo.DEPTH = 1;
defparam rnode_380to381_bb3_shr_i193_0_reg_381_fifo.DATA_WIDTH = 32;
defparam rnode_380to381_bb3_shr_i193_0_reg_381_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_380to381_bb3_shr_i193_0_reg_381_fifo.IMPL = "shift_reg";

assign rnode_380to381_bb3_shr_i193_0_reg_381_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr_i193_stall_in = 1'b0;
assign rnode_380to381_bb3_shr_i193_0_NO_SHIFT_REG = rnode_380to381_bb3_shr_i193_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_shr_i193_0_stall_in_reg_381_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_shr_i193_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_380to381_bb3_and5_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and5_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_and5_i_0_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and5_i_0_reg_381_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_380to381_bb3_and5_i_0_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and5_i_0_valid_out_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and5_i_0_stall_in_reg_381_NO_SHIFT_REG;
 logic rnode_380to381_bb3_and5_i_0_stall_out_reg_381_NO_SHIFT_REG;

acl_data_fifo rnode_380to381_bb3_and5_i_0_reg_381_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_380to381_bb3_and5_i_0_reg_381_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_380to381_bb3_and5_i_0_stall_in_reg_381_NO_SHIFT_REG),
	.valid_out(rnode_380to381_bb3_and5_i_0_valid_out_reg_381_NO_SHIFT_REG),
	.stall_out(rnode_380to381_bb3_and5_i_0_stall_out_reg_381_NO_SHIFT_REG),
	.data_in((local_bb3_and5_i & 32'h7FFFFF)),
	.data_out(rnode_380to381_bb3_and5_i_0_reg_381_NO_SHIFT_REG)
);

defparam rnode_380to381_bb3_and5_i_0_reg_381_fifo.DEPTH = 1;
defparam rnode_380to381_bb3_and5_i_0_reg_381_fifo.DATA_WIDTH = 32;
defparam rnode_380to381_bb3_and5_i_0_reg_381_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_380to381_bb3_and5_i_0_reg_381_fifo.IMPL = "shift_reg";

assign rnode_380to381_bb3_and5_i_0_reg_381_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and5_i_stall_in_1 = 1'b0;
assign rnode_380to381_bb3_and5_i_0_NO_SHIFT_REG = rnode_380to381_bb3_and5_i_0_reg_381_NO_SHIFT_REG;
assign rnode_380to381_bb3_and5_i_0_stall_in_reg_381_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_and5_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb3_mul_i_i_inputs_ready;
 reg local_bb3_mul_i_i_valid_out_0_NO_SHIFT_REG;
wire local_bb3_mul_i_i_stall_in_0;
 reg local_bb3_mul_i_i_valid_out_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i_stall_in_1;
wire local_bb3_mul_i_i_output_regs_ready;
wire [63:0] local_bb3_mul_i_i;
 reg local_bb3_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_mul_i_i_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_mul_i_i_causedstall;

acl_int_mult int_module_local_bb3_mul_i_i (
	.clock(clock),
	.dataa(((local_bb3_conv1_i_i & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb3_conv_i_i & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb3_mul_i_i_output_regs_ready),
	.result(local_bb3_mul_i_i)
);

defparam int_module_local_bb3_mul_i_i.INPUT1_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i.INPUT2_WIDTH = 24;
defparam int_module_local_bb3_mul_i_i.OUTPUT_WIDTH = 64;
defparam int_module_local_bb3_mul_i_i.LATENCY = 3;
defparam int_module_local_bb3_mul_i_i.SIGNED = 0;

assign local_bb3_mul_i_i_inputs_ready = 1'b1;
assign local_bb3_mul_i_i_output_regs_ready = 1'b1;
assign local_bb3_conv1_i_i_stall_in = 1'b0;
assign local_bb3_conv_i_i_stall_in = 1'b0;
assign local_bb3_mul_i_i_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i_output_regs_ready)
		begin
			local_bb3_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= local_bb3_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul_i_i_output_regs_ready)
		begin
			local_bb3_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_mul_i_i_stall_in_0))
			begin
				local_bb3_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_mul_i_i_stall_in_1))
			begin
				local_bb3_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_and3_i_stall_local;
wire [31:0] local_bb3_and3_i;

assign local_bb3_and3_i = ((rnode_380to381_bb3_shr2_i_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_381to384_bb3_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_381to384_bb3_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_381to384_bb3_xor_i195_0_NO_SHIFT_REG;
 logic rnode_381to384_bb3_xor_i195_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_381to384_bb3_xor_i195_0_reg_384_NO_SHIFT_REG;
 logic rnode_381to384_bb3_xor_i195_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_381to384_bb3_xor_i195_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_381to384_bb3_xor_i195_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_381to384_bb3_xor_i195_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to384_bb3_xor_i195_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to384_bb3_xor_i195_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_381to384_bb3_xor_i195_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_381to384_bb3_xor_i195_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(rnode_380to381_bb3_xor_i195_0_NO_SHIFT_REG),
	.data_out(rnode_381to384_bb3_xor_i195_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_381to384_bb3_xor_i195_0_reg_384_fifo.DEPTH = 3;
defparam rnode_381to384_bb3_xor_i195_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_381to384_bb3_xor_i195_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to384_bb3_xor_i195_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_381to384_bb3_xor_i195_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_380to381_bb3_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_381to384_bb3_xor_i195_0_NO_SHIFT_REG = rnode_381to384_bb3_xor_i195_0_reg_384_NO_SHIFT_REG;
assign rnode_381to384_bb3_xor_i195_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_381to384_bb3_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_i_stall_local;
wire local_bb3_lnot17_i;

assign local_bb3_lnot17_i = ((rnode_380to381_bb3_and6_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u64_stall_local;
wire [31:0] local_bb3_var__u64;

assign local_bb3_var__u64 = rnode_380to381_bb3_var__u62_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_and_i194_stall_local;
wire [31:0] local_bb3_and_i194;

assign local_bb3_and_i194 = ((rnode_380to381_bb3_shr_i193_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_i_stall_local;
wire local_bb3_lnot14_i;

assign local_bb3_lnot14_i = ((rnode_380to381_bb3_and5_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_conv3_i_i_stall_local;
wire [31:0] local_bb3_conv3_i_i;
wire [63:0] local_bb3_conv3_i_i$ps;

assign local_bb3_conv3_i_i$ps = (local_bb3_mul_i_i & 64'hFFFFFFFFFFFF);
assign local_bb3_conv3_i_i = local_bb3_conv3_i_i$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_var__u65_stall_local;
wire [63:0] local_bb3_var__u65;

assign local_bb3_var__u65 = ((local_bb3_mul_i_i & 64'hFFFFFFFFFFFF) >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot8_i_stall_local;
wire local_bb3_lnot8_i;

assign local_bb3_lnot8_i = ((local_bb3_and3_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_i_stall_local;
wire local_bb3_cmp11_i;

assign local_bb3_cmp11_i = ((local_bb3_and3_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u66_stall_local;
wire [31:0] local_bb3_var__u66;

assign local_bb3_var__u66 = ((local_bb3_and3_i & 32'hFF) | (rnode_380to381_bb3_and6_i_1_NO_SHIFT_REG & 32'h7FFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_xor_i195_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_xor_i195_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_xor_i195_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_xor_i195_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_xor_i195_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_xor_i195_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_xor_i195_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_xor_i195_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_xor_i195_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_xor_i195_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_xor_i195_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(rnode_381to384_bb3_xor_i195_0_NO_SHIFT_REG),
	.data_out(rnode_384to385_bb3_xor_i195_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_xor_i195_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_xor_i195_0_reg_385_fifo.DATA_WIDTH = 32;
defparam rnode_384to385_bb3_xor_i195_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_xor_i195_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_xor_i195_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_381to384_bb3_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_xor_i195_0_NO_SHIFT_REG = rnode_384to385_bb3_xor_i195_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_xor_i195_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_lnot17_not_i_stall_local;
wire local_bb3_lnot17_not_i;

assign local_bb3_lnot17_not_i = (local_bb3_lnot17_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_and_i_stall_local;
wire [31:0] local_bb3_and_i;

assign local_bb3_and_i = (local_bb3_var__u64 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and10_i_stall_local;
wire [31:0] local_bb3_and10_i;

assign local_bb3_and10_i = (local_bb3_var__u64 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_i196_stall_local;
wire local_bb3_lnot_i196;

assign local_bb3_lnot_i196 = ((local_bb3_and_i194 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i197_stall_local;
wire local_bb3_cmp_i197;

assign local_bb3_cmp_i197 = ((local_bb3_and_i194 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u67_stall_local;
wire [31:0] local_bb3_var__u67;

assign local_bb3_var__u67 = ((rnode_380to381_bb3_and6_i_2_NO_SHIFT_REG & 32'h7FFFFF) | (local_bb3_and_i194 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_add_i206_stall_local;
wire [31:0] local_bb3_add_i206;

assign local_bb3_add_i206 = ((local_bb3_and3_i & 32'hFF) + (local_bb3_and_i194 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot14_not_i_stall_local;
wire local_bb3_lnot14_not_i;

assign local_bb3_lnot14_not_i = (local_bb3_lnot14_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i16_i_stall_local;
wire [31:0] local_bb3_shr_i16_i;

assign local_bb3_shr_i16_i = (local_bb3_conv3_i_i >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i18_i_stall_local;
wire [31:0] local_bb3_shl1_i18_i;

assign local_bb3_shl1_i18_i = (local_bb3_conv3_i_i << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u68_stall_local;
wire [31:0] local_bb3_var__u68;

assign local_bb3_var__u68 = (local_bb3_conv3_i_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shl1_i_i_stall_local;
wire [31:0] local_bb3_shl1_i_i;

assign local_bb3_shl1_i_i = (local_bb3_conv3_i_i << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb3__tr_i_stall_local;
wire [31:0] local_bb3__tr_i;
wire [63:0] local_bb3__tr_i$ps;

assign local_bb3__tr_i$ps = (local_bb3_var__u65 & 64'hFFFFFF);
assign local_bb3__tr_i = local_bb3__tr_i$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge8_demorgan_i_stall_local;
wire local_bb3_brmerge8_demorgan_i;

assign local_bb3_brmerge8_demorgan_i = (local_bb3_cmp11_i & local_bb3_lnot17_i);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp11_not_i_stall_local;
wire local_bb3_cmp11_not_i;

assign local_bb3_cmp11_not_i = (local_bb3_cmp11_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u69_stall_local;
wire local_bb3_var__u69;

assign local_bb3_var__u69 = ((local_bb3_var__u66 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and4_i_stall_local;
wire [31:0] local_bb3_and4_i;

assign local_bb3_and4_i = (rnode_384to385_bb3_xor_i195_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i1_stall_local;
wire [31:0] local_bb3_shr_i1;

assign local_bb3_shr_i1 = ((local_bb3_and_i & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp13_i_stall_local;
wire local_bb3_cmp13_i;

assign local_bb3_cmp13_i = ((local_bb3_and10_i & 32'hFFFF) > (local_bb3_and12_i & 32'hFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_0_i212_stall_local;
wire local_bb3_reduction_0_i212;

assign local_bb3_reduction_0_i212 = (local_bb3_lnot_i196 | local_bb3_lnot8_i);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u70_stall_local;
wire local_bb3_var__u70;

assign local_bb3_var__u70 = (local_bb3_cmp_i197 | local_bb3_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u71_stall_local;
wire local_bb3_var__u71;

assign local_bb3_var__u71 = ((local_bb3_var__u67 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__28_i203_stall_local;
wire local_bb3__28_i203;

assign local_bb3__28_i203 = (local_bb3_cmp_i197 & local_bb3_lnot14_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i_i207_stall_local;
wire [31:0] local_bb3_shr_i_i207;

assign local_bb3_shr_i_i207 = ((local_bb3_var__u68 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i15_i_stall_local;
wire [31:0] local_bb3_shl_i15_i;

assign local_bb3_shl_i15_i = ((local_bb3__tr_i & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb3_and48_i_stall_local;
wire [31:0] local_bb3_and48_i;

assign local_bb3_and48_i = ((local_bb3__tr_i & 32'hFFFFFF) & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge10_demorgan_i_stall_local;
wire local_bb3_brmerge10_demorgan_i;

assign local_bb3_brmerge10_demorgan_i = (local_bb3_brmerge8_demorgan_i & local_bb3_lnot_i196);

// This section implements an unregistered operation.
// 
wire local_bb3__mux9_mux_i_stall_local;
wire local_bb3__mux9_mux_i;

assign local_bb3__mux9_mux_i = (local_bb3_brmerge8_demorgan_i ^ local_bb3_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge3_i_stall_local;
wire local_bb3_brmerge3_i;

assign local_bb3_brmerge3_i = (local_bb3_var__u69 | local_bb3_cmp11_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_i_stall_local;
wire local_bb3__mux_mux_i;

assign local_bb3__mux_mux_i = (local_bb3_var__u69 | local_bb3_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb3__not_i_stall_local;
wire local_bb3__not_i;

assign local_bb3__not_i = (local_bb3_var__u69 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i3_stall_local;
wire local_bb3_cmp_i3;

assign local_bb3_cmp_i3 = ((local_bb3_shr_i1 & 32'h7FFF) > (local_bb3_shr3_i & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp8_i_stall_local;
wire local_bb3_cmp8_i;

assign local_bb3_cmp8_i = ((local_bb3_shr_i1 & 32'h7FFF) == (local_bb3_shr3_i & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb3_or_i17_i_stall_local;
wire [31:0] local_bb3_or_i17_i;

assign local_bb3_or_i17_i = ((local_bb3_shl_i15_i & 32'hFFFF00) | (local_bb3_shr_i16_i & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool49_i_stall_local;
wire local_bb3_tobool49_i;

assign local_bb3_tobool49_i = ((local_bb3_and48_i & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__26_demorgan_i_stall_local;
wire local_bb3__26_demorgan_i;

assign local_bb3__26_demorgan_i = (local_bb3_cmp_i197 | local_bb3_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge5_i_stall_local;
wire local_bb3_brmerge5_i;

assign local_bb3_brmerge5_i = (local_bb3_brmerge3_i | local_bb3_lnot17_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_3_i198_stall_local;
wire local_bb3_reduction_3_i198;

assign local_bb3_reduction_3_i198 = (local_bb3_cmp11_i & local_bb3__not_i);

// This section implements an unregistered operation.
// 
wire local_bb3___i4_stall_local;
wire local_bb3___i4;

assign local_bb3___i4 = (local_bb3_cmp8_i & local_bb3_cmp13_i);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i_i_stall_local;
wire [31:0] local_bb3_shl_i_i;

assign local_bb3_shl_i_i = ((local_bb3_or_i17_i & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__mux_mux_mux_i_stall_local;
wire local_bb3__mux_mux_mux_i;

assign local_bb3__mux_mux_mux_i = (local_bb3_brmerge5_i & local_bb3__mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_5_i199_stall_local;
wire local_bb3_reduction_5_i199;

assign local_bb3_reduction_5_i199 = (local_bb3_lnot14_i & local_bb3_reduction_3_i198);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u21_valid_out_2;
wire local_bb3_var__u21_stall_in_2;
wire local_bb3__21_i_valid_out;
wire local_bb3__21_i_stall_in;
wire local_bb3_var__u64_valid_out_2;
wire local_bb3_var__u64_stall_in_2;
wire local_bb3__21_i_inputs_ready;
wire local_bb3__21_i_stall_local;
wire local_bb3__21_i;

assign local_bb3__21_i_inputs_ready = (rnode_380to381_bb3_c0_ene6_0_valid_out_0_NO_SHIFT_REG & rnode_380to381_bb3_var__u62_0_valid_out_NO_SHIFT_REG);
assign local_bb3__21_i = (local_bb3_cmp_i3 | local_bb3___i4);
assign local_bb3_var__u21_valid_out_2 = 1'b1;
assign local_bb3__21_i_valid_out = 1'b1;
assign local_bb3_var__u64_valid_out_2 = 1'b1;
assign rnode_380to381_bb3_c0_ene6_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_var__u62_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_or_i_i208_stall_local;
wire [31:0] local_bb3_or_i_i208;

assign local_bb3_or_i_i208 = ((local_bb3_shl_i_i & 32'h1FFFFFE) | (local_bb3_shr_i_i207 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_6_i200_stall_local;
wire local_bb3_reduction_6_i200;

assign local_bb3_reduction_6_i200 = (local_bb3_var__u71 & local_bb3_reduction_5_i199);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_381to382_bb3_var__u21_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u21_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_var__u21_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u21_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u21_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_var__u21_1_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u21_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_var__u21_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u21_0_valid_out_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u21_0_stall_in_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u21_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_381to382_bb3_var__u21_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to382_bb3_var__u21_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to382_bb3_var__u21_0_stall_in_0_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_381to382_bb3_var__u21_0_valid_out_0_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_381to382_bb3_var__u21_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(local_bb3_var__u21),
	.data_out(rnode_381to382_bb3_var__u21_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_381to382_bb3_var__u21_0_reg_382_fifo.DEPTH = 1;
defparam rnode_381to382_bb3_var__u21_0_reg_382_fifo.DATA_WIDTH = 32;
defparam rnode_381to382_bb3_var__u21_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to382_bb3_var__u21_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_381to382_bb3_var__u21_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u21_stall_in_2 = 1'b0;
assign rnode_381to382_bb3_var__u21_0_stall_in_0_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_var__u21_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3_var__u21_0_NO_SHIFT_REG = rnode_381to382_bb3_var__u21_0_reg_382_NO_SHIFT_REG;
assign rnode_381to382_bb3_var__u21_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3_var__u21_1_NO_SHIFT_REG = rnode_381to382_bb3_var__u21_0_reg_382_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_381to382_bb3__21_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_1_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_valid_out_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_stall_in_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3__21_i_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_381to382_bb3__21_i_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to382_bb3__21_i_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to382_bb3__21_i_0_stall_in_0_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_381to382_bb3__21_i_0_valid_out_0_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_381to382_bb3__21_i_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(local_bb3__21_i),
	.data_out(rnode_381to382_bb3__21_i_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_381to382_bb3__21_i_0_reg_382_fifo.DEPTH = 1;
defparam rnode_381to382_bb3__21_i_0_reg_382_fifo.DATA_WIDTH = 1;
defparam rnode_381to382_bb3__21_i_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to382_bb3__21_i_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_381to382_bb3__21_i_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__21_i_stall_in = 1'b0;
assign rnode_381to382_bb3__21_i_0_stall_in_0_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3__21_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3__21_i_0_NO_SHIFT_REG = rnode_381to382_bb3__21_i_0_reg_382_NO_SHIFT_REG;
assign rnode_381to382_bb3__21_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3__21_i_1_NO_SHIFT_REG = rnode_381to382_bb3__21_i_0_reg_382_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_381to382_bb3_var__u64_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u64_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_var__u64_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u64_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u64_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_var__u64_1_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u64_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_381to382_bb3_var__u64_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u64_0_valid_out_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u64_0_stall_in_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u64_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_381to382_bb3_var__u64_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to382_bb3_var__u64_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to382_bb3_var__u64_0_stall_in_0_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_381to382_bb3_var__u64_0_valid_out_0_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_381to382_bb3_var__u64_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(local_bb3_var__u64),
	.data_out(rnode_381to382_bb3_var__u64_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_381to382_bb3_var__u64_0_reg_382_fifo.DEPTH = 1;
defparam rnode_381to382_bb3_var__u64_0_reg_382_fifo.DATA_WIDTH = 32;
defparam rnode_381to382_bb3_var__u64_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to382_bb3_var__u64_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_381to382_bb3_var__u64_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u64_stall_in_2 = 1'b0;
assign rnode_381to382_bb3_var__u64_0_stall_in_0_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_var__u64_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3_var__u64_0_NO_SHIFT_REG = rnode_381to382_bb3_var__u64_0_reg_382_NO_SHIFT_REG;
assign rnode_381to382_bb3_var__u64_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3_var__u64_1_NO_SHIFT_REG = rnode_381to382_bb3_var__u64_0_reg_382_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__24_i201_stall_local;
wire local_bb3__24_i201;

assign local_bb3__24_i201 = (local_bb3_cmp_i197 ? local_bb3_reduction_6_i200 : local_bb3_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb3__22_i_stall_local;
wire [31:0] local_bb3__22_i;

assign local_bb3__22_i = (rnode_381to382_bb3__21_i_0_NO_SHIFT_REG ? rnode_381to382_bb3_var__u21_0_NO_SHIFT_REG : rnode_381to382_bb3_var__u64_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3__23_i_stall_local;
wire [31:0] local_bb3__23_i;

assign local_bb3__23_i = (rnode_381to382_bb3__21_i_1_NO_SHIFT_REG ? rnode_381to382_bb3_var__u64_1_NO_SHIFT_REG : rnode_381to382_bb3_var__u21_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3__25_i_stall_local;
wire local_bb3__25_i;

assign local_bb3__25_i = (local_bb3__24_i201 ? local_bb3_lnot14_i : local_bb3__mux_mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb3_shr18_i_stall_local;
wire [31:0] local_bb3_shr18_i;

assign local_bb3_shr18_i = (local_bb3__22_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shr16_i_stall_local;
wire [31:0] local_bb3_shr16_i;

assign local_bb3_shr16_i = (local_bb3__23_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3__27_i202_stall_local;
wire local_bb3__27_i202;

assign local_bb3__27_i202 = (local_bb3__26_demorgan_i ? local_bb3__25_i : local_bb3__mux9_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb3_and19_i_stall_local;
wire [31:0] local_bb3_and19_i;

assign local_bb3_and19_i = ((local_bb3_shr18_i & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_sub_i_stall_local;
wire [31:0] local_bb3_sub_i;

assign local_bb3_sub_i = ((local_bb3_shr16_i & 32'h1FF) - (local_bb3_shr18_i & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb3_add_i206_valid_out;
wire local_bb3_add_i206_stall_in;
wire local_bb3_reduction_0_i212_valid_out;
wire local_bb3_reduction_0_i212_stall_in;
wire local_bb3_var__u70_valid_out;
wire local_bb3_var__u70_stall_in;
wire local_bb3__29_i204_valid_out;
wire local_bb3__29_i204_stall_in;
wire local_bb3__29_i204_inputs_ready;
wire local_bb3__29_i204_stall_local;
wire local_bb3__29_i204;

assign local_bb3__29_i204_inputs_ready = (rnode_380to381_bb3_shr2_i_0_valid_out_NO_SHIFT_REG & rnode_380to381_bb3_and6_i_0_valid_out_1_NO_SHIFT_REG & rnode_380to381_bb3_and6_i_0_valid_out_0_NO_SHIFT_REG & rnode_380to381_bb3_and6_i_0_valid_out_2_NO_SHIFT_REG & rnode_380to381_bb3_shr_i193_0_valid_out_NO_SHIFT_REG & rnode_380to381_bb3_and5_i_0_valid_out_NO_SHIFT_REG);
assign local_bb3__29_i204 = (local_bb3__28_i203 | local_bb3__27_i202);
assign local_bb3_add_i206_valid_out = 1'b1;
assign local_bb3_reduction_0_i212_valid_out = 1'b1;
assign local_bb3_var__u70_valid_out = 1'b1;
assign local_bb3__29_i204_valid_out = 1'b1;
assign rnode_380to381_bb3_shr2_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_and6_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_and6_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_and6_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_shr_i193_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_380to381_bb3_and5_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_lnot23_i_stall_local;
wire local_bb3_lnot23_i;

assign local_bb3_lnot23_i = ((local_bb3_and19_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp27_i_stall_local;
wire local_bb3_cmp27_i;

assign local_bb3_cmp27_i = ((local_bb3_and19_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and68_i_stall_local;
wire [31:0] local_bb3_and68_i;

assign local_bb3_and68_i = (local_bb3_sub_i & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_381to383_bb3_add_i206_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_381to383_bb3_add_i206_0_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_381to383_bb3_add_i206_1_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_381to383_bb3_add_i206_2_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_reg_383_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_381to383_bb3_add_i206_0_reg_383_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_valid_out_0_reg_383_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_stall_in_0_reg_383_NO_SHIFT_REG;
 logic rnode_381to383_bb3_add_i206_0_stall_out_reg_383_NO_SHIFT_REG;

acl_data_fifo rnode_381to383_bb3_add_i206_0_reg_383_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to383_bb3_add_i206_0_reg_383_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to383_bb3_add_i206_0_stall_in_0_reg_383_NO_SHIFT_REG),
	.valid_out(rnode_381to383_bb3_add_i206_0_valid_out_0_reg_383_NO_SHIFT_REG),
	.stall_out(rnode_381to383_bb3_add_i206_0_stall_out_reg_383_NO_SHIFT_REG),
	.data_in((local_bb3_add_i206 & 32'h1FF)),
	.data_out(rnode_381to383_bb3_add_i206_0_reg_383_NO_SHIFT_REG)
);

defparam rnode_381to383_bb3_add_i206_0_reg_383_fifo.DEPTH = 2;
defparam rnode_381to383_bb3_add_i206_0_reg_383_fifo.DATA_WIDTH = 32;
defparam rnode_381to383_bb3_add_i206_0_reg_383_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to383_bb3_add_i206_0_reg_383_fifo.IMPL = "shift_reg";

assign rnode_381to383_bb3_add_i206_0_reg_383_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add_i206_stall_in = 1'b0;
assign rnode_381to383_bb3_add_i206_0_stall_in_0_reg_383_NO_SHIFT_REG = 1'b0;
assign rnode_381to383_bb3_add_i206_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_381to383_bb3_add_i206_0_NO_SHIFT_REG = rnode_381to383_bb3_add_i206_0_reg_383_NO_SHIFT_REG;
assign rnode_381to383_bb3_add_i206_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_381to383_bb3_add_i206_1_NO_SHIFT_REG = rnode_381to383_bb3_add_i206_0_reg_383_NO_SHIFT_REG;
assign rnode_381to383_bb3_add_i206_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_381to383_bb3_add_i206_2_NO_SHIFT_REG = rnode_381to383_bb3_add_i206_0_reg_383_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_381to382_bb3_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_381to382_bb3_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_381to382_bb3_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3_reduction_0_i212_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic rnode_381to382_bb3_reduction_0_i212_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_reduction_0_i212_0_valid_out_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_reduction_0_i212_0_stall_in_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_reduction_0_i212_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_381to382_bb3_reduction_0_i212_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to382_bb3_reduction_0_i212_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to382_bb3_reduction_0_i212_0_stall_in_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_381to382_bb3_reduction_0_i212_0_valid_out_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_381to382_bb3_reduction_0_i212_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(local_bb3_reduction_0_i212),
	.data_out(rnode_381to382_bb3_reduction_0_i212_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_381to382_bb3_reduction_0_i212_0_reg_382_fifo.DEPTH = 1;
defparam rnode_381to382_bb3_reduction_0_i212_0_reg_382_fifo.DATA_WIDTH = 1;
defparam rnode_381to382_bb3_reduction_0_i212_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to382_bb3_reduction_0_i212_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_381to382_bb3_reduction_0_i212_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_reduction_0_i212_stall_in = 1'b0;
assign rnode_381to382_bb3_reduction_0_i212_0_NO_SHIFT_REG = rnode_381to382_bb3_reduction_0_i212_0_reg_382_NO_SHIFT_REG;
assign rnode_381to382_bb3_reduction_0_i212_0_stall_in_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_381to382_bb3_var__u70_0_valid_out_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u70_0_stall_in_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u70_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u70_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u70_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u70_0_valid_out_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u70_0_stall_in_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3_var__u70_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_381to382_bb3_var__u70_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to382_bb3_var__u70_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to382_bb3_var__u70_0_stall_in_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_381to382_bb3_var__u70_0_valid_out_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_381to382_bb3_var__u70_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(local_bb3_var__u70),
	.data_out(rnode_381to382_bb3_var__u70_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_381to382_bb3_var__u70_0_reg_382_fifo.DEPTH = 1;
defparam rnode_381to382_bb3_var__u70_0_reg_382_fifo.DATA_WIDTH = 1;
defparam rnode_381to382_bb3_var__u70_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to382_bb3_var__u70_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_381to382_bb3_var__u70_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u70_stall_in = 1'b0;
assign rnode_381to382_bb3_var__u70_0_NO_SHIFT_REG = rnode_381to382_bb3_var__u70_0_reg_382_NO_SHIFT_REG;
assign rnode_381to382_bb3_var__u70_0_stall_in_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_var__u70_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_381to382_bb3__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_381to382_bb3__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_381to382_bb3__29_i204_0_NO_SHIFT_REG;
 logic rnode_381to382_bb3__29_i204_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic rnode_381to382_bb3__29_i204_0_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3__29_i204_0_valid_out_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3__29_i204_0_stall_in_reg_382_NO_SHIFT_REG;
 logic rnode_381to382_bb3__29_i204_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_381to382_bb3__29_i204_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_381to382_bb3__29_i204_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_381to382_bb3__29_i204_0_stall_in_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_381to382_bb3__29_i204_0_valid_out_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_381to382_bb3__29_i204_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(local_bb3__29_i204),
	.data_out(rnode_381to382_bb3__29_i204_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_381to382_bb3__29_i204_0_reg_382_fifo.DEPTH = 1;
defparam rnode_381to382_bb3__29_i204_0_reg_382_fifo.DATA_WIDTH = 1;
defparam rnode_381to382_bb3__29_i204_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_381to382_bb3__29_i204_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_381to382_bb3__29_i204_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__29_i204_stall_in = 1'b0;
assign rnode_381to382_bb3__29_i204_0_NO_SHIFT_REG = rnode_381to382_bb3__29_i204_0_reg_382_NO_SHIFT_REG;
assign rnode_381to382_bb3__29_i204_0_stall_in_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp69_i_stall_local;
wire local_bb3_cmp69_i;

assign local_bb3_cmp69_i = ((local_bb3_and68_i & 32'hFF) > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_inc_i_stall_local;
wire [31:0] local_bb3_inc_i;

assign local_bb3_inc_i = ((rnode_381to383_bb3_add_i206_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp50_not_i_stall_local;
wire local_bb3_cmp50_not_i;

assign local_bb3_cmp50_not_i = ((rnode_381to383_bb3_add_i206_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_382to384_bb3_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_382to384_bb3_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_382to384_bb3_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_382to384_bb3_reduction_0_i212_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_382to384_bb3_reduction_0_i212_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_reduction_0_i212_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_reduction_0_i212_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_reduction_0_i212_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_382to384_bb3_reduction_0_i212_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to384_bb3_reduction_0_i212_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to384_bb3_reduction_0_i212_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_382to384_bb3_reduction_0_i212_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_382to384_bb3_reduction_0_i212_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(rnode_381to382_bb3_reduction_0_i212_0_NO_SHIFT_REG),
	.data_out(rnode_382to384_bb3_reduction_0_i212_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_382to384_bb3_reduction_0_i212_0_reg_384_fifo.DEPTH = 2;
defparam rnode_382to384_bb3_reduction_0_i212_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_382to384_bb3_reduction_0_i212_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to384_bb3_reduction_0_i212_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_382to384_bb3_reduction_0_i212_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3_reduction_0_i212_0_NO_SHIFT_REG = rnode_382to384_bb3_reduction_0_i212_0_reg_384_NO_SHIFT_REG;
assign rnode_382to384_bb3_reduction_0_i212_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_382to383_bb3_var__u70_0_valid_out_NO_SHIFT_REG;
 logic rnode_382to383_bb3_var__u70_0_stall_in_NO_SHIFT_REG;
 logic rnode_382to383_bb3_var__u70_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3_var__u70_0_reg_383_inputs_ready_NO_SHIFT_REG;
 logic rnode_382to383_bb3_var__u70_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_var__u70_0_valid_out_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_var__u70_0_stall_in_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_var__u70_0_stall_out_reg_383_NO_SHIFT_REG;

acl_data_fifo rnode_382to383_bb3_var__u70_0_reg_383_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to383_bb3_var__u70_0_reg_383_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to383_bb3_var__u70_0_stall_in_reg_383_NO_SHIFT_REG),
	.valid_out(rnode_382to383_bb3_var__u70_0_valid_out_reg_383_NO_SHIFT_REG),
	.stall_out(rnode_382to383_bb3_var__u70_0_stall_out_reg_383_NO_SHIFT_REG),
	.data_in(rnode_381to382_bb3_var__u70_0_NO_SHIFT_REG),
	.data_out(rnode_382to383_bb3_var__u70_0_reg_383_NO_SHIFT_REG)
);

defparam rnode_382to383_bb3_var__u70_0_reg_383_fifo.DEPTH = 1;
defparam rnode_382to383_bb3_var__u70_0_reg_383_fifo.DATA_WIDTH = 1;
defparam rnode_382to383_bb3_var__u70_0_reg_383_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to383_bb3_var__u70_0_reg_383_fifo.IMPL = "shift_reg";

assign rnode_382to383_bb3_var__u70_0_reg_383_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3_var__u70_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_var__u70_0_NO_SHIFT_REG = rnode_382to383_bb3_var__u70_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3_var__u70_0_stall_in_reg_383_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_var__u70_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_382to384_bb3__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_382to384_bb3__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_382to384_bb3__29_i204_0_NO_SHIFT_REG;
 logic rnode_382to384_bb3__29_i204_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_382to384_bb3__29_i204_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3__29_i204_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3__29_i204_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3__29_i204_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_382to384_bb3__29_i204_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to384_bb3__29_i204_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to384_bb3__29_i204_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_382to384_bb3__29_i204_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_382to384_bb3__29_i204_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(rnode_381to382_bb3__29_i204_0_NO_SHIFT_REG),
	.data_out(rnode_382to384_bb3__29_i204_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_382to384_bb3__29_i204_0_reg_384_fifo.DEPTH = 2;
defparam rnode_382to384_bb3__29_i204_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_382to384_bb3__29_i204_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to384_bb3__29_i204_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_382to384_bb3__29_i204_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_381to382_bb3__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3__29_i204_0_NO_SHIFT_REG = rnode_382to384_bb3__29_i204_0_reg_384_NO_SHIFT_REG;
assign rnode_382to384_bb3__29_i204_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__22_i_valid_out_1;
wire local_bb3__22_i_stall_in_1;
wire local_bb3__23_i_valid_out_1;
wire local_bb3__23_i_stall_in_1;
wire local_bb3_shr16_i_valid_out_1;
wire local_bb3_shr16_i_stall_in_1;
wire local_bb3_lnot23_i_valid_out;
wire local_bb3_lnot23_i_stall_in;
wire local_bb3_cmp27_i_valid_out;
wire local_bb3_cmp27_i_stall_in;
wire local_bb3_align_0_i_valid_out;
wire local_bb3_align_0_i_stall_in;
wire local_bb3_align_0_i_inputs_ready;
wire local_bb3_align_0_i_stall_local;
wire [31:0] local_bb3_align_0_i;

assign local_bb3_align_0_i_inputs_ready = (rnode_381to382_bb3__21_i_0_valid_out_0_NO_SHIFT_REG & rnode_381to382_bb3_var__u21_0_valid_out_0_NO_SHIFT_REG & rnode_381to382_bb3_var__u64_0_valid_out_0_NO_SHIFT_REG & rnode_381to382_bb3__21_i_0_valid_out_1_NO_SHIFT_REG & rnode_381to382_bb3_var__u64_0_valid_out_1_NO_SHIFT_REG & rnode_381to382_bb3_var__u21_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_align_0_i = (local_bb3_cmp69_i ? 32'h1F : (local_bb3_and68_i & 32'hFF));
assign local_bb3__22_i_valid_out_1 = 1'b1;
assign local_bb3__23_i_valid_out_1 = 1'b1;
assign local_bb3_shr16_i_valid_out_1 = 1'b1;
assign local_bb3_lnot23_i_valid_out = 1'b1;
assign local_bb3_cmp27_i_valid_out = 1'b1;
assign local_bb3_align_0_i_valid_out = 1'b1;
assign rnode_381to382_bb3__21_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_var__u21_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_var__u64_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3__21_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_var__u64_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_381to382_bb3_var__u21_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__31_i209_stall_local;
wire local_bb3__31_i209;

assign local_bb3__31_i209 = (local_bb3_tobool49_i & local_bb3_cmp50_not_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb3_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_reduction_0_i212_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3_reduction_0_i212_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_reduction_0_i212_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_reduction_0_i212_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_reduction_0_i212_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_reduction_0_i212_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_reduction_0_i212_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_reduction_0_i212_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_reduction_0_i212_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_reduction_0_i212_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(rnode_382to384_bb3_reduction_0_i212_0_NO_SHIFT_REG),
	.data_out(rnode_384to385_bb3_reduction_0_i212_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_reduction_0_i212_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_reduction_0_i212_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3_reduction_0_i212_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_reduction_0_i212_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_reduction_0_i212_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_reduction_0_i212_0_NO_SHIFT_REG = rnode_384to385_bb3_reduction_0_i212_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_reduction_0_i212_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_var__u70_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb3_var__u70_0_stall_in_NO_SHIFT_REG;
 logic rnode_383to384_bb3_var__u70_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_var__u70_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb3_var__u70_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_var__u70_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_var__u70_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_var__u70_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_var__u70_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_var__u70_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_var__u70_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_var__u70_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_var__u70_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(rnode_382to383_bb3_var__u70_0_NO_SHIFT_REG),
	.data_out(rnode_383to384_bb3_var__u70_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_var__u70_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_var__u70_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb3_var__u70_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_var__u70_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_var__u70_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3_var__u70_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_var__u70_0_NO_SHIFT_REG = rnode_383to384_bb3_var__u70_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_var__u70_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_var__u70_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb3__29_i204_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3__29_i204_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3__29_i204_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__29_i204_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__29_i204_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__29_i204_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3__29_i204_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3__29_i204_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3__29_i204_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3__29_i204_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3__29_i204_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(rnode_382to384_bb3__29_i204_0_NO_SHIFT_REG),
	.data_out(rnode_384to385_bb3__29_i204_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3__29_i204_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3__29_i204_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3__29_i204_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3__29_i204_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3__29_i204_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3__29_i204_0_NO_SHIFT_REG = rnode_384to385_bb3__29_i204_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3__29_i204_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_382to383_bb3__22_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3__22_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3__22_i_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3__22_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_382to383_bb3__22_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3__22_i_1_NO_SHIFT_REG;
 logic rnode_382to383_bb3__22_i_0_reg_383_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3__22_i_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3__22_i_0_valid_out_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3__22_i_0_stall_in_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3__22_i_0_stall_out_reg_383_NO_SHIFT_REG;

acl_data_fifo rnode_382to383_bb3__22_i_0_reg_383_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to383_bb3__22_i_0_reg_383_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to383_bb3__22_i_0_stall_in_0_reg_383_NO_SHIFT_REG),
	.valid_out(rnode_382to383_bb3__22_i_0_valid_out_0_reg_383_NO_SHIFT_REG),
	.stall_out(rnode_382to383_bb3__22_i_0_stall_out_reg_383_NO_SHIFT_REG),
	.data_in(local_bb3__22_i),
	.data_out(rnode_382to383_bb3__22_i_0_reg_383_NO_SHIFT_REG)
);

defparam rnode_382to383_bb3__22_i_0_reg_383_fifo.DEPTH = 1;
defparam rnode_382to383_bb3__22_i_0_reg_383_fifo.DATA_WIDTH = 32;
defparam rnode_382to383_bb3__22_i_0_reg_383_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to383_bb3__22_i_0_reg_383_fifo.IMPL = "shift_reg";

assign rnode_382to383_bb3__22_i_0_reg_383_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__22_i_stall_in_1 = 1'b0;
assign rnode_382to383_bb3__22_i_0_stall_in_0_reg_383_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3__22_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3__22_i_0_NO_SHIFT_REG = rnode_382to383_bb3__22_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3__22_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3__22_i_1_NO_SHIFT_REG = rnode_382to383_bb3__22_i_0_reg_383_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_382to383_bb3__23_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3__23_i_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3__23_i_1_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3__23_i_2_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_reg_383_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3__23_i_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_valid_out_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_stall_in_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3__23_i_0_stall_out_reg_383_NO_SHIFT_REG;

acl_data_fifo rnode_382to383_bb3__23_i_0_reg_383_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to383_bb3__23_i_0_reg_383_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to383_bb3__23_i_0_stall_in_0_reg_383_NO_SHIFT_REG),
	.valid_out(rnode_382to383_bb3__23_i_0_valid_out_0_reg_383_NO_SHIFT_REG),
	.stall_out(rnode_382to383_bb3__23_i_0_stall_out_reg_383_NO_SHIFT_REG),
	.data_in(local_bb3__23_i),
	.data_out(rnode_382to383_bb3__23_i_0_reg_383_NO_SHIFT_REG)
);

defparam rnode_382to383_bb3__23_i_0_reg_383_fifo.DEPTH = 1;
defparam rnode_382to383_bb3__23_i_0_reg_383_fifo.DATA_WIDTH = 32;
defparam rnode_382to383_bb3__23_i_0_reg_383_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to383_bb3__23_i_0_reg_383_fifo.IMPL = "shift_reg";

assign rnode_382to383_bb3__23_i_0_reg_383_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__23_i_stall_in_1 = 1'b0;
assign rnode_382to383_bb3__23_i_0_stall_in_0_reg_383_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3__23_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3__23_i_0_NO_SHIFT_REG = rnode_382to383_bb3__23_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3__23_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3__23_i_1_NO_SHIFT_REG = rnode_382to383_bb3__23_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3__23_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3__23_i_2_NO_SHIFT_REG = rnode_382to383_bb3__23_i_0_reg_383_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_382to384_bb3_shr16_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_382to384_bb3_shr16_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_382to384_bb3_shr16_i_0_NO_SHIFT_REG;
 logic rnode_382to384_bb3_shr16_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_382to384_bb3_shr16_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_382to384_bb3_shr16_i_1_NO_SHIFT_REG;
 logic rnode_382to384_bb3_shr16_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_382to384_bb3_shr16_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_shr16_i_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_shr16_i_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_shr16_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_382to384_bb3_shr16_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to384_bb3_shr16_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to384_bb3_shr16_i_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_382to384_bb3_shr16_i_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_382to384_bb3_shr16_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb3_shr16_i & 32'h1FF)),
	.data_out(rnode_382to384_bb3_shr16_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_382to384_bb3_shr16_i_0_reg_384_fifo.DEPTH = 2;
defparam rnode_382to384_bb3_shr16_i_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_382to384_bb3_shr16_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to384_bb3_shr16_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_382to384_bb3_shr16_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr16_i_stall_in_1 = 1'b0;
assign rnode_382to384_bb3_shr16_i_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3_shr16_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3_shr16_i_0_NO_SHIFT_REG = rnode_382to384_bb3_shr16_i_0_reg_384_NO_SHIFT_REG;
assign rnode_382to384_bb3_shr16_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3_shr16_i_1_NO_SHIFT_REG = rnode_382to384_bb3_shr16_i_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_382to383_bb3_lnot23_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_382to383_bb3_lnot23_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_382to383_bb3_lnot23_i_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3_lnot23_i_0_reg_383_inputs_ready_NO_SHIFT_REG;
 logic rnode_382to383_bb3_lnot23_i_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_lnot23_i_0_valid_out_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_lnot23_i_0_stall_in_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_lnot23_i_0_stall_out_reg_383_NO_SHIFT_REG;

acl_data_fifo rnode_382to383_bb3_lnot23_i_0_reg_383_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to383_bb3_lnot23_i_0_reg_383_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to383_bb3_lnot23_i_0_stall_in_reg_383_NO_SHIFT_REG),
	.valid_out(rnode_382to383_bb3_lnot23_i_0_valid_out_reg_383_NO_SHIFT_REG),
	.stall_out(rnode_382to383_bb3_lnot23_i_0_stall_out_reg_383_NO_SHIFT_REG),
	.data_in(local_bb3_lnot23_i),
	.data_out(rnode_382to383_bb3_lnot23_i_0_reg_383_NO_SHIFT_REG)
);

defparam rnode_382to383_bb3_lnot23_i_0_reg_383_fifo.DEPTH = 1;
defparam rnode_382to383_bb3_lnot23_i_0_reg_383_fifo.DATA_WIDTH = 1;
defparam rnode_382to383_bb3_lnot23_i_0_reg_383_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to383_bb3_lnot23_i_0_reg_383_fifo.IMPL = "shift_reg";

assign rnode_382to383_bb3_lnot23_i_0_reg_383_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_lnot23_i_stall_in = 1'b0;
assign rnode_382to383_bb3_lnot23_i_0_NO_SHIFT_REG = rnode_382to383_bb3_lnot23_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3_lnot23_i_0_stall_in_reg_383_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_lnot23_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_382to384_bb3_cmp27_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_1_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_2_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_382to384_bb3_cmp27_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_382to384_bb3_cmp27_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to384_bb3_cmp27_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to384_bb3_cmp27_i_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_382to384_bb3_cmp27_i_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_382to384_bb3_cmp27_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb3_cmp27_i),
	.data_out(rnode_382to384_bb3_cmp27_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_382to384_bb3_cmp27_i_0_reg_384_fifo.DEPTH = 2;
defparam rnode_382to384_bb3_cmp27_i_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_382to384_bb3_cmp27_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to384_bb3_cmp27_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_382to384_bb3_cmp27_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp27_i_stall_in = 1'b0;
assign rnode_382to384_bb3_cmp27_i_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3_cmp27_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3_cmp27_i_0_NO_SHIFT_REG = rnode_382to384_bb3_cmp27_i_0_reg_384_NO_SHIFT_REG;
assign rnode_382to384_bb3_cmp27_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3_cmp27_i_1_NO_SHIFT_REG = rnode_382to384_bb3_cmp27_i_0_reg_384_NO_SHIFT_REG;
assign rnode_382to384_bb3_cmp27_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3_cmp27_i_2_NO_SHIFT_REG = rnode_382to384_bb3_cmp27_i_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_382to383_bb3_align_0_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3_align_0_i_0_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3_align_0_i_1_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3_align_0_i_2_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3_align_0_i_3_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3_align_0_i_4_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_reg_383_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb3_align_0_i_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_valid_out_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_stall_in_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb3_align_0_i_0_stall_out_reg_383_NO_SHIFT_REG;

acl_data_fifo rnode_382to383_bb3_align_0_i_0_reg_383_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to383_bb3_align_0_i_0_reg_383_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to383_bb3_align_0_i_0_stall_in_0_reg_383_NO_SHIFT_REG),
	.valid_out(rnode_382to383_bb3_align_0_i_0_valid_out_0_reg_383_NO_SHIFT_REG),
	.stall_out(rnode_382to383_bb3_align_0_i_0_stall_out_reg_383_NO_SHIFT_REG),
	.data_in((local_bb3_align_0_i & 32'hFF)),
	.data_out(rnode_382to383_bb3_align_0_i_0_reg_383_NO_SHIFT_REG)
);

defparam rnode_382to383_bb3_align_0_i_0_reg_383_fifo.DEPTH = 1;
defparam rnode_382to383_bb3_align_0_i_0_reg_383_fifo.DATA_WIDTH = 32;
defparam rnode_382to383_bb3_align_0_i_0_reg_383_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to383_bb3_align_0_i_0_reg_383_fifo.IMPL = "shift_reg";

assign rnode_382to383_bb3_align_0_i_0_reg_383_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_align_0_i_stall_in = 1'b0;
assign rnode_382to383_bb3_align_0_i_0_stall_in_0_reg_383_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_align_0_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3_align_0_i_0_NO_SHIFT_REG = rnode_382to383_bb3_align_0_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3_align_0_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3_align_0_i_1_NO_SHIFT_REG = rnode_382to383_bb3_align_0_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3_align_0_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3_align_0_i_2_NO_SHIFT_REG = rnode_382to383_bb3_align_0_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3_align_0_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3_align_0_i_3_NO_SHIFT_REG = rnode_382to383_bb3_align_0_i_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb3_align_0_i_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb3_align_0_i_4_NO_SHIFT_REG = rnode_382to383_bb3_align_0_i_0_reg_383_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__32_i210_stall_local;
wire [31:0] local_bb3__32_i210;

assign local_bb3__32_i210 = (local_bb3__31_i209 ? (local_bb3_shl1_i_i & 32'hFFFFFE00) : (local_bb3_shl1_i18_i & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__34_i_stall_local;
wire [31:0] local_bb3__34_i;

assign local_bb3__34_i = (local_bb3__31_i209 ? (local_bb3_or_i_i208 & 32'h1FFFFFF) : (local_bb3_or_i17_i & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__36_i_stall_local;
wire [31:0] local_bb3__36_i;

assign local_bb3__36_i = (local_bb3__31_i209 ? (rnode_381to383_bb3_add_i206_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb3_and21_i_stall_local;
wire [31:0] local_bb3_and21_i;

assign local_bb3_and21_i = (rnode_382to383_bb3__22_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and20_i_valid_out;
wire local_bb3_and20_i_stall_in;
wire local_bb3_and20_i_inputs_ready;
wire local_bb3_and20_i_stall_local;
wire [31:0] local_bb3_and20_i;

assign local_bb3_and20_i_inputs_ready = rnode_382to383_bb3__23_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_and20_i = (rnode_382to383_bb3__23_i_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb3_and20_i_valid_out = 1'b1;
assign rnode_382to383_bb3__23_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and35_i_valid_out;
wire local_bb3_and35_i_stall_in;
wire local_bb3_and35_i_inputs_ready;
wire local_bb3_and35_i_stall_local;
wire [31:0] local_bb3_and35_i;

assign local_bb3_and35_i_inputs_ready = rnode_382to383_bb3__23_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_and35_i = (rnode_382to383_bb3__23_i_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb3_and35_i_valid_out = 1'b1;
assign rnode_382to383_bb3__23_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_xor_i_stall_local;
wire [31:0] local_bb3_xor_i;

assign local_bb3_xor_i = (rnode_382to383_bb3__23_i_2_NO_SHIFT_REG ^ rnode_382to383_bb3__22_i_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_and17_i_stall_local;
wire [31:0] local_bb3_and17_i;

assign local_bb3_and17_i = ((rnode_382to384_bb3_shr16_i_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_384to386_bb3_shr16_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to386_bb3_shr16_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_384to386_bb3_shr16_i_0_NO_SHIFT_REG;
 logic rnode_384to386_bb3_shr16_i_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to386_bb3_shr16_i_0_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_shr16_i_0_valid_out_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_shr16_i_0_stall_in_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_shr16_i_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_384to386_bb3_shr16_i_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to386_bb3_shr16_i_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to386_bb3_shr16_i_0_stall_in_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_384to386_bb3_shr16_i_0_valid_out_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_384to386_bb3_shr16_i_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((rnode_382to384_bb3_shr16_i_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_384to386_bb3_shr16_i_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_384to386_bb3_shr16_i_0_reg_386_fifo.DEPTH = 2;
defparam rnode_384to386_bb3_shr16_i_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_384to386_bb3_shr16_i_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to386_bb3_shr16_i_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_384to386_bb3_shr16_i_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_382to384_bb3_shr16_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_shr16_i_0_NO_SHIFT_REG = rnode_384to386_bb3_shr16_i_0_reg_386_NO_SHIFT_REG;
assign rnode_384to386_bb3_shr16_i_0_stall_in_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_shr16_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and93_i_stall_local;
wire [31:0] local_bb3_and93_i;

assign local_bb3_and93_i = ((rnode_382to383_bb3_align_0_i_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb3_and95_i_stall_local;
wire [31:0] local_bb3_and95_i;

assign local_bb3_and95_i = ((rnode_382to383_bb3_align_0_i_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and115_i_stall_local;
wire [31:0] local_bb3_and115_i;

assign local_bb3_and115_i = ((rnode_382to383_bb3_align_0_i_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_and130_i_stall_local;
wire [31:0] local_bb3_and130_i;

assign local_bb3_and130_i = ((rnode_382to383_bb3_align_0_i_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb3_and149_i_stall_local;
wire [31:0] local_bb3_and149_i;

assign local_bb3_and149_i = ((rnode_382to383_bb3_align_0_i_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb3__33_i211_stall_local;
wire [31:0] local_bb3__33_i211;

assign local_bb3__33_i211 = (local_bb3_tobool49_i ? (local_bb3__32_i210 & 32'hFFFFFF00) : (local_bb3_shl1_i18_i & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb3__35_i_stall_local;
wire [31:0] local_bb3__35_i;

assign local_bb3__35_i = (local_bb3_tobool49_i ? (local_bb3__34_i & 32'h1FFFFFF) : (local_bb3_or_i17_i & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__37_i_stall_local;
wire [31:0] local_bb3__37_i;

assign local_bb3__37_i = (local_bb3_tobool49_i ? (local_bb3__36_i & 32'h1FF) : (local_bb3_inc_i & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot33_not_i_stall_local;
wire local_bb3_lnot33_not_i;

assign local_bb3_lnot33_not_i = ((local_bb3_and21_i & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or64_i_stall_local;
wire [31:0] local_bb3_or64_i;

assign local_bb3_or64_i = ((local_bb3_and21_i & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_and20_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and20_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and20_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and20_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and20_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and20_i_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and20_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and20_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and20_i_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and20_i_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and20_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_and20_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_and20_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_and20_i_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_and20_i_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_and20_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb3_and20_i & 32'h7FFFFF)),
	.data_out(rnode_383to384_bb3_and20_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_and20_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_and20_i_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb3_and20_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_and20_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_and20_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and20_i_stall_in = 1'b0;
assign rnode_383to384_bb3_and20_i_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and20_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3_and20_i_0_NO_SHIFT_REG = rnode_383to384_bb3_and20_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_and20_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3_and20_i_1_NO_SHIFT_REG = rnode_383to384_bb3_and20_i_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and35_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and35_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and35_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and35_i_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and35_i_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and35_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_and35_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_and35_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_and35_i_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_and35_i_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_and35_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb3_and35_i & 32'h80000000)),
	.data_out(rnode_383to384_bb3_and35_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_and35_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_and35_i_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb3_and35_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_and35_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_and35_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and35_i_stall_in = 1'b0;
assign rnode_383to384_bb3_and35_i_0_NO_SHIFT_REG = rnode_383to384_bb3_and35_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_and35_i_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp37_i_stall_local;
wire local_bb3_cmp37_i;

assign local_bb3_cmp37_i = ($signed(local_bb3_xor_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb3_xor_lobit_i_stall_local;
wire [31:0] local_bb3_xor_lobit_i;

assign local_bb3_xor_lobit_i = ($signed(local_bb3_xor_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_and36_lobit_i_stall_local;
wire [31:0] local_bb3_and36_lobit_i;

assign local_bb3_and36_lobit_i = (local_bb3_xor_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_i_stall_local;
wire local_bb3_lnot_i;

assign local_bb3_lnot_i = ((local_bb3_and17_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_i5_stall_local;
wire local_bb3_cmp25_i5;

assign local_bb3_cmp25_i5 = ((local_bb3_and17_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp96_i_stall_local;
wire local_bb3_cmp96_i;

assign local_bb3_cmp96_i = ((local_bb3_and95_i & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp116_i_stall_local;
wire local_bb3_cmp116_i;

assign local_bb3_cmp116_i = ((local_bb3_and115_i & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp131_not_i_stall_local;
wire local_bb3_cmp131_not_i;

assign local_bb3_cmp131_not_i = ((local_bb3_and130_i & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_Pivot20_i_stall_local;
wire local_bb3_Pivot20_i;

assign local_bb3_Pivot20_i = ((local_bb3_and149_i & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_SwitchLeaf_i_stall_local;
wire local_bb3_SwitchLeaf_i;

assign local_bb3_SwitchLeaf_i = ((local_bb3_and149_i & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and75_i214_stall_local;
wire [31:0] local_bb3_and75_i214;

assign local_bb3_and75_i214 = ((local_bb3__35_i & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3__33_i211_valid_out;
wire local_bb3__33_i211_stall_in;
wire local_bb3__37_i_valid_out;
wire local_bb3__37_i_stall_in;
wire local_bb3_and75_i214_valid_out;
wire local_bb3_and75_i214_stall_in;
wire local_bb3_and83_i_valid_out;
wire local_bb3_and83_i_stall_in;
wire local_bb3_and83_i_inputs_ready;
wire local_bb3_and83_i_stall_local;
wire [31:0] local_bb3_and83_i;

assign local_bb3_and83_i_inputs_ready = (local_bb3_mul_i_i_valid_out_0_NO_SHIFT_REG & rnode_381to383_bb3_add_i206_0_valid_out_1_NO_SHIFT_REG & rnode_381to383_bb3_add_i206_0_valid_out_0_NO_SHIFT_REG & rnode_381to383_bb3_add_i206_0_valid_out_2_NO_SHIFT_REG & local_bb3_mul_i_i_valid_out_1_NO_SHIFT_REG);
assign local_bb3_and83_i = ((local_bb3__35_i & 32'h1FFFFFF) & 32'h1);
assign local_bb3__33_i211_valid_out = 1'b1;
assign local_bb3__37_i_valid_out = 1'b1;
assign local_bb3_and75_i214_valid_out = 1'b1;
assign local_bb3_and83_i_valid_out = 1'b1;
assign local_bb3_mul_i_i_stall_in_0 = 1'b0;
assign rnode_381to383_bb3_add_i206_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_381to383_bb3_add_i206_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_381to383_bb3_add_i206_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign local_bb3_mul_i_i_stall_in_1 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_shl65_i_stall_local;
wire [31:0] local_bb3_shl65_i;

assign local_bb3_shl65_i = ((local_bb3_or64_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot30_i_stall_local;
wire local_bb3_lnot30_i;

assign local_bb3_lnot30_i = ((rnode_383to384_bb3_and20_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i6_stall_local;
wire [31:0] local_bb3_or_i6;

assign local_bb3_or_i6 = ((rnode_383to384_bb3_and20_i_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_384to386_bb3_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_384to386_bb3_and35_i_0_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and35_i_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to386_bb3_and35_i_0_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and35_i_0_valid_out_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and35_i_0_stall_in_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and35_i_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_384to386_bb3_and35_i_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to386_bb3_and35_i_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to386_bb3_and35_i_0_stall_in_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_384to386_bb3_and35_i_0_valid_out_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_384to386_bb3_and35_i_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((rnode_383to384_bb3_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_384to386_bb3_and35_i_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_384to386_bb3_and35_i_0_reg_386_fifo.DEPTH = 2;
defparam rnode_384to386_bb3_and35_i_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_384to386_bb3_and35_i_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to386_bb3_and35_i_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_384to386_bb3_and35_i_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_and35_i_0_NO_SHIFT_REG = rnode_384to386_bb3_and35_i_0_reg_386_NO_SHIFT_REG;
assign rnode_384to386_bb3_and35_i_0_stall_in_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_not_i_stall_local;
wire local_bb3_cmp25_not_i;

assign local_bb3_cmp25_not_i = (local_bb3_cmp25_i5 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u72_stall_local;
wire local_bb3_var__u72;

assign local_bb3_var__u72 = (local_bb3_cmp25_i5 | rnode_382to384_bb3_cmp27_i_2_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3__33_i211_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3__33_i211_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__33_i211_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3__33_i211_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3__33_i211_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__33_i211_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3__33_i211_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__33_i211_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3__33_i211_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3__33_i211_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3__33_i211_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3__33_i211_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3__33_i211_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3__33_i211_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3__33_i211_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3__33_i211_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb3__33_i211 & 32'hFFFFFF00)),
	.data_out(rnode_383to384_bb3__33_i211_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3__33_i211_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3__33_i211_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb3__33_i211_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3__33_i211_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3__33_i211_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__33_i211_stall_in = 1'b0;
assign rnode_383to384_bb3__33_i211_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3__33_i211_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3__33_i211_0_NO_SHIFT_REG = rnode_383to384_bb3__33_i211_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3__33_i211_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3__33_i211_1_NO_SHIFT_REG = rnode_383to384_bb3__33_i211_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3__37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__37_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__37_i_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__37_i_2_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__37_i_3_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3__37_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3__37_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3__37_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3__37_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3__37_i_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3__37_i_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3__37_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb3__37_i & 32'h3FF)),
	.data_out(rnode_383to384_bb3__37_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3__37_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3__37_i_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb3__37_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3__37_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3__37_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__37_i_stall_in = 1'b0;
assign rnode_383to384_bb3__37_i_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3__37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3__37_i_0_NO_SHIFT_REG = rnode_383to384_bb3__37_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3__37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3__37_i_1_NO_SHIFT_REG = rnode_383to384_bb3__37_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3__37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3__37_i_2_NO_SHIFT_REG = rnode_383to384_bb3__37_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3__37_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3__37_i_3_NO_SHIFT_REG = rnode_383to384_bb3__37_i_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_383to385_bb3_and75_i214_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to385_bb3_and75_i214_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_383to385_bb3_and75_i214_0_NO_SHIFT_REG;
 logic rnode_383to385_bb3_and75_i214_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to385_bb3_and75_i214_0_reg_385_NO_SHIFT_REG;
 logic rnode_383to385_bb3_and75_i214_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_383to385_bb3_and75_i214_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_383to385_bb3_and75_i214_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_383to385_bb3_and75_i214_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to385_bb3_and75_i214_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to385_bb3_and75_i214_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_383to385_bb3_and75_i214_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_383to385_bb3_and75_i214_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in((local_bb3_and75_i214 & 32'h7FFFFF)),
	.data_out(rnode_383to385_bb3_and75_i214_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_383to385_bb3_and75_i214_0_reg_385_fifo.DEPTH = 2;
defparam rnode_383to385_bb3_and75_i214_0_reg_385_fifo.DATA_WIDTH = 32;
defparam rnode_383to385_bb3_and75_i214_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to385_bb3_and75_i214_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_383to385_bb3_and75_i214_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and75_i214_stall_in = 1'b0;
assign rnode_383to385_bb3_and75_i214_0_NO_SHIFT_REG = rnode_383to385_bb3_and75_i214_0_reg_385_NO_SHIFT_REG;
assign rnode_383to385_bb3_and75_i214_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_383to385_bb3_and75_i214_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_and83_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and83_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and83_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and83_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and83_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and83_i_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and83_i_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and83_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_and83_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_and83_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_and83_i_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_and83_i_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_and83_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb3_and83_i & 32'h1)),
	.data_out(rnode_383to384_bb3_and83_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_and83_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_and83_i_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb3_and83_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_and83_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_and83_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and83_i_stall_in = 1'b0;
assign rnode_383to384_bb3_and83_i_0_NO_SHIFT_REG = rnode_383to384_bb3_and83_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_and83_i_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and83_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__28_i_stall_local;
wire [31:0] local_bb3__28_i;

assign local_bb3__28_i = (rnode_382to383_bb3_lnot23_i_0_NO_SHIFT_REG ? 32'h0 : ((local_bb3_shl65_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot30_not_i_stall_local;
wire local_bb3_lnot30_not_i;

assign local_bb3_lnot30_not_i = (local_bb3_lnot30_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i7_stall_local;
wire [31:0] local_bb3_shl_i7;

assign local_bb3_shl_i7 = ((local_bb3_or_i6 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_and35_i_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and35_i_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_and35_i_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and35_i_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and35_i_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and35_i_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_and35_i_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_and35_i_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_and35_i_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_and35_i_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_and35_i_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in((rnode_384to386_bb3_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_386to387_bb3_and35_i_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_and35_i_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_and35_i_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb3_and35_i_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_and35_i_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_and35_i_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_384to386_bb3_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_and35_i_0_NO_SHIFT_REG = rnode_386to387_bb3_and35_i_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_and35_i_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_or_cond_i_stall_local;
wire local_bb3_or_cond_i;

assign local_bb3_or_cond_i = (local_bb3_lnot30_i | local_bb3_cmp25_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp77_i_stall_local;
wire local_bb3_cmp77_i;

assign local_bb3_cmp77_i = ((rnode_383to384_bb3__33_i211_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u73_stall_local;
wire local_bb3_var__u73;

assign local_bb3_var__u73 = ($signed((rnode_383to384_bb3__33_i211_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp53_i_stall_local;
wire local_bb3_cmp53_i;

assign local_bb3_cmp53_i = ((rnode_383to384_bb3__37_i_0_NO_SHIFT_REG & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp68_i_valid_out;
wire local_bb3_cmp68_i_stall_in;
wire local_bb3_cmp68_i_inputs_ready;
wire local_bb3_cmp68_i_stall_local;
wire local_bb3_cmp68_i;

assign local_bb3_cmp68_i_inputs_ready = rnode_383to384_bb3__37_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_cmp68_i = ((rnode_383to384_bb3__37_i_1_NO_SHIFT_REG & 32'h3FF) < 32'h80);
assign local_bb3_cmp68_i_valid_out = 1'b1;
assign rnode_383to384_bb3__37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_sub_i215_stall_local;
wire [31:0] local_bb3_sub_i215;

assign local_bb3_sub_i215 = ((rnode_383to384_bb3__37_i_2_NO_SHIFT_REG & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp71_not_i_valid_out;
wire local_bb3_cmp71_not_i_stall_in;
wire local_bb3_cmp71_not_i_inputs_ready;
wire local_bb3_cmp71_not_i_stall_local;
wire local_bb3_cmp71_not_i;

assign local_bb3_cmp71_not_i_inputs_ready = rnode_383to384_bb3__37_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb3_cmp71_not_i = ((rnode_383to384_bb3__37_i_3_NO_SHIFT_REG & 32'h3FF) != 32'h7F);
assign local_bb3_cmp71_not_i_valid_out = 1'b1;
assign rnode_383to384_bb3__37_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_tobool84_i_stall_local;
wire local_bb3_tobool84_i;

assign local_bb3_tobool84_i = ((rnode_383to384_bb3_and83_i_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and72_i_stall_local;
wire [31:0] local_bb3_and72_i;

assign local_bb3_and72_i = ((local_bb3__28_i & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb3_and75_i_stall_local;
wire [31:0] local_bb3_and75_i;

assign local_bb3_and75_i = ((local_bb3__28_i & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb3_and78_i_stall_local;
wire [31:0] local_bb3_and78_i;

assign local_bb3_and78_i = ((local_bb3__28_i & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb3_shr94_i_stall_local;
wire [31:0] local_bb3_shr94_i;

assign local_bb3_shr94_i = ((local_bb3__28_i & 32'h7FFFFF8) >> (local_bb3_and93_i & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb3_and90_i_stall_local;
wire [31:0] local_bb3_and90_i;

assign local_bb3_and90_i = ((local_bb3__28_i & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb3_and87_i_stall_local;
wire [31:0] local_bb3_and87_i;

assign local_bb3_and87_i = ((local_bb3__28_i & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb3_and84_i_stall_local;
wire [31:0] local_bb3_and84_i;

assign local_bb3_and84_i = ((local_bb3__28_i & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u74_stall_local;
wire [31:0] local_bb3_var__u74;

assign local_bb3_var__u74 = ((local_bb3__28_i & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb3_or_cond_not_i_stall_local;
wire local_bb3_or_cond_not_i;

assign local_bb3_or_cond_not_i = (local_bb3_cmp25_i5 & local_bb3_lnot30_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3__27_i_stall_local;
wire [31:0] local_bb3__27_i;

assign local_bb3__27_i = (local_bb3_lnot_i ? 32'h0 : ((local_bb3_shl_i7 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_8_i_stall_local;
wire local_bb3_reduction_8_i;

assign local_bb3_reduction_8_i = (rnode_382to384_bb3_cmp27_i_1_NO_SHIFT_REG & local_bb3_or_cond_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or581_i_valid_out;
wire local_bb3_or581_i_stall_in;
wire local_bb3_or581_i_inputs_ready;
wire local_bb3_or581_i_stall_local;
wire local_bb3_or581_i;

assign local_bb3_or581_i_inputs_ready = (rnode_383to384_bb3_var__u70_0_valid_out_NO_SHIFT_REG & rnode_383to384_bb3__37_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3_or581_i = (rnode_383to384_bb3_var__u70_0_NO_SHIFT_REG | local_bb3_cmp53_i);
assign local_bb3_or581_i_valid_out = 1'b1;
assign rnode_383to384_bb3_var__u70_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3__37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_cmp68_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp68_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp68_i_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp68_i_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp68_i_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp68_i_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp68_i_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp68_i_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_cmp68_i_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_cmp68_i_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_cmp68_i_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_cmp68_i_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_cmp68_i_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb3_cmp68_i),
	.data_out(rnode_384to385_bb3_cmp68_i_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_cmp68_i_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_cmp68_i_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3_cmp68_i_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_cmp68_i_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_cmp68_i_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp68_i_stall_in = 1'b0;
assign rnode_384to385_bb3_cmp68_i_0_NO_SHIFT_REG = rnode_384to385_bb3_cmp68_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_cmp68_i_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_cmp68_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and74_i_stall_local;
wire [31:0] local_bb3_and74_i;

assign local_bb3_and74_i = ((local_bb3_sub_i215 & 32'hFF800000) + 32'h40800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_cmp71_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp71_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp71_not_i_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp71_not_i_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp71_not_i_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp71_not_i_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp71_not_i_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_cmp71_not_i_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_cmp71_not_i_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_cmp71_not_i_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_cmp71_not_i_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_cmp71_not_i_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_cmp71_not_i_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb3_cmp71_not_i),
	.data_out(rnode_384to385_bb3_cmp71_not_i_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_cmp71_not_i_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_cmp71_not_i_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3_cmp71_not_i_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_cmp71_not_i_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_cmp71_not_i_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp71_not_i_stall_in = 1'b0;
assign rnode_384to385_bb3_cmp71_not_i_0_NO_SHIFT_REG = rnode_384to385_bb3_cmp71_not_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_cmp71_not_i_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_cmp71_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__39_i_stall_local;
wire local_bb3__39_i;

assign local_bb3__39_i = (local_bb3_tobool84_i & local_bb3_var__u73);

// This section implements an unregistered operation.
// 
wire local_bb3_and72_tr_i_stall_local;
wire [7:0] local_bb3_and72_tr_i;
wire [31:0] local_bb3_and72_tr_i$ps;

assign local_bb3_and72_tr_i$ps = (local_bb3_and72_i & 32'hFFFFFF);
assign local_bb3_and72_tr_i = local_bb3_and72_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb3_cmp76_i_stall_local;
wire local_bb3_cmp76_i;

assign local_bb3_cmp76_i = ((local_bb3_and75_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp79_i_stall_local;
wire local_bb3_cmp79_i;

assign local_bb3_cmp79_i = ((local_bb3_and78_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and142_i_stall_local;
wire [31:0] local_bb3_and142_i;

assign local_bb3_and142_i = (local_bb3_shr94_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_shr150_i_stall_local;
wire [31:0] local_bb3_shr150_i;

assign local_bb3_shr150_i = (local_bb3_shr94_i >> (local_bb3_and149_i & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u75_stall_local;
wire [31:0] local_bb3_var__u75;

assign local_bb3_var__u75 = (local_bb3_shr94_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and146_i_stall_local;
wire [31:0] local_bb3_and146_i;

assign local_bb3_and146_i = (local_bb3_shr94_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp91_i_stall_local;
wire local_bb3_cmp91_i;

assign local_bb3_cmp91_i = ((local_bb3_and90_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp88_i_stall_local;
wire local_bb3_cmp88_i;

assign local_bb3_cmp88_i = ((local_bb3_and87_i & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp85_i_stall_local;
wire local_bb3_cmp85_i;

assign local_bb3_cmp85_i = ((local_bb3_and84_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u76_stall_local;
wire local_bb3_var__u76;

assign local_bb3_var__u76 = ((local_bb3_var__u74 & 32'hFFF8) != 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_or581_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_1_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_valid_out_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_stall_in_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_or581_i_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_or581_i_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_or581_i_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_or581_i_0_stall_in_0_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_or581_i_0_valid_out_0_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_or581_i_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb3_or581_i),
	.data_out(rnode_384to385_bb3_or581_i_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_or581_i_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_or581_i_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3_or581_i_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_or581_i_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_or581_i_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or581_i_stall_in = 1'b0;
assign rnode_384to385_bb3_or581_i_0_stall_in_0_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_or581_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3_or581_i_0_NO_SHIFT_REG = rnode_384to385_bb3_or581_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_or581_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3_or581_i_1_NO_SHIFT_REG = rnode_384to385_bb3_or581_i_0_reg_385_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u77_stall_local;
wire [31:0] local_bb3_var__u77;

assign local_bb3_var__u77[31:1] = 31'h0;
assign local_bb3_var__u77[0] = rnode_384to385_bb3_cmp68_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i216_valid_out;
wire local_bb3_shl_i216_stall_in;
wire local_bb3_shl_i216_inputs_ready;
wire local_bb3_shl_i216_stall_local;
wire [31:0] local_bb3_shl_i216;

assign local_bb3_shl_i216_inputs_ready = rnode_383to384_bb3__37_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_shl_i216 = ((local_bb3_and74_i & 32'hFF800000) & 32'h7F800000);
assign local_bb3_shl_i216_valid_out = 1'b1;
assign rnode_383to384_bb3__37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__40_i_valid_out;
wire local_bb3__40_i_stall_in;
wire local_bb3__40_i_inputs_ready;
wire local_bb3__40_i_stall_local;
wire local_bb3__40_i;

assign local_bb3__40_i_inputs_ready = (rnode_383to384_bb3__33_i211_0_valid_out_0_NO_SHIFT_REG & rnode_383to384_bb3__33_i211_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb3_and83_i_0_valid_out_NO_SHIFT_REG);
assign local_bb3__40_i = (local_bb3_cmp77_i | local_bb3__39_i);
assign local_bb3__40_i_valid_out = 1'b1;
assign rnode_383to384_bb3__33_i211_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3__33_i211_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and83_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_frombool74_i_stall_local;
wire [7:0] local_bb3_frombool74_i;

assign local_bb3_frombool74_i = (local_bb3_and72_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u78_stall_local;
wire [31:0] local_bb3_var__u78;

assign local_bb3_var__u78 = ((local_bb3_and146_i & 32'h3FFFFFFF) | local_bb3_shr94_i);

// This section implements an unregistered operation.
// 
wire local_bb3__31_v_i_stall_local;
wire local_bb3__31_v_i;

assign local_bb3__31_v_i = (local_bb3_cmp96_i ? local_bb3_cmp79_i : local_bb3_cmp91_i);

// This section implements an unregistered operation.
// 
wire local_bb3__30_v_i_stall_local;
wire local_bb3__30_v_i;

assign local_bb3__30_v_i = (local_bb3_cmp96_i ? local_bb3_cmp76_i : local_bb3_cmp88_i);

// This section implements an unregistered operation.
// 
wire local_bb3_frombool109_i_stall_local;
wire [7:0] local_bb3_frombool109_i;

assign local_bb3_frombool109_i[7:1] = 7'h0;
assign local_bb3_frombool109_i[0] = local_bb3_cmp85_i;

// This section implements an unregistered operation.
// 
wire local_bb3_or107_i_stall_local;
wire [31:0] local_bb3_or107_i;

assign local_bb3_or107_i[31:1] = 31'h0;
assign local_bb3_or107_i[0] = local_bb3_var__u76;

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_2_i213_stall_local;
wire local_bb3_reduction_2_i213;

assign local_bb3_reduction_2_i213 = (rnode_384to385_bb3_reduction_0_i212_0_NO_SHIFT_REG | rnode_384to385_bb3_or581_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_cond111_i_stall_local;
wire [31:0] local_bb3_cond111_i;

assign local_bb3_cond111_i = (rnode_384to385_bb3_or581_i_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_shl_i216_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3_shl_i216_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_shl_i216_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_shl_i216_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_shl_i216_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_shl_i216_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_shl_i216_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_shl_i216_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_shl_i216_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_shl_i216_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_shl_i216_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_shl_i216_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_shl_i216_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in((local_bb3_shl_i216 & 32'h7F800000)),
	.data_out(rnode_384to385_bb3_shl_i216_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_shl_i216_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_shl_i216_0_reg_385_fifo.DATA_WIDTH = 32;
defparam rnode_384to385_bb3_shl_i216_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_shl_i216_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_shl_i216_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shl_i216_stall_in = 1'b0;
assign rnode_384to385_bb3_shl_i216_0_NO_SHIFT_REG = rnode_384to385_bb3_shl_i216_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_shl_i216_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_shl_i216_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3__40_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3__40_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb3__40_i_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3__40_i_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3__40_i_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__40_i_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__40_i_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__40_i_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3__40_i_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3__40_i_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3__40_i_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3__40_i_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3__40_i_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb3__40_i),
	.data_out(rnode_384to385_bb3__40_i_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3__40_i_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3__40_i_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3__40_i_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3__40_i_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3__40_i_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__40_i_stall_in = 1'b0;
assign rnode_384to385_bb3__40_i_0_NO_SHIFT_REG = rnode_384to385_bb3__40_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3__40_i_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3__40_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_or1596_i_stall_local;
wire [31:0] local_bb3_or1596_i;

assign local_bb3_or1596_i = (local_bb3_var__u78 | (local_bb3_and142_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__31_i_stall_local;
wire [7:0] local_bb3__31_i;

assign local_bb3__31_i[7:1] = 7'h0;
assign local_bb3__31_i[0] = local_bb3__31_v_i;

// This section implements an unregistered operation.
// 
wire local_bb3__30_i_stall_local;
wire [7:0] local_bb3__30_i;

assign local_bb3__30_i[7:1] = 7'h0;
assign local_bb3__30_i[0] = local_bb3__30_v_i;

// This section implements an unregistered operation.
// 
wire local_bb3__29_i_stall_local;
wire [7:0] local_bb3__29_i;

assign local_bb3__29_i = (local_bb3_cmp96_i ? (local_bb3_frombool74_i & 8'h1) : (local_bb3_frombool109_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__32_i_stall_local;
wire [31:0] local_bb3__32_i;

assign local_bb3__32_i = (local_bb3_cmp96_i ? 32'h0 : (local_bb3_or107_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_conv101_i_stall_local;
wire [31:0] local_bb3_conv101_i;

assign local_bb3_conv101_i[31:1] = 31'h0;
assign local_bb3_conv101_i[0] = local_bb3_reduction_2_i213;

// This section implements an unregistered operation.
// 
wire local_bb3_or76_i_stall_local;
wire [31:0] local_bb3_or76_i;

assign local_bb3_or76_i = ((rnode_384to385_bb3_shl_i216_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_383to385_bb3_and75_i214_0_NO_SHIFT_REG & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cond_i217_stall_local;
wire [31:0] local_bb3_cond_i217;

assign local_bb3_cond_i217[31:1] = 31'h0;
assign local_bb3_cond_i217[0] = rnode_384to385_bb3__40_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or162_i_stall_local;
wire [31:0] local_bb3_or162_i;

assign local_bb3_or162_i = (local_bb3_or1596_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or1237_i_stall_local;
wire [7:0] local_bb3_or1237_i;

assign local_bb3_or1237_i = ((local_bb3__30_i & 8'h1) | (local_bb3__29_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__33_i_stall_local;
wire [7:0] local_bb3__33_i;

assign local_bb3__33_i = (local_bb3_cmp116_i ? (local_bb3__29_i & 8'h1) : (local_bb3__31_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_add87_i_stall_local;
wire [31:0] local_bb3_add87_i;

assign local_bb3_add87_i = ((local_bb3_cond_i217 & 32'h1) + (local_bb3_or76_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__37_v_i_stall_local;
wire [31:0] local_bb3__37_v_i;

assign local_bb3__37_v_i = (local_bb3_Pivot20_i ? 32'h0 : (local_bb3_or162_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or123_i_stall_local;
wire [31:0] local_bb3_or123_i;

assign local_bb3_or123_i[31:8] = 24'h0;
assign local_bb3_or123_i[7:0] = (local_bb3_or1237_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u79_stall_local;
wire [7:0] local_bb3_var__u79;

assign local_bb3_var__u79 = ((local_bb3__33_i & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and88_i_stall_local;
wire [31:0] local_bb3_and88_i;

assign local_bb3_and88_i = (local_bb3_add87_i & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and90_i218_stall_local;
wire [31:0] local_bb3_and90_i218;

assign local_bb3_and90_i218 = (local_bb3_add87_i & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb3__39_v_i_stall_local;
wire [31:0] local_bb3__39_v_i;

assign local_bb3__39_v_i = (local_bb3_SwitchLeaf_i ? (local_bb3_var__u75 & 32'h1) : (local_bb3__37_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or124_i_stall_local;
wire [31:0] local_bb3_or124_i;

assign local_bb3_or124_i = (local_bb3_cmp116_i ? 32'h0 : (local_bb3_or123_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_conv135_i_stall_local;
wire [31:0] local_bb3_conv135_i;

assign local_bb3_conv135_i[31:8] = 24'h0;
assign local_bb3_conv135_i[7:0] = (local_bb3_var__u79 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or89_i_stall_local;
wire [31:0] local_bb3_or89_i;

assign local_bb3_or89_i = ((local_bb3_and88_i & 32'h7FFFFFFF) | (local_bb3_and4_i & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp91_i219_stall_local;
wire local_bb3_cmp91_i219;

assign local_bb3_cmp91_i219 = ((local_bb3_and90_i218 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_3_i_stall_local;
wire [31:0] local_bb3_reduction_3_i;

assign local_bb3_reduction_3_i = ((local_bb3__32_i & 32'h1) | (local_bb3_or124_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or136_i_stall_local;
wire [31:0] local_bb3_or136_i;

assign local_bb3_or136_i = (local_bb3_cmp131_not_i ? (local_bb3_conv135_i & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge14_i_stall_local;
wire local_bb3_brmerge14_i;

assign local_bb3_brmerge14_i = (local_bb3_cmp91_i219 | rnode_384to385_bb3_cmp71_not_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_5_i_stall_local;
wire [31:0] local_bb3_reduction_5_i;

assign local_bb3_reduction_5_i = (local_bb3_shr150_i | (local_bb3_reduction_3_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_4_i_stall_local;
wire [31:0] local_bb3_reduction_4_i;

assign local_bb3_reduction_4_i = ((local_bb3_or136_i & 32'h1) | (local_bb3__39_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_conv99_i_stall_local;
wire [31:0] local_bb3_conv99_i;

assign local_bb3_conv99_i = (local_bb3_brmerge14_i ? (local_bb3_var__u77 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_6_i_stall_local;
wire [31:0] local_bb3_reduction_6_i;

assign local_bb3_reduction_6_i = ((local_bb3_reduction_4_i & 32'h1) | local_bb3_reduction_5_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or102_i_stall_local;
wire [31:0] local_bb3_or102_i;

assign local_bb3_or102_i = ((local_bb3_conv99_i & 32'h1) | (local_bb3_conv101_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot33_not_i_valid_out;
wire local_bb3_lnot33_not_i_stall_in;
wire local_bb3_cmp37_i_valid_out;
wire local_bb3_cmp37_i_stall_in;
wire local_bb3_and36_lobit_i_valid_out;
wire local_bb3_and36_lobit_i_stall_in;
wire local_bb3_xor188_i_valid_out;
wire local_bb3_xor188_i_stall_in;
wire local_bb3_xor188_i_inputs_ready;
wire local_bb3_xor188_i_stall_local;
wire [31:0] local_bb3_xor188_i;

assign local_bb3_xor188_i_inputs_ready = (rnode_382to383_bb3__22_i_0_valid_out_0_NO_SHIFT_REG & rnode_382to383_bb3_lnot23_i_0_valid_out_NO_SHIFT_REG & rnode_382to383_bb3_align_0_i_0_valid_out_0_NO_SHIFT_REG & rnode_382to383_bb3_align_0_i_0_valid_out_4_NO_SHIFT_REG & rnode_382to383_bb3_align_0_i_0_valid_out_1_NO_SHIFT_REG & rnode_382to383_bb3_align_0_i_0_valid_out_2_NO_SHIFT_REG & rnode_382to383_bb3_align_0_i_0_valid_out_3_NO_SHIFT_REG & rnode_382to383_bb3__23_i_0_valid_out_2_NO_SHIFT_REG & rnode_382to383_bb3__22_i_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_xor188_i = (local_bb3_reduction_6_i ^ local_bb3_xor_lobit_i);
assign local_bb3_lnot33_not_i_valid_out = 1'b1;
assign local_bb3_cmp37_i_valid_out = 1'b1;
assign local_bb3_and36_lobit_i_valid_out = 1'b1;
assign local_bb3_xor188_i_valid_out = 1'b1;
assign rnode_382to383_bb3__22_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_lnot23_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_align_0_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_align_0_i_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_align_0_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_align_0_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3_align_0_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3__23_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb3__22_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_tobool103_i_stall_local;
wire local_bb3_tobool103_i;

assign local_bb3_tobool103_i = ((local_bb3_or102_i & 32'h1) != 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_lnot33_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb3_lnot33_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_383to384_bb3_lnot33_not_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_lnot33_not_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb3_lnot33_not_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_lnot33_not_i_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_lnot33_not_i_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_lnot33_not_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_lnot33_not_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_lnot33_not_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_lnot33_not_i_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_lnot33_not_i_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_lnot33_not_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb3_lnot33_not_i),
	.data_out(rnode_383to384_bb3_lnot33_not_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_lnot33_not_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_lnot33_not_i_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb3_lnot33_not_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_lnot33_not_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_lnot33_not_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_lnot33_not_i_stall_in = 1'b0;
assign rnode_383to384_bb3_lnot33_not_i_0_NO_SHIFT_REG = rnode_383to384_bb3_lnot33_not_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_lnot33_not_i_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_lnot33_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_cmp37_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_cmp37_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_cmp37_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_cmp37_i_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_cmp37_i_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_cmp37_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb3_cmp37_i),
	.data_out(rnode_383to384_bb3_cmp37_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_cmp37_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_cmp37_i_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb3_cmp37_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_cmp37_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_cmp37_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp37_i_stall_in = 1'b0;
assign rnode_383to384_bb3_cmp37_i_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3_cmp37_i_0_NO_SHIFT_REG = rnode_383to384_bb3_cmp37_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3_cmp37_i_1_NO_SHIFT_REG = rnode_383to384_bb3_cmp37_i_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_and36_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and36_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and36_lobit_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and36_lobit_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_and36_lobit_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and36_lobit_i_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and36_lobit_i_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_and36_lobit_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_and36_lobit_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_and36_lobit_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_and36_lobit_i_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_and36_lobit_i_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_and36_lobit_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb3_and36_lobit_i & 32'h1)),
	.data_out(rnode_383to384_bb3_and36_lobit_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_and36_lobit_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_and36_lobit_i_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb3_and36_lobit_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_and36_lobit_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_and36_lobit_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and36_lobit_i_stall_in = 1'b0;
assign rnode_383to384_bb3_and36_lobit_i_0_NO_SHIFT_REG = rnode_383to384_bb3_and36_lobit_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_and36_lobit_i_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and36_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb3_xor188_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb3_xor188_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_xor188_i_0_NO_SHIFT_REG;
 logic rnode_383to384_bb3_xor188_i_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb3_xor188_i_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_xor188_i_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_xor188_i_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb3_xor188_i_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb3_xor188_i_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb3_xor188_i_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb3_xor188_i_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb3_xor188_i_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb3_xor188_i_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb3_xor188_i),
	.data_out(rnode_383to384_bb3_xor188_i_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb3_xor188_i_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb3_xor188_i_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb3_xor188_i_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb3_xor188_i_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb3_xor188_i_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_xor188_i_stall_in = 1'b0;
assign rnode_383to384_bb3_xor188_i_0_NO_SHIFT_REG = rnode_383to384_bb3_xor188_i_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb3_xor188_i_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_xor188_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cond107_i_stall_local;
wire [31:0] local_bb3_cond107_i;

assign local_bb3_cond107_i = (local_bb3_tobool103_i ? (local_bb3_and4_i & 32'h80000000) : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge_not_i_stall_local;
wire local_bb3_brmerge_not_i;

assign local_bb3_brmerge_not_i = (rnode_382to384_bb3_cmp27_i_0_NO_SHIFT_REG & rnode_383to384_bb3_lnot33_not_i_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_384to386_bb3_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_2_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_valid_out_0_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_stall_in_0_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_cmp37_i_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_384to386_bb3_cmp37_i_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to386_bb3_cmp37_i_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to386_bb3_cmp37_i_0_stall_in_0_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_384to386_bb3_cmp37_i_0_valid_out_0_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_384to386_bb3_cmp37_i_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in(rnode_383to384_bb3_cmp37_i_1_NO_SHIFT_REG),
	.data_out(rnode_384to386_bb3_cmp37_i_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_384to386_bb3_cmp37_i_0_reg_386_fifo.DEPTH = 2;
defparam rnode_384to386_bb3_cmp37_i_0_reg_386_fifo.DATA_WIDTH = 1;
defparam rnode_384to386_bb3_cmp37_i_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to386_bb3_cmp37_i_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_384to386_bb3_cmp37_i_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb3_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_cmp37_i_0_stall_in_0_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_384to386_bb3_cmp37_i_0_NO_SHIFT_REG = rnode_384to386_bb3_cmp37_i_0_reg_386_NO_SHIFT_REG;
assign rnode_384to386_bb3_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_384to386_bb3_cmp37_i_1_NO_SHIFT_REG = rnode_384to386_bb3_cmp37_i_0_reg_386_NO_SHIFT_REG;
assign rnode_384to386_bb3_cmp37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_384to386_bb3_cmp37_i_2_NO_SHIFT_REG = rnode_384to386_bb3_cmp37_i_0_reg_386_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_add_i8_stall_local;
wire [31:0] local_bb3_add_i8;

assign local_bb3_add_i8 = ((local_bb3__27_i & 32'h7FFFFF8) | (rnode_383to384_bb3_and36_lobit_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and108_i_stall_local;
wire [31:0] local_bb3_and108_i;

assign local_bb3_and108_i = (local_bb3_cond107_i & local_bb3_or89_i);

// This section implements an unregistered operation.
// 
wire local_bb3__24_i_stall_local;
wire local_bb3__24_i;

assign local_bb3__24_i = (local_bb3_or_cond_not_i | local_bb3_brmerge_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge_not_not_i_stall_local;
wire local_bb3_brmerge_not_not_i;

assign local_bb3_brmerge_not_not_i = (local_bb3_brmerge_not_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_not_cmp37_i_stall_local;
wire local_bb3_not_cmp37_i;

assign local_bb3_not_cmp37_i = (rnode_384to386_bb3_cmp37_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_add192_i_stall_local;
wire [31:0] local_bb3_add192_i;

assign local_bb3_add192_i = ((local_bb3_add_i8 & 32'h7FFFFF9) + rnode_383to384_bb3_xor188_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_or112_i_stall_local;
wire [31:0] local_bb3_or112_i;

assign local_bb3_or112_i = (local_bb3_and108_i | (local_bb3_cond111_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_7_i_stall_local;
wire local_bb3_reduction_7_i;

assign local_bb3_reduction_7_i = (local_bb3_cmp25_i5 & local_bb3_brmerge_not_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u80_valid_out;
wire local_bb3_var__u80_stall_in;
wire local_bb3_var__u80_inputs_ready;
wire local_bb3_var__u80_stall_local;
wire [31:0] local_bb3_var__u80;

assign local_bb3_var__u80_inputs_ready = (rnode_384to385_bb3_xor_i195_0_valid_out_NO_SHIFT_REG & rnode_384to385_bb3__29_i204_0_valid_out_NO_SHIFT_REG & rnode_384to385_bb3_or581_i_0_valid_out_1_NO_SHIFT_REG & rnode_384to385_bb3_or581_i_0_valid_out_0_NO_SHIFT_REG & rnode_384to385_bb3_reduction_0_i212_0_valid_out_NO_SHIFT_REG & rnode_384to385_bb3_cmp68_i_0_valid_out_NO_SHIFT_REG & rnode_384to385_bb3_cmp71_not_i_0_valid_out_NO_SHIFT_REG & rnode_384to385_bb3_shl_i216_0_valid_out_NO_SHIFT_REG & rnode_383to385_bb3_and75_i214_0_valid_out_NO_SHIFT_REG & rnode_384to385_bb3__40_i_0_valid_out_NO_SHIFT_REG);
assign local_bb3_var__u80 = (rnode_384to385_bb3__29_i204_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb3_or112_i);
assign local_bb3_var__u80_valid_out = 1'b1;
assign rnode_384to385_bb3_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_or581_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_or581_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_cmp68_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_cmp71_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_shl_i216_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_383to385_bb3_and75_i214_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3__40_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_9_i_stall_local;
wire local_bb3_reduction_9_i;

assign local_bb3_reduction_9_i = (local_bb3_reduction_7_i & local_bb3_reduction_8_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb3_var__u80_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_var__u80_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_var__u80_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_var__u80_2_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_var__u80_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_valid_out_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_stall_in_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u80_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb3_var__u80_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb3_var__u80_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb3_var__u80_0_stall_in_0_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb3_var__u80_0_valid_out_0_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb3_var__u80_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in(local_bb3_var__u80),
	.data_out(rnode_385to386_bb3_var__u80_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb3_var__u80_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb3_var__u80_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_385to386_bb3_var__u80_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb3_var__u80_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb3_var__u80_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u80_stall_in = 1'b0;
assign rnode_385to386_bb3_var__u80_0_stall_in_0_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_var__u80_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_var__u80_0_NO_SHIFT_REG = rnode_385to386_bb3_var__u80_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_var__u80_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_var__u80_1_NO_SHIFT_REG = rnode_385to386_bb3_var__u80_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_var__u80_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_var__u80_2_NO_SHIFT_REG = rnode_385to386_bb3_var__u80_0_reg_386_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_and17_i_valid_out_2;
wire local_bb3_and17_i_stall_in_2;
wire local_bb3_var__u72_valid_out;
wire local_bb3_var__u72_stall_in;
wire local_bb3_add192_i_valid_out;
wire local_bb3_add192_i_stall_in;
wire local_bb3__26_i_valid_out;
wire local_bb3__26_i_stall_in;
wire local_bb3__26_i_inputs_ready;
wire local_bb3__26_i_stall_local;
wire local_bb3__26_i;

assign local_bb3__26_i_inputs_ready = (rnode_382to384_bb3_shr16_i_0_valid_out_0_NO_SHIFT_REG & rnode_382to384_bb3_cmp27_i_0_valid_out_2_NO_SHIFT_REG & rnode_383to384_bb3_and36_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_383to384_bb3_xor188_i_0_valid_out_NO_SHIFT_REG & rnode_383to384_bb3_and20_i_0_valid_out_0_NO_SHIFT_REG & rnode_382to384_bb3_cmp27_i_0_valid_out_0_NO_SHIFT_REG & rnode_383to384_bb3_lnot33_not_i_0_valid_out_NO_SHIFT_REG & rnode_382to384_bb3_cmp27_i_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb3_and20_i_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb3_cmp37_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3__26_i = (local_bb3_reduction_9_i ? rnode_383to384_bb3_cmp37_i_0_NO_SHIFT_REG : local_bb3__24_i);
assign local_bb3_and17_i_valid_out_2 = 1'b1;
assign local_bb3_var__u72_valid_out = 1'b1;
assign local_bb3_add192_i_valid_out = 1'b1;
assign local_bb3__26_i_valid_out = 1'b1;
assign rnode_382to384_bb3_shr16_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3_cmp27_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and36_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_xor188_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and20_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3_cmp27_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_lnot33_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_382to384_bb3_cmp27_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_and20_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb3_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and_i11_stall_local;
wire [31:0] local_bb3_and_i11;

assign local_bb3_and_i11 = (rnode_385to386_bb3_var__u80_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and10_i17_stall_local;
wire [31:0] local_bb3_and10_i17;

assign local_bb3_and10_i17 = (rnode_385to386_bb3_var__u80_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_var__u80_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u80_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_var__u80_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u80_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u80_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_var__u80_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u80_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_var__u80_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u80_0_valid_out_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u80_0_stall_in_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u80_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_var__u80_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_var__u80_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_var__u80_0_stall_in_0_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_var__u80_0_valid_out_0_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_var__u80_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_385to386_bb3_var__u80_2_NO_SHIFT_REG),
	.data_out(rnode_386to387_bb3_var__u80_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_var__u80_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_var__u80_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb3_var__u80_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_var__u80_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_var__u80_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_var__u80_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u80_0_stall_in_0_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u80_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3_var__u80_0_NO_SHIFT_REG = rnode_386to387_bb3_var__u80_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_var__u80_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3_var__u80_1_NO_SHIFT_REG = rnode_386to387_bb3_var__u80_0_reg_387_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_384to386_bb3_and17_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and17_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_384to386_bb3_and17_i_0_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and17_i_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to386_bb3_and17_i_0_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and17_i_0_valid_out_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and17_i_0_stall_in_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb3_and17_i_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_384to386_bb3_and17_i_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to386_bb3_and17_i_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to386_bb3_and17_i_0_stall_in_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_384to386_bb3_and17_i_0_valid_out_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_384to386_bb3_and17_i_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((local_bb3_and17_i & 32'hFF)),
	.data_out(rnode_384to386_bb3_and17_i_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_384to386_bb3_and17_i_0_reg_386_fifo.DEPTH = 2;
defparam rnode_384to386_bb3_and17_i_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_384to386_bb3_and17_i_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to386_bb3_and17_i_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_384to386_bb3_and17_i_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and17_i_stall_in_2 = 1'b0;
assign rnode_384to386_bb3_and17_i_0_NO_SHIFT_REG = rnode_384to386_bb3_and17_i_0_reg_386_NO_SHIFT_REG;
assign rnode_384to386_bb3_and17_i_0_stall_in_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_and17_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_var__u72_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3_var__u72_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb3_var__u72_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_var__u72_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3_var__u72_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_var__u72_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_var__u72_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_var__u72_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_var__u72_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_var__u72_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_var__u72_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_var__u72_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_var__u72_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb3_var__u72),
	.data_out(rnode_384to385_bb3_var__u72_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_var__u72_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_var__u72_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3_var__u72_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_var__u72_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_var__u72_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u72_stall_in = 1'b0;
assign rnode_384to385_bb3_var__u72_0_NO_SHIFT_REG = rnode_384to385_bb3_var__u72_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_var__u72_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_var__u72_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3_add192_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_add192_i_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_add192_i_1_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_add192_i_2_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_add192_i_3_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb3_add192_i_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_valid_out_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_stall_in_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3_add192_i_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3_add192_i_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3_add192_i_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3_add192_i_0_stall_in_0_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3_add192_i_0_valid_out_0_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3_add192_i_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb3_add192_i),
	.data_out(rnode_384to385_bb3_add192_i_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3_add192_i_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3_add192_i_0_reg_385_fifo.DATA_WIDTH = 32;
defparam rnode_384to385_bb3_add192_i_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3_add192_i_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3_add192_i_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add192_i_stall_in = 1'b0;
assign rnode_384to385_bb3_add192_i_0_stall_in_0_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3_add192_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3_add192_i_0_NO_SHIFT_REG = rnode_384to385_bb3_add192_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_add192_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3_add192_i_1_NO_SHIFT_REG = rnode_384to385_bb3_add192_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_add192_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3_add192_i_2_NO_SHIFT_REG = rnode_384to385_bb3_add192_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3_add192_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3_add192_i_3_NO_SHIFT_REG = rnode_384to385_bb3_add192_i_0_reg_385_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb3__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb3__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb3__26_i_0_NO_SHIFT_REG;
 logic rnode_384to385_bb3__26_i_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb3__26_i_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__26_i_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__26_i_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb3__26_i_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb3__26_i_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb3__26_i_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb3__26_i_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb3__26_i_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb3__26_i_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb3__26_i),
	.data_out(rnode_384to385_bb3__26_i_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb3__26_i_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb3__26_i_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb3__26_i_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb3__26_i_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb3__26_i_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__26_i_stall_in = 1'b0;
assign rnode_384to385_bb3__26_i_0_NO_SHIFT_REG = rnode_384to385_bb3__26_i_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb3__26_i_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb3__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i12_stall_local;
wire [31:0] local_bb3_shr_i12;

assign local_bb3_shr_i12 = ((local_bb3_and_i11 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp13_i19_stall_local;
wire local_bb3_cmp13_i19;

assign local_bb3_cmp13_i19 = ((local_bb3_and10_i17 & 32'hFFFF) > (local_bb3_and12_i18 & 32'hFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb3_var__u72_0_valid_out_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u72_0_stall_in_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u72_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u72_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u72_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u72_0_valid_out_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u72_0_stall_in_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_var__u72_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb3_var__u72_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb3_var__u72_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb3_var__u72_0_stall_in_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb3_var__u72_0_valid_out_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb3_var__u72_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in(rnode_384to385_bb3_var__u72_0_NO_SHIFT_REG),
	.data_out(rnode_385to386_bb3_var__u72_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb3_var__u72_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb3_var__u72_0_reg_386_fifo.DATA_WIDTH = 1;
defparam rnode_385to386_bb3_var__u72_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb3_var__u72_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb3_var__u72_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3_var__u72_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_var__u72_0_NO_SHIFT_REG = rnode_385to386_bb3_var__u72_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_var__u72_0_stall_in_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_var__u72_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and193_i_valid_out;
wire local_bb3_and193_i_stall_in;
wire local_bb3_and193_i_inputs_ready;
wire local_bb3_and193_i_stall_local;
wire [31:0] local_bb3_and193_i;

assign local_bb3_and193_i_inputs_ready = rnode_384to385_bb3_add192_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_and193_i = (rnode_384to385_bb3_add192_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb3_and193_i_valid_out = 1'b1;
assign rnode_384to385_bb3_add192_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and195_i_valid_out;
wire local_bb3_and195_i_stall_in;
wire local_bb3_and195_i_inputs_ready;
wire local_bb3_and195_i_stall_local;
wire [31:0] local_bb3_and195_i;

assign local_bb3_and195_i_inputs_ready = rnode_384to385_bb3_add192_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_and195_i = (rnode_384to385_bb3_add192_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb3_and195_i_valid_out = 1'b1;
assign rnode_384to385_bb3_add192_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and198_i_valid_out;
wire local_bb3_and198_i_stall_in;
wire local_bb3_and198_i_inputs_ready;
wire local_bb3_and198_i_stall_local;
wire [31:0] local_bb3_and198_i;

assign local_bb3_and198_i_inputs_ready = rnode_384to385_bb3_add192_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_and198_i = (rnode_384to385_bb3_add192_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb3_and198_i_valid_out = 1'b1;
assign rnode_384to385_bb3_add192_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and201_i_stall_local;
wire [31:0] local_bb3_and201_i;

assign local_bb3_and201_i = (rnode_384to385_bb3_add192_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_385to387_bb3__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_385to387_bb3__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_385to387_bb3__26_i_0_NO_SHIFT_REG;
 logic rnode_385to387_bb3__26_i_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_385to387_bb3__26_i_0_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb3__26_i_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb3__26_i_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb3__26_i_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_385to387_bb3__26_i_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to387_bb3__26_i_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to387_bb3__26_i_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_385to387_bb3__26_i_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_385to387_bb3__26_i_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_384to385_bb3__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_385to387_bb3__26_i_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_385to387_bb3__26_i_0_reg_387_fifo.DEPTH = 2;
defparam rnode_385to387_bb3__26_i_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_385to387_bb3__26_i_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to387_bb3__26_i_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_385to387_bb3__26_i_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb3__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to387_bb3__26_i_0_NO_SHIFT_REG = rnode_385to387_bb3__26_i_0_reg_387_NO_SHIFT_REG;
assign rnode_385to387_bb3__26_i_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_385to387_bb3__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i15_stall_local;
wire local_bb3_cmp_i15;

assign local_bb3_cmp_i15 = ((local_bb3_shr_i12 & 32'h7FFF) > (local_bb3_shr3_i14 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp8_i16_stall_local;
wire local_bb3_cmp8_i16;

assign local_bb3_cmp8_i16 = ((local_bb3_shr_i12 & 32'h7FFF) == (local_bb3_shr3_i14 & 32'h7FFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_var__u72_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u72_0_stall_in_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u72_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u72_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u72_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u72_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u72_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u72_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_var__u72_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_var__u72_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_var__u72_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_var__u72_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_var__u72_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_385to386_bb3_var__u72_0_NO_SHIFT_REG),
	.data_out(rnode_386to387_bb3_var__u72_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_var__u72_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_var__u72_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_386to387_bb3_var__u72_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_var__u72_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_var__u72_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_var__u72_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u72_0_NO_SHIFT_REG = rnode_386to387_bb3_var__u72_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_var__u72_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u72_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb3_and193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and193_i_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and193_i_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and193_i_2_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and193_i_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_valid_out_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_stall_in_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and193_i_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb3_and193_i_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb3_and193_i_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb3_and193_i_0_stall_in_0_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb3_and193_i_0_valid_out_0_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb3_and193_i_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((local_bb3_and193_i & 32'hFFFFFFF)),
	.data_out(rnode_385to386_bb3_and193_i_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb3_and193_i_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb3_and193_i_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_385to386_bb3_and193_i_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb3_and193_i_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb3_and193_i_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and193_i_stall_in = 1'b0;
assign rnode_385to386_bb3_and193_i_0_stall_in_0_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_and193_i_0_NO_SHIFT_REG = rnode_385to386_bb3_and193_i_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_and193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_and193_i_1_NO_SHIFT_REG = rnode_385to386_bb3_and193_i_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_and193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3_and193_i_2_NO_SHIFT_REG = rnode_385to386_bb3_and193_i_0_reg_386_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb3_and195_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and195_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and195_i_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and195_i_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and195_i_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and195_i_0_valid_out_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and195_i_0_stall_in_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and195_i_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb3_and195_i_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb3_and195_i_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb3_and195_i_0_stall_in_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb3_and195_i_0_valid_out_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb3_and195_i_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((local_bb3_and195_i & 32'h1F)),
	.data_out(rnode_385to386_bb3_and195_i_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb3_and195_i_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb3_and195_i_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_385to386_bb3_and195_i_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb3_and195_i_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb3_and195_i_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and195_i_stall_in = 1'b0;
assign rnode_385to386_bb3_and195_i_0_NO_SHIFT_REG = rnode_385to386_bb3_and195_i_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_and195_i_0_stall_in_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and195_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb3_and198_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and198_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and198_i_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and198_i_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3_and198_i_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and198_i_0_valid_out_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and198_i_0_stall_in_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3_and198_i_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb3_and198_i_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb3_and198_i_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb3_and198_i_0_stall_in_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb3_and198_i_0_valid_out_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb3_and198_i_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((local_bb3_and198_i & 32'h1)),
	.data_out(rnode_385to386_bb3_and198_i_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb3_and198_i_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb3_and198_i_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_385to386_bb3_and198_i_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb3_and198_i_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb3_and198_i_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and198_i_stall_in = 1'b0;
assign rnode_385to386_bb3_and198_i_0_NO_SHIFT_REG = rnode_385to386_bb3_and198_i_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3_and198_i_0_stall_in_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and198_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i_i_stall_local;
wire [31:0] local_bb3_shr_i_i;

assign local_bb3_shr_i_i = ((local_bb3_and201_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3__26_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__26_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3__26_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3__26_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3__26_i_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3__26_i_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3__26_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_385to387_bb3__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb3__26_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3__26_i_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3__26_i_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb3__26_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3__26_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3__26_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_385to387_bb3__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__26_i_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__26_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__26_i_0_NO_SHIFT_REG = rnode_387to388_bb3__26_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3__26_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__26_i_1_NO_SHIFT_REG = rnode_387to388_bb3__26_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3__26_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__26_i_2_NO_SHIFT_REG = rnode_387to388_bb3__26_i_0_reg_388_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3___i20_stall_local;
wire local_bb3___i20;

assign local_bb3___i20 = (local_bb3_cmp8_i16 & local_bb3_cmp13_i19);

// This section implements an unregistered operation.
// 
wire local_bb3_shr216_i_stall_local;
wire [31:0] local_bb3_shr216_i;

assign local_bb3_shr216_i = ((rnode_385to386_bb3_and193_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__pre_i_stall_local;
wire [31:0] local_bb3__pre_i;

assign local_bb3__pre_i = ((rnode_385to386_bb3_and195_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i_i_stall_local;
wire [31:0] local_bb3_or_i_i;

assign local_bb3_or_i_i = ((local_bb3_shr_i_i & 32'h3FFFFFF) | (local_bb3_and201_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cond292_i_stall_local;
wire [31:0] local_bb3_cond292_i;

assign local_bb3_cond292_i = (rnode_387to388_bb3__26_i_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u81_stall_local;
wire [31:0] local_bb3_var__u81;

assign local_bb3_var__u81[31:1] = 31'h0;
assign local_bb3_var__u81[0] = rnode_387to388_bb3__26_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u20_valid_out_2;
wire local_bb3_var__u20_stall_in_2;
wire local_bb3__21_i21_valid_out;
wire local_bb3__21_i21_stall_in;
wire local_bb3__21_i21_inputs_ready;
wire local_bb3__21_i21_stall_local;
wire local_bb3__21_i21;

assign local_bb3__21_i21_inputs_ready = (rnode_385to386_bb3_c0_ene5_0_valid_out_0_NO_SHIFT_REG & rnode_385to386_bb3_var__u80_0_valid_out_1_NO_SHIFT_REG & rnode_385to386_bb3_var__u80_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3__21_i21 = (local_bb3_cmp_i15 | local_bb3___i20);
assign local_bb3_var__u20_valid_out_2 = 1'b1;
assign local_bb3__21_i21_valid_out = 1'b1;
assign rnode_385to386_bb3_c0_ene5_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_var__u80_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_var__u80_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_or219_i_stall_local;
wire [31:0] local_bb3_or219_i;

assign local_bb3_or219_i = ((local_bb3_shr216_i & 32'h7FFFFFF) | (rnode_385to386_bb3_and198_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool213_i_stall_local;
wire local_bb3_tobool213_i;

assign local_bb3_tobool213_i = ((local_bb3__pre_i & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_shr1_i_i_stall_local;
wire [31:0] local_bb3_shr1_i_i;

assign local_bb3_shr1_i_i = ((local_bb3_or_i_i & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext_i_stall_local;
wire [31:0] local_bb3_lnot_ext_i;

assign local_bb3_lnot_ext_i = ((local_bb3_var__u81 & 32'h1) ^ 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_var__u20_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u20_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_var__u20_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u20_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u20_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_var__u20_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u20_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_var__u20_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u20_0_valid_out_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u20_0_stall_in_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_var__u20_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_var__u20_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_var__u20_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_var__u20_0_stall_in_0_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_var__u20_0_valid_out_0_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_var__u20_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(local_bb3_var__u20),
	.data_out(rnode_386to387_bb3_var__u20_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_var__u20_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_var__u20_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb3_var__u20_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_var__u20_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_var__u20_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u20_stall_in_2 = 1'b0;
assign rnode_386to387_bb3_var__u20_0_stall_in_0_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u20_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3_var__u20_0_NO_SHIFT_REG = rnode_386to387_bb3_var__u20_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_var__u20_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3_var__u20_1_NO_SHIFT_REG = rnode_386to387_bb3_var__u20_0_reg_387_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3__21_i21_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_valid_out_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_stall_in_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3__21_i21_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3__21_i21_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3__21_i21_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3__21_i21_0_stall_in_0_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3__21_i21_0_valid_out_0_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3__21_i21_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(local_bb3__21_i21),
	.data_out(rnode_386to387_bb3__21_i21_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3__21_i21_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3__21_i21_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_386to387_bb3__21_i21_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3__21_i21_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3__21_i21_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__21_i21_stall_in = 1'b0;
assign rnode_386to387_bb3__21_i21_0_stall_in_0_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3__21_i21_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3__21_i21_0_NO_SHIFT_REG = rnode_386to387_bb3__21_i21_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3__21_i21_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3__21_i21_1_NO_SHIFT_REG = rnode_386to387_bb3__21_i21_0_reg_387_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__40_demorgan_i_stall_local;
wire local_bb3__40_demorgan_i;

assign local_bb3__40_demorgan_i = (rnode_384to386_bb3_cmp37_i_0_NO_SHIFT_REG | local_bb3_tobool213_i);

// This section implements an unregistered operation.
// 
wire local_bb3__42_i_stall_local;
wire local_bb3__42_i;

assign local_bb3__42_i = (local_bb3_tobool213_i & local_bb3_not_cmp37_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or2_i_i_stall_local;
wire [31:0] local_bb3_or2_i_i;

assign local_bb3_or2_i_i = ((local_bb3_shr1_i_i & 32'h1FFFFFF) | (local_bb3_or_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__22_i22_stall_local;
wire [31:0] local_bb3__22_i22;

assign local_bb3__22_i22 = (rnode_386to387_bb3__21_i21_0_NO_SHIFT_REG ? rnode_386to387_bb3_var__u20_0_NO_SHIFT_REG : rnode_386to387_bb3_var__u80_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3__23_i23_stall_local;
wire [31:0] local_bb3__23_i23;

assign local_bb3__23_i23 = (rnode_386to387_bb3__21_i21_1_NO_SHIFT_REG ? rnode_386to387_bb3_var__u80_1_NO_SHIFT_REG : rnode_386to387_bb3_var__u20_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3__43_i_stall_local;
wire [31:0] local_bb3__43_i;

assign local_bb3__43_i = (local_bb3__42_i ? 32'h0 : (local_bb3__pre_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_shr3_i_i_stall_local;
wire [31:0] local_bb3_shr3_i_i;

assign local_bb3_shr3_i_i = ((local_bb3_or2_i_i & 32'h7FFFFFF) >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb3_shr18_i26_stall_local;
wire [31:0] local_bb3_shr18_i26;

assign local_bb3_shr18_i26 = (local_bb3__22_i22 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_shr16_i24_stall_local;
wire [31:0] local_bb3_shr16_i24;

assign local_bb3_shr16_i24 = (local_bb3__23_i23 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_or4_i_i_stall_local;
wire [31:0] local_bb3_or4_i_i;

assign local_bb3_or4_i_i = ((local_bb3_shr3_i_i & 32'h7FFFFF) | (local_bb3_or2_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_and19_i27_stall_local;
wire [31:0] local_bb3_and19_i27;

assign local_bb3_and19_i27 = ((local_bb3_shr18_i26 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_sub_i56_stall_local;
wire [31:0] local_bb3_sub_i56;

assign local_bb3_sub_i56 = ((local_bb3_shr16_i24 & 32'h1FF) - (local_bb3_shr18_i26 & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb3_shr5_i_i_stall_local;
wire [31:0] local_bb3_shr5_i_i;

assign local_bb3_shr5_i_i = ((local_bb3_or4_i_i & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot23_i31_stall_local;
wire local_bb3_lnot23_i31;

assign local_bb3_lnot23_i31 = ((local_bb3_and19_i27 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp27_i33_stall_local;
wire local_bb3_cmp27_i33;

assign local_bb3_cmp27_i33 = ((local_bb3_and19_i27 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and68_i57_stall_local;
wire [31:0] local_bb3_and68_i57;

assign local_bb3_and68_i57 = (local_bb3_sub_i56 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_or6_i_i_stall_local;
wire [31:0] local_bb3_or6_i_i;

assign local_bb3_or6_i_i = ((local_bb3_shr5_i_i & 32'h7FFFF) | (local_bb3_or4_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cmp69_i58_stall_local;
wire local_bb3_cmp69_i58;

assign local_bb3_cmp69_i58 = ((local_bb3_and68_i57 & 32'hFF) > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_shr7_i_i_stall_local;
wire [31:0] local_bb3_shr7_i_i;

assign local_bb3_shr7_i_i = ((local_bb3_or6_i_i & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_or6_masked_i_i_stall_local;
wire [31:0] local_bb3_or6_masked_i_i;

assign local_bb3_or6_masked_i_i = ((local_bb3_or6_i_i & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3__22_i22_valid_out_1;
wire local_bb3__22_i22_stall_in_1;
wire local_bb3__23_i23_valid_out_1;
wire local_bb3__23_i23_stall_in_1;
wire local_bb3_shr16_i24_valid_out_1;
wire local_bb3_shr16_i24_stall_in_1;
wire local_bb3_lnot23_i31_valid_out;
wire local_bb3_lnot23_i31_stall_in;
wire local_bb3_cmp27_i33_valid_out;
wire local_bb3_cmp27_i33_stall_in;
wire local_bb3_align_0_i59_valid_out;
wire local_bb3_align_0_i59_stall_in;
wire local_bb3_align_0_i59_inputs_ready;
wire local_bb3_align_0_i59_stall_local;
wire [31:0] local_bb3_align_0_i59;

assign local_bb3_align_0_i59_inputs_ready = (rnode_386to387_bb3__21_i21_0_valid_out_0_NO_SHIFT_REG & rnode_386to387_bb3_var__u20_0_valid_out_0_NO_SHIFT_REG & rnode_386to387_bb3_var__u80_0_valid_out_0_NO_SHIFT_REG & rnode_386to387_bb3__21_i21_0_valid_out_1_NO_SHIFT_REG & rnode_386to387_bb3_var__u20_0_valid_out_1_NO_SHIFT_REG & rnode_386to387_bb3_var__u80_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_align_0_i59 = (local_bb3_cmp69_i58 ? 32'h1F : (local_bb3_and68_i57 & 32'hFF));
assign local_bb3__22_i22_valid_out_1 = 1'b1;
assign local_bb3__23_i23_valid_out_1 = 1'b1;
assign local_bb3_shr16_i24_valid_out_1 = 1'b1;
assign local_bb3_lnot23_i31_valid_out = 1'b1;
assign local_bb3_cmp27_i33_valid_out = 1'b1;
assign local_bb3_align_0_i59_valid_out = 1'b1;
assign rnode_386to387_bb3__21_i21_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u20_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u80_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3__21_i21_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u20_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u80_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_neg_i_i_stall_local;
wire [31:0] local_bb3_neg_i_i;

assign local_bb3_neg_i_i = ((local_bb3_or6_masked_i_i & 32'h7FFFFFF) | (local_bb3_shr7_i_i & 32'h7FF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3__22_i22_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__22_i22_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3__22_i22_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__22_i22_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__22_i22_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3__22_i22_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__22_i22_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3__22_i22_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__22_i22_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__22_i22_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__22_i22_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3__22_i22_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3__22_i22_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3__22_i22_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3__22_i22_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3__22_i22_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb3__22_i22),
	.data_out(rnode_387to388_bb3__22_i22_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3__22_i22_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3__22_i22_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb3__22_i22_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3__22_i22_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3__22_i22_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__22_i22_stall_in_1 = 1'b0;
assign rnode_387to388_bb3__22_i22_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__22_i22_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__22_i22_0_NO_SHIFT_REG = rnode_387to388_bb3__22_i22_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3__22_i22_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__22_i22_1_NO_SHIFT_REG = rnode_387to388_bb3__22_i22_0_reg_388_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3__23_i23_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3__23_i23_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3__23_i23_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3__23_i23_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3__23_i23_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__23_i23_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3__23_i23_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3__23_i23_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3__23_i23_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3__23_i23_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3__23_i23_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb3__23_i23),
	.data_out(rnode_387to388_bb3__23_i23_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3__23_i23_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3__23_i23_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb3__23_i23_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3__23_i23_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3__23_i23_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__23_i23_stall_in_1 = 1'b0;
assign rnode_387to388_bb3__23_i23_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__23_i23_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__23_i23_0_NO_SHIFT_REG = rnode_387to388_bb3__23_i23_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3__23_i23_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__23_i23_1_NO_SHIFT_REG = rnode_387to388_bb3__23_i23_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3__23_i23_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__23_i23_2_NO_SHIFT_REG = rnode_387to388_bb3__23_i23_0_reg_388_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_387to389_bb3_shr16_i24_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to389_bb3_shr16_i24_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_387to389_bb3_shr16_i24_0_NO_SHIFT_REG;
 logic rnode_387to389_bb3_shr16_i24_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to389_bb3_shr16_i24_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_387to389_bb3_shr16_i24_1_NO_SHIFT_REG;
 logic rnode_387to389_bb3_shr16_i24_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to389_bb3_shr16_i24_0_reg_389_NO_SHIFT_REG;
 logic rnode_387to389_bb3_shr16_i24_0_valid_out_0_reg_389_NO_SHIFT_REG;
 logic rnode_387to389_bb3_shr16_i24_0_stall_in_0_reg_389_NO_SHIFT_REG;
 logic rnode_387to389_bb3_shr16_i24_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_387to389_bb3_shr16_i24_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to389_bb3_shr16_i24_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to389_bb3_shr16_i24_0_stall_in_0_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_387to389_bb3_shr16_i24_0_valid_out_0_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_387to389_bb3_shr16_i24_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb3_shr16_i24 & 32'h1FF)),
	.data_out(rnode_387to389_bb3_shr16_i24_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_387to389_bb3_shr16_i24_0_reg_389_fifo.DEPTH = 2;
defparam rnode_387to389_bb3_shr16_i24_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_387to389_bb3_shr16_i24_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to389_bb3_shr16_i24_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_387to389_bb3_shr16_i24_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr16_i24_stall_in_1 = 1'b0;
assign rnode_387to389_bb3_shr16_i24_0_stall_in_0_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_387to389_bb3_shr16_i24_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to389_bb3_shr16_i24_0_NO_SHIFT_REG = rnode_387to389_bb3_shr16_i24_0_reg_389_NO_SHIFT_REG;
assign rnode_387to389_bb3_shr16_i24_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to389_bb3_shr16_i24_1_NO_SHIFT_REG = rnode_387to389_bb3_shr16_i24_0_reg_389_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_lnot23_i31_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb3_lnot23_i31_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb3_lnot23_i31_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_lnot23_i31_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb3_lnot23_i31_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_lnot23_i31_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_lnot23_i31_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_lnot23_i31_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_lnot23_i31_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_lnot23_i31_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_lnot23_i31_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_lnot23_i31_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_lnot23_i31_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb3_lnot23_i31),
	.data_out(rnode_387to388_bb3_lnot23_i31_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_lnot23_i31_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_lnot23_i31_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb3_lnot23_i31_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_lnot23_i31_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_lnot23_i31_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_lnot23_i31_stall_in = 1'b0;
assign rnode_387to388_bb3_lnot23_i31_0_NO_SHIFT_REG = rnode_387to388_bb3_lnot23_i31_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_lnot23_i31_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_lnot23_i31_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_387to389_bb3_cmp27_i33_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_1_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_2_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_reg_389_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_valid_out_0_reg_389_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_stall_in_0_reg_389_NO_SHIFT_REG;
 logic rnode_387to389_bb3_cmp27_i33_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_387to389_bb3_cmp27_i33_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to389_bb3_cmp27_i33_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to389_bb3_cmp27_i33_0_stall_in_0_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_387to389_bb3_cmp27_i33_0_valid_out_0_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_387to389_bb3_cmp27_i33_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb3_cmp27_i33),
	.data_out(rnode_387to389_bb3_cmp27_i33_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_387to389_bb3_cmp27_i33_0_reg_389_fifo.DEPTH = 2;
defparam rnode_387to389_bb3_cmp27_i33_0_reg_389_fifo.DATA_WIDTH = 1;
defparam rnode_387to389_bb3_cmp27_i33_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to389_bb3_cmp27_i33_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_387to389_bb3_cmp27_i33_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp27_i33_stall_in = 1'b0;
assign rnode_387to389_bb3_cmp27_i33_0_stall_in_0_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_387to389_bb3_cmp27_i33_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to389_bb3_cmp27_i33_0_NO_SHIFT_REG = rnode_387to389_bb3_cmp27_i33_0_reg_389_NO_SHIFT_REG;
assign rnode_387to389_bb3_cmp27_i33_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to389_bb3_cmp27_i33_1_NO_SHIFT_REG = rnode_387to389_bb3_cmp27_i33_0_reg_389_NO_SHIFT_REG;
assign rnode_387to389_bb3_cmp27_i33_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_387to389_bb3_cmp27_i33_2_NO_SHIFT_REG = rnode_387to389_bb3_cmp27_i33_0_reg_389_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_align_0_i59_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_align_0_i59_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_align_0_i59_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_align_0_i59_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_align_0_i59_3_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_align_0_i59_4_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_align_0_i59_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_align_0_i59_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_align_0_i59_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_align_0_i59_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_align_0_i59_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_align_0_i59_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_align_0_i59_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in((local_bb3_align_0_i59 & 32'hFF)),
	.data_out(rnode_387to388_bb3_align_0_i59_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_align_0_i59_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_align_0_i59_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb3_align_0_i59_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_align_0_i59_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_align_0_i59_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_align_0_i59_stall_in = 1'b0;
assign rnode_387to388_bb3_align_0_i59_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_align_0_i59_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_align_0_i59_0_NO_SHIFT_REG = rnode_387to388_bb3_align_0_i59_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_align_0_i59_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_align_0_i59_1_NO_SHIFT_REG = rnode_387to388_bb3_align_0_i59_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_align_0_i59_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_align_0_i59_2_NO_SHIFT_REG = rnode_387to388_bb3_align_0_i59_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_align_0_i59_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_align_0_i59_3_NO_SHIFT_REG = rnode_387to388_bb3_align_0_i59_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_align_0_i59_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_align_0_i59_4_NO_SHIFT_REG = rnode_387to388_bb3_align_0_i59_0_reg_388_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_and_i_i9_stall_local;
wire [31:0] local_bb3_and_i_i9;

assign local_bb3_and_i_i9 = ((local_bb3_neg_i_i & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and21_i29_stall_local;
wire [31:0] local_bb3_and21_i29;

assign local_bb3_and21_i29 = (rnode_387to388_bb3__22_i22_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and20_i28_valid_out;
wire local_bb3_and20_i28_stall_in;
wire local_bb3_and20_i28_inputs_ready;
wire local_bb3_and20_i28_stall_local;
wire [31:0] local_bb3_and20_i28;

assign local_bb3_and20_i28_inputs_ready = rnode_387to388_bb3__23_i23_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_and20_i28 = (rnode_387to388_bb3__23_i23_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb3_and20_i28_valid_out = 1'b1;
assign rnode_387to388_bb3__23_i23_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and35_i34_valid_out;
wire local_bb3_and35_i34_stall_in;
wire local_bb3_and35_i34_inputs_ready;
wire local_bb3_and35_i34_stall_local;
wire [31:0] local_bb3_and35_i34;

assign local_bb3_and35_i34_inputs_ready = rnode_387to388_bb3__23_i23_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_and35_i34 = (rnode_387to388_bb3__23_i23_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb3_and35_i34_valid_out = 1'b1;
assign rnode_387to388_bb3__23_i23_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_xor_i35_stall_local;
wire [31:0] local_bb3_xor_i35;

assign local_bb3_xor_i35 = (rnode_387to388_bb3__23_i23_2_NO_SHIFT_REG ^ rnode_387to388_bb3__22_i22_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_and17_i25_stall_local;
wire [31:0] local_bb3_and17_i25;

assign local_bb3_and17_i25 = ((rnode_387to389_bb3_shr16_i24_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_389to391_bb3_shr16_i24_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to391_bb3_shr16_i24_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb3_shr16_i24_0_NO_SHIFT_REG;
 logic rnode_389to391_bb3_shr16_i24_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb3_shr16_i24_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_shr16_i24_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_shr16_i24_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_shr16_i24_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_389to391_bb3_shr16_i24_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to391_bb3_shr16_i24_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to391_bb3_shr16_i24_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_389to391_bb3_shr16_i24_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_389to391_bb3_shr16_i24_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((rnode_387to389_bb3_shr16_i24_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_389to391_bb3_shr16_i24_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_389to391_bb3_shr16_i24_0_reg_391_fifo.DEPTH = 2;
defparam rnode_389to391_bb3_shr16_i24_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_389to391_bb3_shr16_i24_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to391_bb3_shr16_i24_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_389to391_bb3_shr16_i24_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_387to389_bb3_shr16_i24_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_shr16_i24_0_NO_SHIFT_REG = rnode_389to391_bb3_shr16_i24_0_reg_391_NO_SHIFT_REG;
assign rnode_389to391_bb3_shr16_i24_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_shr16_i24_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and93_i67_stall_local;
wire [31:0] local_bb3_and93_i67;

assign local_bb3_and93_i67 = ((rnode_387to388_bb3_align_0_i59_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb3_and95_i69_stall_local;
wire [31:0] local_bb3_and95_i69;

assign local_bb3_and95_i69 = ((rnode_387to388_bb3_align_0_i59_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_and115_i85_stall_local;
wire [31:0] local_bb3_and115_i85;

assign local_bb3_and115_i85 = ((rnode_387to388_bb3_align_0_i59_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_and130_i91_stall_local;
wire [31:0] local_bb3_and130_i91;

assign local_bb3_and130_i91 = ((rnode_387to388_bb3_align_0_i59_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb3_and149_i96_stall_local;
wire [31:0] local_bb3_and149_i96;

assign local_bb3_and149_i96 = ((rnode_387to388_bb3_align_0_i59_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb3__and_i_i9_valid_out;
wire local_bb3__and_i_i9_stall_in;
wire local_bb3__and_i_i9_inputs_ready;
wire local_bb3__and_i_i9_stall_local;
wire [31:0] local_bb3__and_i_i9;

thirtysix_six_comp local_bb3__and_i_i9_popcnt_instance (
	.data((local_bb3_and_i_i9 & 32'h7FFFFFF)),
	.sum(local_bb3__and_i_i9)
);


assign local_bb3__and_i_i9_inputs_ready = rnode_384to385_bb3_add192_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb3__and_i_i9_valid_out = 1'b1;
assign rnode_384to385_bb3_add192_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_lnot33_not_i40_stall_local;
wire local_bb3_lnot33_not_i40;

assign local_bb3_lnot33_not_i40 = ((local_bb3_and21_i29 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or64_i53_stall_local;
wire [31:0] local_bb3_or64_i53;

assign local_bb3_or64_i53 = ((local_bb3_and21_i29 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3_and20_i28_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and20_i28_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_and20_i28_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and20_i28_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and20_i28_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_and20_i28_1_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and20_i28_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_and20_i28_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and20_i28_0_valid_out_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and20_i28_0_stall_in_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and20_i28_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3_and20_i28_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3_and20_i28_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3_and20_i28_0_stall_in_0_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3_and20_i28_0_valid_out_0_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3_and20_i28_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb3_and20_i28 & 32'h7FFFFF)),
	.data_out(rnode_388to389_bb3_and20_i28_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3_and20_i28_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3_and20_i28_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb3_and20_i28_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3_and20_i28_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3_and20_i28_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and20_i28_stall_in = 1'b0;
assign rnode_388to389_bb3_and20_i28_0_stall_in_0_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_and20_i28_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3_and20_i28_0_NO_SHIFT_REG = rnode_388to389_bb3_and20_i28_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3_and20_i28_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3_and20_i28_1_NO_SHIFT_REG = rnode_388to389_bb3_and20_i28_0_reg_389_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_and35_i34_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and35_i34_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_and35_i34_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and35_i34_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and35_i34_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and35_i34_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3_and35_i34_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3_and35_i34_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3_and35_i34_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3_and35_i34_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3_and35_i34_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb3_and35_i34 & 32'h80000000)),
	.data_out(rnode_388to389_bb3_and35_i34_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3_and35_i34_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3_and35_i34_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb3_and35_i34_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3_and35_i34_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3_and35_i34_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and35_i34_stall_in = 1'b0;
assign rnode_388to389_bb3_and35_i34_0_NO_SHIFT_REG = rnode_388to389_bb3_and35_i34_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3_and35_i34_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp37_i36_stall_local;
wire local_bb3_cmp37_i36;

assign local_bb3_cmp37_i36 = ($signed(local_bb3_xor_i35) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb3_xor_lobit_i109_stall_local;
wire [31:0] local_bb3_xor_lobit_i109;

assign local_bb3_xor_lobit_i109 = ($signed(local_bb3_xor_i35) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_and36_lobit_i111_stall_local;
wire [31:0] local_bb3_and36_lobit_i111;

assign local_bb3_and36_lobit_i111 = (local_bb3_xor_i35 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_i30_stall_local;
wire local_bb3_lnot_i30;

assign local_bb3_lnot_i30 = ((local_bb3_and17_i25 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_i32_stall_local;
wire local_bb3_cmp25_i32;

assign local_bb3_cmp25_i32 = ((local_bb3_and17_i25 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp96_i70_stall_local;
wire local_bb3_cmp96_i70;

assign local_bb3_cmp96_i70 = ((local_bb3_and95_i69 & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp116_i86_stall_local;
wire local_bb3_cmp116_i86;

assign local_bb3_cmp116_i86 = ((local_bb3_and115_i85 & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp131_not_i93_stall_local;
wire local_bb3_cmp131_not_i93;

assign local_bb3_cmp131_not_i93 = ((local_bb3_and130_i91 & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_Pivot20_i98_stall_local;
wire local_bb3_Pivot20_i98;

assign local_bb3_Pivot20_i98 = ((local_bb3_and149_i96 & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_SwitchLeaf_i99_stall_local;
wire local_bb3_SwitchLeaf_i99;

assign local_bb3_SwitchLeaf_i99 = ((local_bb3_and149_i96 & 32'h3) == 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb3__and_i_i9_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3__and_i_i9_0_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3__and_i_i9_1_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3__and_i_i9_2_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb3__and_i_i9_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_valid_out_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_stall_in_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb3__and_i_i9_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb3__and_i_i9_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb3__and_i_i9_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb3__and_i_i9_0_stall_in_0_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb3__and_i_i9_0_valid_out_0_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb3__and_i_i9_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((local_bb3__and_i_i9 & 32'h3F)),
	.data_out(rnode_385to386_bb3__and_i_i9_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb3__and_i_i9_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb3__and_i_i9_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_385to386_bb3__and_i_i9_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb3__and_i_i9_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb3__and_i_i9_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__and_i_i9_stall_in = 1'b0;
assign rnode_385to386_bb3__and_i_i9_0_stall_in_0_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3__and_i_i9_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3__and_i_i9_0_NO_SHIFT_REG = rnode_385to386_bb3__and_i_i9_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3__and_i_i9_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3__and_i_i9_1_NO_SHIFT_REG = rnode_385to386_bb3__and_i_i9_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb3__and_i_i9_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb3__and_i_i9_2_NO_SHIFT_REG = rnode_385to386_bb3__and_i_i9_0_reg_386_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_shl65_i54_stall_local;
wire [31:0] local_bb3_shl65_i54;

assign local_bb3_shl65_i54 = ((local_bb3_or64_i53 & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot30_i38_stall_local;
wire local_bb3_lnot30_i38;

assign local_bb3_lnot30_i38 = ((rnode_388to389_bb3_and20_i28_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i50_stall_local;
wire [31:0] local_bb3_or_i50;

assign local_bb3_or_i50 = ((rnode_388to389_bb3_and20_i28_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_389to391_bb3_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb3_and35_i34_0_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and35_i34_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb3_and35_i34_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and35_i34_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and35_i34_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and35_i34_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_389to391_bb3_and35_i34_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to391_bb3_and35_i34_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to391_bb3_and35_i34_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_389to391_bb3_and35_i34_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_389to391_bb3_and35_i34_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((rnode_388to389_bb3_and35_i34_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_389to391_bb3_and35_i34_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_389to391_bb3_and35_i34_0_reg_391_fifo.DEPTH = 2;
defparam rnode_389to391_bb3_and35_i34_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_389to391_bb3_and35_i34_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to391_bb3_and35_i34_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_389to391_bb3_and35_i34_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_and35_i34_0_NO_SHIFT_REG = rnode_389to391_bb3_and35_i34_0_reg_391_NO_SHIFT_REG;
assign rnode_389to391_bb3_and35_i34_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_not_i37_stall_local;
wire local_bb3_cmp25_not_i37;

assign local_bb3_cmp25_not_i37 = (local_bb3_cmp25_i32 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u82_stall_local;
wire local_bb3_var__u82;

assign local_bb3_var__u82 = (local_bb3_cmp25_i32 | rnode_387to389_bb3_cmp27_i33_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_and9_i_i_stall_local;
wire [31:0] local_bb3_and9_i_i;

assign local_bb3_and9_i_i = ((rnode_385to386_bb3__and_i_i9_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_and203_i_stall_local;
wire [31:0] local_bb3_and203_i;

assign local_bb3_and203_i = ((rnode_385to386_bb3__and_i_i9_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_and206_i_stall_local;
wire [31:0] local_bb3_and206_i;

assign local_bb3_and206_i = ((rnode_385to386_bb3__and_i_i9_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb3__28_i55_stall_local;
wire [31:0] local_bb3__28_i55;

assign local_bb3__28_i55 = (rnode_387to388_bb3_lnot23_i31_0_NO_SHIFT_REG ? 32'h0 : ((local_bb3_shl65_i54 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot30_not_i42_stall_local;
wire local_bb3_lnot30_not_i42;

assign local_bb3_lnot30_not_i42 = (local_bb3_lnot30_i38 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i51_stall_local;
wire [31:0] local_bb3_shl_i51;

assign local_bb3_shl_i51 = ((local_bb3_or_i50 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb3_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3_and35_i34_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and35_i34_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3_and35_i34_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and35_i34_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and35_i34_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and35_i34_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb3_and35_i34_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb3_and35_i34_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb3_and35_i34_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb3_and35_i34_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb3_and35_i34_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((rnode_389to391_bb3_and35_i34_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_391to392_bb3_and35_i34_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb3_and35_i34_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb3_and35_i34_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb3_and35_i34_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb3_and35_i34_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb3_and35_i34_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to391_bb3_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_and35_i34_0_NO_SHIFT_REG = rnode_391to392_bb3_and35_i34_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb3_and35_i34_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_or_cond_i39_stall_local;
wire local_bb3_or_cond_i39;

assign local_bb3_or_cond_i39 = (local_bb3_lnot30_i38 | local_bb3_cmp25_not_i37);

// This section implements an unregistered operation.
// 
wire local_bb3_sub239_i_stall_local;
wire [31:0] local_bb3_sub239_i;

assign local_bb3_sub239_i = (32'h0 - (local_bb3_and9_i_i & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb3_shl204_i_stall_local;
wire [31:0] local_bb3_shl204_i;

assign local_bb3_shl204_i = ((rnode_385to386_bb3_and193_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb3_and203_i & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb3_and72_i60_stall_local;
wire [31:0] local_bb3_and72_i60;

assign local_bb3_and72_i60 = ((local_bb3__28_i55 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb3_and75_i63_stall_local;
wire [31:0] local_bb3_and75_i63;

assign local_bb3_and75_i63 = ((local_bb3__28_i55 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb3_and78_i65_stall_local;
wire [31:0] local_bb3_and78_i65;

assign local_bb3_and78_i65 = ((local_bb3__28_i55 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb3_shr94_i68_stall_local;
wire [31:0] local_bb3_shr94_i68;

assign local_bb3_shr94_i68 = ((local_bb3__28_i55 & 32'h7FFFFF8) >> (local_bb3_and93_i67 & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb3_and90_i71_stall_local;
wire [31:0] local_bb3_and90_i71;

assign local_bb3_and90_i71 = ((local_bb3__28_i55 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb3_and87_i72_stall_local;
wire [31:0] local_bb3_and87_i72;

assign local_bb3_and87_i72 = ((local_bb3__28_i55 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb3_and84_i73_stall_local;
wire [31:0] local_bb3_and84_i73;

assign local_bb3_and84_i73 = ((local_bb3__28_i55 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u83_stall_local;
wire [31:0] local_bb3_var__u83;

assign local_bb3_var__u83 = ((local_bb3__28_i55 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb3_or_cond_not_i43_stall_local;
wire local_bb3_or_cond_not_i43;

assign local_bb3_or_cond_not_i43 = (local_bb3_cmp25_i32 & local_bb3_lnot30_not_i42);

// This section implements an unregistered operation.
// 
wire local_bb3__27_i52_stall_local;
wire [31:0] local_bb3__27_i52;

assign local_bb3__27_i52 = (local_bb3_lnot_i30 ? 32'h0 : ((local_bb3_shl_i51 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_8_i47_stall_local;
wire local_bb3_reduction_8_i47;

assign local_bb3_reduction_8_i47 = (rnode_387to389_bb3_cmp27_i33_1_NO_SHIFT_REG & local_bb3_or_cond_i39);

// This section implements an unregistered operation.
// 
wire local_bb3_cond244_i_stall_local;
wire [31:0] local_bb3_cond244_i;

assign local_bb3_cond244_i = (rnode_384to386_bb3_cmp37_i_2_NO_SHIFT_REG ? local_bb3_sub239_i : (local_bb3__43_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and205_i_stall_local;
wire [31:0] local_bb3_and205_i;

assign local_bb3_and205_i = (local_bb3_shl204_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and72_tr_i61_stall_local;
wire [7:0] local_bb3_and72_tr_i61;
wire [31:0] local_bb3_and72_tr_i61$ps;

assign local_bb3_and72_tr_i61$ps = (local_bb3_and72_i60 & 32'hFFFFFF);
assign local_bb3_and72_tr_i61 = local_bb3_and72_tr_i61$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb3_cmp76_i64_stall_local;
wire local_bb3_cmp76_i64;

assign local_bb3_cmp76_i64 = ((local_bb3_and75_i63 & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp79_i66_stall_local;
wire local_bb3_cmp79_i66;

assign local_bb3_cmp79_i66 = ((local_bb3_and78_i65 & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and142_i95_stall_local;
wire [31:0] local_bb3_and142_i95;

assign local_bb3_and142_i95 = (local_bb3_shr94_i68 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_shr150_i97_stall_local;
wire [31:0] local_bb3_shr150_i97;

assign local_bb3_shr150_i97 = (local_bb3_shr94_i68 >> (local_bb3_and149_i96 & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u84_stall_local;
wire [31:0] local_bb3_var__u84;

assign local_bb3_var__u84 = (local_bb3_shr94_i68 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and146_i100_stall_local;
wire [31:0] local_bb3_and146_i100;

assign local_bb3_and146_i100 = (local_bb3_shr94_i68 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp91_i74_stall_local;
wire local_bb3_cmp91_i74;

assign local_bb3_cmp91_i74 = ((local_bb3_and90_i71 & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp88_i75_stall_local;
wire local_bb3_cmp88_i75;

assign local_bb3_cmp88_i75 = ((local_bb3_and87_i72 & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp85_i76_stall_local;
wire local_bb3_cmp85_i76;

assign local_bb3_cmp85_i76 = ((local_bb3_and84_i73 & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u85_stall_local;
wire local_bb3_var__u85;

assign local_bb3_var__u85 = ((local_bb3_var__u83 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_add245_i_stall_local;
wire [31:0] local_bb3_add245_i;

assign local_bb3_add245_i = (local_bb3_cond244_i + (rnode_384to386_bb3_and17_i_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_fold_i10_stall_local;
wire [31:0] local_bb3_fold_i10;

assign local_bb3_fold_i10 = (local_bb3_cond244_i + (rnode_384to386_bb3_shr16_i_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb3_shl207_i_stall_local;
wire [31:0] local_bb3_shl207_i;

assign local_bb3_shl207_i = ((local_bb3_and205_i & 32'h7FFFFFF) << (local_bb3_and206_i & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb3_frombool74_i62_stall_local;
wire [7:0] local_bb3_frombool74_i62;

assign local_bb3_frombool74_i62 = (local_bb3_and72_tr_i61 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u86_stall_local;
wire [31:0] local_bb3_var__u86;

assign local_bb3_var__u86 = ((local_bb3_and146_i100 & 32'h3FFFFFFF) | local_bb3_shr94_i68);

// This section implements an unregistered operation.
// 
wire local_bb3__31_v_i82_stall_local;
wire local_bb3__31_v_i82;

assign local_bb3__31_v_i82 = (local_bb3_cmp96_i70 ? local_bb3_cmp79_i66 : local_bb3_cmp91_i74);

// This section implements an unregistered operation.
// 
wire local_bb3__30_v_i80_stall_local;
wire local_bb3__30_v_i80;

assign local_bb3__30_v_i80 = (local_bb3_cmp96_i70 ? local_bb3_cmp76_i64 : local_bb3_cmp88_i75);

// This section implements an unregistered operation.
// 
wire local_bb3_frombool109_i78_stall_local;
wire [7:0] local_bb3_frombool109_i78;

assign local_bb3_frombool109_i78[7:1] = 7'h0;
assign local_bb3_frombool109_i78[0] = local_bb3_cmp85_i76;

// This section implements an unregistered operation.
// 
wire local_bb3_or107_i77_stall_local;
wire [31:0] local_bb3_or107_i77;

assign local_bb3_or107_i77[31:1] = 31'h0;
assign local_bb3_or107_i77[0] = local_bb3_var__u85;

// This section implements an unregistered operation.
// 
wire local_bb3_and250_i_stall_local;
wire [31:0] local_bb3_and250_i;

assign local_bb3_and250_i = (local_bb3_fold_i10 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and269_i_stall_local;
wire [31:0] local_bb3_and269_i;

assign local_bb3_and269_i = (local_bb3_fold_i10 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and208_i_stall_local;
wire [31:0] local_bb3_and208_i;

assign local_bb3_and208_i = (local_bb3_shl207_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_or1596_i101_stall_local;
wire [31:0] local_bb3_or1596_i101;

assign local_bb3_or1596_i101 = (local_bb3_var__u86 | (local_bb3_and142_i95 & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3__31_i83_stall_local;
wire [7:0] local_bb3__31_i83;

assign local_bb3__31_i83[7:1] = 7'h0;
assign local_bb3__31_i83[0] = local_bb3__31_v_i82;

// This section implements an unregistered operation.
// 
wire local_bb3__30_i81_stall_local;
wire [7:0] local_bb3__30_i81;

assign local_bb3__30_i81[7:1] = 7'h0;
assign local_bb3__30_i81[0] = local_bb3__30_v_i80;

// This section implements an unregistered operation.
// 
wire local_bb3__29_i79_stall_local;
wire [7:0] local_bb3__29_i79;

assign local_bb3__29_i79 = (local_bb3_cmp96_i70 ? (local_bb3_frombool74_i62 & 8'h1) : (local_bb3_frombool109_i78 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__32_i84_stall_local;
wire [31:0] local_bb3__32_i84;

assign local_bb3__32_i84 = (local_bb3_cmp96_i70 ? 32'h0 : (local_bb3_or107_i77 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__44_i_stall_local;
wire [31:0] local_bb3__44_i;

assign local_bb3__44_i = (local_bb3__40_demorgan_i ? (local_bb3_and208_i & 32'h7FFFFFF) : (local_bb3_or219_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_or162_i102_stall_local;
wire [31:0] local_bb3_or162_i102;

assign local_bb3_or162_i102 = (local_bb3_or1596_i101 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or1237_i87_stall_local;
wire [7:0] local_bb3_or1237_i87;

assign local_bb3_or1237_i87 = ((local_bb3__30_i81 & 8'h1) | (local_bb3__29_i79 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3__33_i89_stall_local;
wire [7:0] local_bb3__33_i89;

assign local_bb3__33_i89 = (local_bb3_cmp116_i86 ? (local_bb3__29_i79 & 8'h1) : (local_bb3__31_i83 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and250_i_valid_out;
wire local_bb3_and250_i_stall_in;
wire local_bb3_and269_i_valid_out;
wire local_bb3_and269_i_stall_in;
wire local_bb3_add245_i_valid_out;
wire local_bb3_add245_i_stall_in;
wire local_bb3__45_i_valid_out;
wire local_bb3__45_i_stall_in;
wire local_bb3_not_cmp37_i_valid_out_1;
wire local_bb3_not_cmp37_i_stall_in_1;
wire local_bb3__45_i_inputs_ready;
wire local_bb3__45_i_stall_local;
wire [31:0] local_bb3__45_i;

assign local_bb3__45_i_inputs_ready = (rnode_384to386_bb3_shr16_i_0_valid_out_NO_SHIFT_REG & rnode_384to386_bb3_and17_i_0_valid_out_NO_SHIFT_REG & rnode_384to386_bb3_cmp37_i_0_valid_out_2_NO_SHIFT_REG & rnode_384to386_bb3_cmp37_i_0_valid_out_0_NO_SHIFT_REG & rnode_385to386_bb3_and193_i_0_valid_out_2_NO_SHIFT_REG & rnode_384to386_bb3_cmp37_i_0_valid_out_1_NO_SHIFT_REG & rnode_385to386_bb3_and195_i_0_valid_out_NO_SHIFT_REG & rnode_385to386_bb3_and193_i_0_valid_out_1_NO_SHIFT_REG & rnode_385to386_bb3_and198_i_0_valid_out_NO_SHIFT_REG & rnode_385to386_bb3_and193_i_0_valid_out_0_NO_SHIFT_REG & rnode_385to386_bb3__and_i_i9_0_valid_out_1_NO_SHIFT_REG & rnode_385to386_bb3__and_i_i9_0_valid_out_2_NO_SHIFT_REG & rnode_385to386_bb3__and_i_i9_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3__45_i = (local_bb3__42_i ? (rnode_385to386_bb3_and193_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb3__44_i & 32'h7FFFFFF));
assign local_bb3_and250_i_valid_out = 1'b1;
assign local_bb3_and269_i_valid_out = 1'b1;
assign local_bb3_add245_i_valid_out = 1'b1;
assign local_bb3__45_i_valid_out = 1'b1;
assign local_bb3_not_cmp37_i_valid_out_1 = 1'b1;
assign rnode_384to386_bb3_shr16_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_and17_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_cmp37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb3_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and195_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and198_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3_and193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3__and_i_i9_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3__and_i_i9_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb3__and_i_i9_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__37_v_i103_stall_local;
wire [31:0] local_bb3__37_v_i103;

assign local_bb3__37_v_i103 = (local_bb3_Pivot20_i98 ? 32'h0 : (local_bb3_or162_i102 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or123_i88_stall_local;
wire [31:0] local_bb3_or123_i88;

assign local_bb3_or123_i88[31:8] = 24'h0;
assign local_bb3_or123_i88[7:0] = (local_bb3_or1237_i87 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u87_stall_local;
wire [7:0] local_bb3_var__u87;

assign local_bb3_var__u87 = ((local_bb3__33_i89 & 8'h1) & 8'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_and250_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and250_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_and250_i_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and250_i_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_and250_i_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and250_i_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and250_i_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_and250_i_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_and250_i_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_and250_i_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_and250_i_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_and250_i_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_and250_i_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in((local_bb3_and250_i & 32'hFF)),
	.data_out(rnode_386to387_bb3_and250_i_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_and250_i_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_and250_i_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb3_and250_i_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_and250_i_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_and250_i_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and250_i_stall_in = 1'b0;
assign rnode_386to387_bb3_and250_i_0_NO_SHIFT_REG = rnode_386to387_bb3_and250_i_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_and250_i_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_and250_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_386to388_bb3_and269_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to388_bb3_and269_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_386to388_bb3_and269_i_0_NO_SHIFT_REG;
 logic rnode_386to388_bb3_and269_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to388_bb3_and269_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_386to388_bb3_and269_i_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_386to388_bb3_and269_i_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_386to388_bb3_and269_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_386to388_bb3_and269_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to388_bb3_and269_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to388_bb3_and269_i_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_386to388_bb3_and269_i_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_386to388_bb3_and269_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in((local_bb3_and269_i & 32'hFF800000)),
	.data_out(rnode_386to388_bb3_and269_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_386to388_bb3_and269_i_0_reg_388_fifo.DEPTH = 2;
defparam rnode_386to388_bb3_and269_i_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_386to388_bb3_and269_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to388_bb3_and269_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_386to388_bb3_and269_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and269_i_stall_in = 1'b0;
assign rnode_386to388_bb3_and269_i_0_NO_SHIFT_REG = rnode_386to388_bb3_and269_i_0_reg_388_NO_SHIFT_REG;
assign rnode_386to388_bb3_and269_i_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_386to388_bb3_and269_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_add245_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_add245_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_add245_i_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_add245_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3_add245_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_add245_i_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3_add245_i_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3_add245_i_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_add245_i_0_valid_out_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_add245_i_0_stall_in_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_add245_i_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_add245_i_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_add245_i_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_add245_i_0_stall_in_0_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_add245_i_0_valid_out_0_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_add245_i_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(local_bb3_add245_i),
	.data_out(rnode_386to387_bb3_add245_i_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_add245_i_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_add245_i_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb3_add245_i_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_add245_i_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_add245_i_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add245_i_stall_in = 1'b0;
assign rnode_386to387_bb3_add245_i_0_stall_in_0_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_add245_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3_add245_i_0_NO_SHIFT_REG = rnode_386to387_bb3_add245_i_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_add245_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3_add245_i_1_NO_SHIFT_REG = rnode_386to387_bb3_add245_i_0_reg_387_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3__45_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3__45_i_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3__45_i_1_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3__45_i_2_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb3__45_i_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_valid_out_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_stall_in_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3__45_i_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3__45_i_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3__45_i_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3__45_i_0_stall_in_0_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3__45_i_0_valid_out_0_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3__45_i_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in((local_bb3__45_i & 32'hFFFFFFF)),
	.data_out(rnode_386to387_bb3__45_i_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3__45_i_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3__45_i_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb3__45_i_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3__45_i_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3__45_i_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__45_i_stall_in = 1'b0;
assign rnode_386to387_bb3__45_i_0_stall_in_0_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3__45_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3__45_i_0_NO_SHIFT_REG = rnode_386to387_bb3__45_i_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3__45_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3__45_i_1_NO_SHIFT_REG = rnode_386to387_bb3__45_i_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3__45_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb3__45_i_2_NO_SHIFT_REG = rnode_386to387_bb3__45_i_0_reg_387_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb3_not_cmp37_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to387_bb3_not_cmp37_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_386to387_bb3_not_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_386to387_bb3_not_cmp37_i_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_386to387_bb3_not_cmp37_i_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_not_cmp37_i_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_not_cmp37_i_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb3_not_cmp37_i_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb3_not_cmp37_i_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb3_not_cmp37_i_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb3_not_cmp37_i_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb3_not_cmp37_i_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb3_not_cmp37_i_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(local_bb3_not_cmp37_i),
	.data_out(rnode_386to387_bb3_not_cmp37_i_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb3_not_cmp37_i_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb3_not_cmp37_i_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_386to387_bb3_not_cmp37_i_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb3_not_cmp37_i_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb3_not_cmp37_i_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_not_cmp37_i_stall_in_1 = 1'b0;
assign rnode_386to387_bb3_not_cmp37_i_0_NO_SHIFT_REG = rnode_386to387_bb3_not_cmp37_i_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb3_not_cmp37_i_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_not_cmp37_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__39_v_i104_stall_local;
wire [31:0] local_bb3__39_v_i104;

assign local_bb3__39_v_i104 = (local_bb3_SwitchLeaf_i99 ? (local_bb3_var__u84 & 32'h1) : (local_bb3__37_v_i103 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or124_i90_stall_local;
wire [31:0] local_bb3_or124_i90;

assign local_bb3_or124_i90 = (local_bb3_cmp116_i86 ? 32'h0 : (local_bb3_or123_i88 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_conv135_i92_stall_local;
wire [31:0] local_bb3_conv135_i92;

assign local_bb3_conv135_i92[31:8] = 24'h0;
assign local_bb3_conv135_i92[7:0] = (local_bb3_var__u87 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_notrhs_i_stall_local;
wire local_bb3_notrhs_i;

assign local_bb3_notrhs_i = ((rnode_386to387_bb3_and250_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_shl273_i_stall_local;
wire [31:0] local_bb3_shl273_i;

assign local_bb3_shl273_i = ((rnode_386to388_bb3_and269_i_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb3_and247_i_stall_local;
wire [31:0] local_bb3_and247_i;

assign local_bb3_and247_i = (rnode_386to387_bb3_add245_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp258_i_stall_local;
wire local_bb3_cmp258_i;

assign local_bb3_cmp258_i = ($signed(rnode_386to387_bb3_add245_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb3_and225_i_stall_local;
wire [31:0] local_bb3_and225_i;

assign local_bb3_and225_i = ((rnode_386to387_bb3__45_i_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and270_i_stall_local;
wire [31:0] local_bb3_and270_i;

assign local_bb3_and270_i = ((rnode_386to387_bb3__45_i_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb3_shr271_i_valid_out;
wire local_bb3_shr271_i_stall_in;
wire local_bb3_shr271_i_inputs_ready;
wire local_bb3_shr271_i_stall_local;
wire [31:0] local_bb3_shr271_i;

assign local_bb3_shr271_i_inputs_ready = rnode_386to387_bb3__45_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_shr271_i = ((rnode_386to387_bb3__45_i_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb3_shr271_i_valid_out = 1'b1;
assign rnode_386to387_bb3__45_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_3_i105_stall_local;
wire [31:0] local_bb3_reduction_3_i105;

assign local_bb3_reduction_3_i105 = ((local_bb3__32_i84 & 32'h1) | (local_bb3_or124_i90 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or136_i94_stall_local;
wire [31:0] local_bb3_or136_i94;

assign local_bb3_or136_i94 = (local_bb3_cmp131_not_i93 ? (local_bb3_conv135_i92 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_notlhs_i_stall_local;
wire local_bb3_notlhs_i;

assign local_bb3_notlhs_i = ((local_bb3_and247_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp226_i_stall_local;
wire local_bb3_cmp226_i;

assign local_bb3_cmp226_i = ((local_bb3_and225_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp296_i_stall_local;
wire local_bb3_cmp296_i;

assign local_bb3_cmp296_i = ((local_bb3_and270_i & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp296_i_valid_out;
wire local_bb3_cmp296_i_stall_in;
wire local_bb3_cmp299_i_valid_out;
wire local_bb3_cmp299_i_stall_in;
wire local_bb3_cmp299_i_inputs_ready;
wire local_bb3_cmp299_i_stall_local;
wire local_bb3_cmp299_i;

assign local_bb3_cmp299_i_inputs_ready = rnode_386to387_bb3__45_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_cmp299_i = ((local_bb3_and270_i & 32'h7) == 32'h4);
assign local_bb3_cmp296_i_valid_out = 1'b1;
assign local_bb3_cmp299_i_valid_out = 1'b1;
assign rnode_386to387_bb3__45_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_shr271_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb3_shr271_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_shr271_i_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_shr271_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_shr271_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_shr271_i_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_shr271_i_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_shr271_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_shr271_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_shr271_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_shr271_i_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_shr271_i_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_shr271_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in((local_bb3_shr271_i & 32'h1FFFFFF)),
	.data_out(rnode_387to388_bb3_shr271_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_shr271_i_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_shr271_i_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb3_shr271_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_shr271_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_shr271_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr271_i_stall_in = 1'b0;
assign rnode_387to388_bb3_shr271_i_0_NO_SHIFT_REG = rnode_387to388_bb3_shr271_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_shr271_i_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_shr271_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_5_i107_stall_local;
wire [31:0] local_bb3_reduction_5_i107;

assign local_bb3_reduction_5_i107 = (local_bb3_shr150_i97 | (local_bb3_reduction_3_i105 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_4_i106_stall_local;
wire [31:0] local_bb3_reduction_4_i106;

assign local_bb3_reduction_4_i106 = ((local_bb3_or136_i94 & 32'h1) | (local_bb3__39_v_i104 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_not__46_i_stall_local;
wire local_bb3_not__46_i;

assign local_bb3_not__46_i = (local_bb3_notrhs_i | local_bb3_notlhs_i);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp226_not_i_stall_local;
wire local_bb3_cmp226_not_i;

assign local_bb3_cmp226_not_i = (local_bb3_cmp226_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_cmp296_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp296_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp296_i_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp296_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp296_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp296_i_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp296_i_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp296_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_cmp296_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_cmp296_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_cmp296_i_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_cmp296_i_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_cmp296_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb3_cmp296_i),
	.data_out(rnode_387to388_bb3_cmp296_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_cmp296_i_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_cmp296_i_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb3_cmp296_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_cmp296_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_cmp296_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp296_i_stall_in = 1'b0;
assign rnode_387to388_bb3_cmp296_i_0_NO_SHIFT_REG = rnode_387to388_bb3_cmp296_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_cmp296_i_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_cmp296_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_cmp299_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp299_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp299_i_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp299_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp299_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp299_i_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp299_i_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_cmp299_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_cmp299_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_cmp299_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_cmp299_i_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_cmp299_i_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_cmp299_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb3_cmp299_i),
	.data_out(rnode_387to388_bb3_cmp299_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_cmp299_i_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_cmp299_i_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb3_cmp299_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_cmp299_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_cmp299_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp299_i_stall_in = 1'b0;
assign rnode_387to388_bb3_cmp299_i_0_NO_SHIFT_REG = rnode_387to388_bb3_cmp299_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_cmp299_i_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_cmp299_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and272_i_stall_local;
wire [31:0] local_bb3_and272_i;

assign local_bb3_and272_i = ((rnode_387to388_bb3_shr271_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_6_i108_stall_local;
wire [31:0] local_bb3_reduction_6_i108;

assign local_bb3_reduction_6_i108 = ((local_bb3_reduction_4_i106 & 32'h1) | local_bb3_reduction_5_i107);

// This section implements an unregistered operation.
// 
wire local_bb3__47_i_stall_local;
wire local_bb3__47_i;

assign local_bb3__47_i = (local_bb3_cmp226_i | local_bb3_not__46_i);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge12_i_stall_local;
wire local_bb3_brmerge12_i;

assign local_bb3_brmerge12_i = (local_bb3_cmp226_not_i | rnode_386to387_bb3_not_cmp37_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot262__i_stall_local;
wire local_bb3_lnot262__i;

assign local_bb3_lnot262__i = (local_bb3_cmp258_i & local_bb3_cmp226_not_i);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp29649_i_stall_local;
wire [31:0] local_bb3_cmp29649_i;

assign local_bb3_cmp29649_i[31:1] = 31'h0;
assign local_bb3_cmp29649_i[0] = rnode_387to388_bb3_cmp296_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_conv300_i_stall_local;
wire [31:0] local_bb3_conv300_i;

assign local_bb3_conv300_i[31:1] = 31'h0;
assign local_bb3_conv300_i[0] = rnode_387to388_bb3_cmp299_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or274_i_stall_local;
wire [31:0] local_bb3_or274_i;

assign local_bb3_or274_i = ((local_bb3_and272_i & 32'h7FFFFF) | (local_bb3_shl273_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb3_lnot33_not_i40_valid_out;
wire local_bb3_lnot33_not_i40_stall_in;
wire local_bb3_cmp37_i36_valid_out;
wire local_bb3_cmp37_i36_stall_in;
wire local_bb3_and36_lobit_i111_valid_out;
wire local_bb3_and36_lobit_i111_stall_in;
wire local_bb3_xor188_i110_valid_out;
wire local_bb3_xor188_i110_stall_in;
wire local_bb3_xor188_i110_inputs_ready;
wire local_bb3_xor188_i110_stall_local;
wire [31:0] local_bb3_xor188_i110;

assign local_bb3_xor188_i110_inputs_ready = (rnode_387to388_bb3__22_i22_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb3_lnot23_i31_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb3_align_0_i59_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb3_align_0_i59_0_valid_out_4_NO_SHIFT_REG & rnode_387to388_bb3_align_0_i59_0_valid_out_1_NO_SHIFT_REG & rnode_387to388_bb3_align_0_i59_0_valid_out_2_NO_SHIFT_REG & rnode_387to388_bb3_align_0_i59_0_valid_out_3_NO_SHIFT_REG & rnode_387to388_bb3__23_i23_0_valid_out_2_NO_SHIFT_REG & rnode_387to388_bb3__22_i22_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_xor188_i110 = (local_bb3_reduction_6_i108 ^ local_bb3_xor_lobit_i109);
assign local_bb3_lnot33_not_i40_valid_out = 1'b1;
assign local_bb3_cmp37_i36_valid_out = 1'b1;
assign local_bb3_and36_lobit_i111_valid_out = 1'b1;
assign local_bb3_xor188_i110_valid_out = 1'b1;
assign rnode_387to388_bb3__22_i22_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_lnot23_i31_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_align_0_i59_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_align_0_i59_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_align_0_i59_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_align_0_i59_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_align_0_i59_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__23_i23_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__22_i22_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_resultSign_0_i_stall_local;
wire [31:0] local_bb3_resultSign_0_i;

assign local_bb3_resultSign_0_i = (local_bb3_brmerge12_i ? (rnode_386to387_bb3_and35_i_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_resultSign_0_i_valid_out;
wire local_bb3_resultSign_0_i_stall_in;
wire local_bb3__47_i_valid_out;
wire local_bb3__47_i_stall_in;
wire local_bb3_or2662_i_valid_out;
wire local_bb3_or2662_i_stall_in;
wire local_bb3_or2662_i_inputs_ready;
wire local_bb3_or2662_i_stall_local;
wire local_bb3_or2662_i;

assign local_bb3_or2662_i_inputs_ready = (rnode_386to387_bb3_and35_i_0_valid_out_NO_SHIFT_REG & rnode_386to387_bb3_not_cmp37_i_0_valid_out_NO_SHIFT_REG & rnode_386to387_bb3_add245_i_0_valid_out_0_NO_SHIFT_REG & rnode_386to387_bb3_and250_i_0_valid_out_NO_SHIFT_REG & rnode_386to387_bb3__45_i_0_valid_out_0_NO_SHIFT_REG & rnode_386to387_bb3_add245_i_0_valid_out_1_NO_SHIFT_REG & rnode_386to387_bb3_var__u72_0_valid_out_NO_SHIFT_REG);
assign local_bb3_or2662_i = (rnode_386to387_bb3_var__u72_0_NO_SHIFT_REG | local_bb3_lnot262__i);
assign local_bb3_resultSign_0_i_valid_out = 1'b1;
assign local_bb3__47_i_valid_out = 1'b1;
assign local_bb3_or2662_i_valid_out = 1'b1;
assign rnode_386to387_bb3_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_not_cmp37_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_add245_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_and250_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3__45_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_add245_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb3_var__u72_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3_lnot33_not_i40_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb3_lnot33_not_i40_0_stall_in_NO_SHIFT_REG;
 logic rnode_388to389_bb3_lnot33_not_i40_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_lnot33_not_i40_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic rnode_388to389_bb3_lnot33_not_i40_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_lnot33_not_i40_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_lnot33_not_i40_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_lnot33_not_i40_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3_lnot33_not_i40_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3_lnot33_not_i40_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3_lnot33_not_i40_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3_lnot33_not_i40_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3_lnot33_not_i40_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb3_lnot33_not_i40),
	.data_out(rnode_388to389_bb3_lnot33_not_i40_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3_lnot33_not_i40_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3_lnot33_not_i40_0_reg_389_fifo.DATA_WIDTH = 1;
defparam rnode_388to389_bb3_lnot33_not_i40_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3_lnot33_not_i40_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3_lnot33_not_i40_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_lnot33_not_i40_stall_in = 1'b0;
assign rnode_388to389_bb3_lnot33_not_i40_0_NO_SHIFT_REG = rnode_388to389_bb3_lnot33_not_i40_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3_lnot33_not_i40_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_lnot33_not_i40_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3_cmp37_i36_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_1_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_valid_out_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_stall_in_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_cmp37_i36_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3_cmp37_i36_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3_cmp37_i36_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3_cmp37_i36_0_stall_in_0_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3_cmp37_i36_0_valid_out_0_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3_cmp37_i36_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb3_cmp37_i36),
	.data_out(rnode_388to389_bb3_cmp37_i36_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3_cmp37_i36_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3_cmp37_i36_0_reg_389_fifo.DATA_WIDTH = 1;
defparam rnode_388to389_bb3_cmp37_i36_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3_cmp37_i36_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3_cmp37_i36_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp37_i36_stall_in = 1'b0;
assign rnode_388to389_bb3_cmp37_i36_0_stall_in_0_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_cmp37_i36_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3_cmp37_i36_0_NO_SHIFT_REG = rnode_388to389_bb3_cmp37_i36_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3_cmp37_i36_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3_cmp37_i36_1_NO_SHIFT_REG = rnode_388to389_bb3_cmp37_i36_0_reg_389_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3_and36_lobit_i111_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and36_lobit_i111_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_and36_lobit_i111_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and36_lobit_i111_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_and36_lobit_i111_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and36_lobit_i111_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and36_lobit_i111_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_and36_lobit_i111_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3_and36_lobit_i111_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3_and36_lobit_i111_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3_and36_lobit_i111_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3_and36_lobit_i111_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3_and36_lobit_i111_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb3_and36_lobit_i111 & 32'h1)),
	.data_out(rnode_388to389_bb3_and36_lobit_i111_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3_and36_lobit_i111_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3_and36_lobit_i111_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb3_and36_lobit_i111_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3_and36_lobit_i111_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3_and36_lobit_i111_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and36_lobit_i111_stall_in = 1'b0;
assign rnode_388to389_bb3_and36_lobit_i111_0_NO_SHIFT_REG = rnode_388to389_bb3_and36_lobit_i111_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3_and36_lobit_i111_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_and36_lobit_i111_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3_xor188_i110_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb3_xor188_i110_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_xor188_i110_0_NO_SHIFT_REG;
 logic rnode_388to389_bb3_xor188_i110_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3_xor188_i110_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_xor188_i110_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_xor188_i110_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3_xor188_i110_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3_xor188_i110_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3_xor188_i110_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3_xor188_i110_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3_xor188_i110_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3_xor188_i110_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb3_xor188_i110),
	.data_out(rnode_388to389_bb3_xor188_i110_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3_xor188_i110_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3_xor188_i110_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb3_xor188_i110_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3_xor188_i110_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3_xor188_i110_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_xor188_i110_stall_in = 1'b0;
assign rnode_388to389_bb3_xor188_i110_0_NO_SHIFT_REG = rnode_388to389_bb3_xor188_i110_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3_xor188_i110_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_xor188_i110_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_resultSign_0_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb3_resultSign_0_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_resultSign_0_i_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_resultSign_0_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb3_resultSign_0_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_resultSign_0_i_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_resultSign_0_i_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_resultSign_0_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_resultSign_0_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_resultSign_0_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_resultSign_0_i_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_resultSign_0_i_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_resultSign_0_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in((local_bb3_resultSign_0_i & 32'h80000000)),
	.data_out(rnode_387to388_bb3_resultSign_0_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_resultSign_0_i_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_resultSign_0_i_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb3_resultSign_0_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_resultSign_0_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_resultSign_0_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_resultSign_0_i_stall_in = 1'b0;
assign rnode_387to388_bb3_resultSign_0_i_0_NO_SHIFT_REG = rnode_387to388_bb3_resultSign_0_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_resultSign_0_i_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_resultSign_0_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3__47_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3__47_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3__47_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3__47_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3__47_i_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3__47_i_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3__47_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb3__47_i),
	.data_out(rnode_387to388_bb3__47_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3__47_i_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3__47_i_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb3__47_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3__47_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3__47_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__47_i_stall_in = 1'b0;
assign rnode_387to388_bb3__47_i_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__47_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__47_i_0_NO_SHIFT_REG = rnode_387to388_bb3__47_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3__47_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3__47_i_1_NO_SHIFT_REG = rnode_387to388_bb3__47_i_0_reg_388_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb3_or2662_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_1_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_2_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb3_or2662_i_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb3_or2662_i_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb3_or2662_i_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb3_or2662_i_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb3_or2662_i_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb3_or2662_i_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb3_or2662_i),
	.data_out(rnode_387to388_bb3_or2662_i_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb3_or2662_i_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb3_or2662_i_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb3_or2662_i_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb3_or2662_i_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb3_or2662_i_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or2662_i_stall_in = 1'b0;
assign rnode_387to388_bb3_or2662_i_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_or2662_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_or2662_i_0_NO_SHIFT_REG = rnode_387to388_bb3_or2662_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_or2662_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_or2662_i_1_NO_SHIFT_REG = rnode_387to388_bb3_or2662_i_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb3_or2662_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb3_or2662_i_2_NO_SHIFT_REG = rnode_387to388_bb3_or2662_i_0_reg_388_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge_not_i41_stall_local;
wire local_bb3_brmerge_not_i41;

assign local_bb3_brmerge_not_i41 = (rnode_387to389_bb3_cmp27_i33_0_NO_SHIFT_REG & rnode_388to389_bb3_lnot33_not_i40_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_389to391_bb3_cmp37_i36_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_1_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_2_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_valid_out_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_stall_in_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_cmp37_i36_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_389to391_bb3_cmp37_i36_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to391_bb3_cmp37_i36_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to391_bb3_cmp37_i36_0_stall_in_0_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_389to391_bb3_cmp37_i36_0_valid_out_0_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_389to391_bb3_cmp37_i36_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in(rnode_388to389_bb3_cmp37_i36_1_NO_SHIFT_REG),
	.data_out(rnode_389to391_bb3_cmp37_i36_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_389to391_bb3_cmp37_i36_0_reg_391_fifo.DEPTH = 2;
defparam rnode_389to391_bb3_cmp37_i36_0_reg_391_fifo.DATA_WIDTH = 1;
defparam rnode_389to391_bb3_cmp37_i36_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to391_bb3_cmp37_i36_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_389to391_bb3_cmp37_i36_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3_cmp37_i36_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_cmp37_i36_0_stall_in_0_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_cmp37_i36_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_389to391_bb3_cmp37_i36_0_NO_SHIFT_REG = rnode_389to391_bb3_cmp37_i36_0_reg_391_NO_SHIFT_REG;
assign rnode_389to391_bb3_cmp37_i36_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_389to391_bb3_cmp37_i36_1_NO_SHIFT_REG = rnode_389to391_bb3_cmp37_i36_0_reg_391_NO_SHIFT_REG;
assign rnode_389to391_bb3_cmp37_i36_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_389to391_bb3_cmp37_i36_2_NO_SHIFT_REG = rnode_389to391_bb3_cmp37_i36_0_reg_391_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_add_i112_stall_local;
wire [31:0] local_bb3_add_i112;

assign local_bb3_add_i112 = ((local_bb3__27_i52 & 32'h7FFFFF8) | (rnode_388to389_bb3_and36_lobit_i111_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_or275_i_stall_local;
wire [31:0] local_bb3_or275_i;

assign local_bb3_or275_i = ((local_bb3_or274_i & 32'h7FFFFFFF) | (rnode_387to388_bb3_resultSign_0_i_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u88_stall_local;
wire [31:0] local_bb3_var__u88;

assign local_bb3_var__u88[31:1] = 31'h0;
assign local_bb3_var__u88[0] = rnode_387to388_bb3__47_i_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or2804_i_stall_local;
wire local_bb3_or2804_i;

assign local_bb3_or2804_i = (rnode_387to388_bb3__47_i_0_NO_SHIFT_REG | rnode_387to388_bb3_or2662_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_or2875_i_stall_local;
wire local_bb3_or2875_i;

assign local_bb3_or2875_i = (rnode_387to388_bb3_or2662_i_1_NO_SHIFT_REG | rnode_387to388_bb3__26_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u89_stall_local;
wire [31:0] local_bb3_var__u89;

assign local_bb3_var__u89[31:1] = 31'h0;
assign local_bb3_var__u89[0] = rnode_387to388_bb3_or2662_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__24_i44_stall_local;
wire local_bb3__24_i44;

assign local_bb3__24_i44 = (local_bb3_or_cond_not_i43 | local_bb3_brmerge_not_i41);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge_not_not_i45_stall_local;
wire local_bb3_brmerge_not_not_i45;

assign local_bb3_brmerge_not_not_i45 = (local_bb3_brmerge_not_i41 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_not_cmp37_i142_stall_local;
wire local_bb3_not_cmp37_i142;

assign local_bb3_not_cmp37_i142 = (rnode_389to391_bb3_cmp37_i36_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_add192_i113_stall_local;
wire [31:0] local_bb3_add192_i113;

assign local_bb3_add192_i113 = ((local_bb3_add_i112 & 32'h7FFFFF9) + rnode_388to389_bb3_xor188_i110_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext314_i_stall_local;
wire [31:0] local_bb3_lnot_ext314_i;

assign local_bb3_lnot_ext314_i = ((local_bb3_var__u88 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cond282_i_stall_local;
wire [31:0] local_bb3_cond282_i;

assign local_bb3_cond282_i = (local_bb3_or2804_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cond289_i_stall_local;
wire [31:0] local_bb3_cond289_i;

assign local_bb3_cond289_i = (local_bb3_or2875_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext310_i_stall_local;
wire [31:0] local_bb3_lnot_ext310_i;

assign local_bb3_lnot_ext310_i = ((local_bb3_var__u89 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_7_i46_stall_local;
wire local_bb3_reduction_7_i46;

assign local_bb3_reduction_7_i46 = (local_bb3_cmp25_i32 & local_bb3_brmerge_not_not_i45);

// This section implements an unregistered operation.
// 
wire local_bb3_and293_i_stall_local;
wire [31:0] local_bb3_and293_i;

assign local_bb3_and293_i = ((local_bb3_cond282_i | 32'h80000000) & local_bb3_or275_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or294_i_stall_local;
wire [31:0] local_bb3_or294_i;

assign local_bb3_or294_i = ((local_bb3_cond289_i & 32'h7F800000) | (local_bb3_cond292_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_0_i_stall_local;
wire [31:0] local_bb3_reduction_0_i;

assign local_bb3_reduction_0_i = ((local_bb3_lnot_ext310_i & 32'h1) & (local_bb3_lnot_ext_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_9_i48_stall_local;
wire local_bb3_reduction_9_i48;

assign local_bb3_reduction_9_i48 = (local_bb3_reduction_7_i46 & local_bb3_reduction_8_i47);

// This section implements an unregistered operation.
// 
wire local_bb3_and302_i_stall_local;
wire [31:0] local_bb3_and302_i;

assign local_bb3_and302_i = ((local_bb3_conv300_i & 32'h1) & local_bb3_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or295_i_stall_local;
wire [31:0] local_bb3_or295_i;

assign local_bb3_or295_i = ((local_bb3_or294_i & 32'h7FC00000) | local_bb3_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb3_and17_i25_valid_out_2;
wire local_bb3_and17_i25_stall_in_2;
wire local_bb3_var__u82_valid_out;
wire local_bb3_var__u82_stall_in;
wire local_bb3_add192_i113_valid_out;
wire local_bb3_add192_i113_stall_in;
wire local_bb3__26_i49_valid_out;
wire local_bb3__26_i49_stall_in;
wire local_bb3__26_i49_inputs_ready;
wire local_bb3__26_i49_stall_local;
wire local_bb3__26_i49;

assign local_bb3__26_i49_inputs_ready = (rnode_387to389_bb3_shr16_i24_0_valid_out_0_NO_SHIFT_REG & rnode_387to389_bb3_cmp27_i33_0_valid_out_2_NO_SHIFT_REG & rnode_388to389_bb3_and36_lobit_i111_0_valid_out_NO_SHIFT_REG & rnode_388to389_bb3_xor188_i110_0_valid_out_NO_SHIFT_REG & rnode_388to389_bb3_and20_i28_0_valid_out_0_NO_SHIFT_REG & rnode_387to389_bb3_cmp27_i33_0_valid_out_0_NO_SHIFT_REG & rnode_388to389_bb3_lnot33_not_i40_0_valid_out_NO_SHIFT_REG & rnode_387to389_bb3_cmp27_i33_0_valid_out_1_NO_SHIFT_REG & rnode_388to389_bb3_and20_i28_0_valid_out_1_NO_SHIFT_REG & rnode_388to389_bb3_cmp37_i36_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3__26_i49 = (local_bb3_reduction_9_i48 ? rnode_388to389_bb3_cmp37_i36_0_NO_SHIFT_REG : local_bb3__24_i44);
assign local_bb3_and17_i25_valid_out_2 = 1'b1;
assign local_bb3_var__u82_valid_out = 1'b1;
assign local_bb3_add192_i113_valid_out = 1'b1;
assign local_bb3__26_i49_valid_out = 1'b1;
assign rnode_387to389_bb3_shr16_i24_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to389_bb3_cmp27_i33_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_and36_lobit_i111_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_xor188_i110_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_and20_i28_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to389_bb3_cmp27_i33_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_lnot33_not_i40_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to389_bb3_cmp27_i33_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_and20_i28_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3_cmp37_i36_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_lor_ext_i_stall_local;
wire [31:0] local_bb3_lor_ext_i;

assign local_bb3_lor_ext_i = ((local_bb3_cmp29649_i & 32'h1) | (local_bb3_and302_i & 32'h1));

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_389to391_bb3_and17_i25_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and17_i25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb3_and17_i25_0_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and17_i25_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb3_and17_i25_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and17_i25_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and17_i25_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb3_and17_i25_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_389to391_bb3_and17_i25_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to391_bb3_and17_i25_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to391_bb3_and17_i25_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_389to391_bb3_and17_i25_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_389to391_bb3_and17_i25_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb3_and17_i25 & 32'hFF)),
	.data_out(rnode_389to391_bb3_and17_i25_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_389to391_bb3_and17_i25_0_reg_391_fifo.DEPTH = 2;
defparam rnode_389to391_bb3_and17_i25_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_389to391_bb3_and17_i25_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to391_bb3_and17_i25_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_389to391_bb3_and17_i25_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and17_i25_stall_in_2 = 1'b0;
assign rnode_389to391_bb3_and17_i25_0_NO_SHIFT_REG = rnode_389to391_bb3_and17_i25_0_reg_391_NO_SHIFT_REG;
assign rnode_389to391_bb3_and17_i25_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_and17_i25_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb3_var__u82_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to390_bb3_var__u82_0_stall_in_NO_SHIFT_REG;
 logic rnode_389to390_bb3_var__u82_0_NO_SHIFT_REG;
 logic rnode_389to390_bb3_var__u82_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to390_bb3_var__u82_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3_var__u82_0_valid_out_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3_var__u82_0_stall_in_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3_var__u82_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb3_var__u82_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb3_var__u82_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb3_var__u82_0_stall_in_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb3_var__u82_0_valid_out_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb3_var__u82_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb3_var__u82),
	.data_out(rnode_389to390_bb3_var__u82_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb3_var__u82_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb3_var__u82_0_reg_390_fifo.DATA_WIDTH = 1;
defparam rnode_389to390_bb3_var__u82_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb3_var__u82_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb3_var__u82_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u82_stall_in = 1'b0;
assign rnode_389to390_bb3_var__u82_0_NO_SHIFT_REG = rnode_389to390_bb3_var__u82_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb3_var__u82_0_stall_in_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb3_var__u82_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb3_add192_i113_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb3_add192_i113_0_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb3_add192_i113_1_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb3_add192_i113_2_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb3_add192_i113_3_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb3_add192_i113_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_valid_out_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_stall_in_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3_add192_i113_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb3_add192_i113_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb3_add192_i113_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb3_add192_i113_0_stall_in_0_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb3_add192_i113_0_valid_out_0_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb3_add192_i113_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb3_add192_i113),
	.data_out(rnode_389to390_bb3_add192_i113_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb3_add192_i113_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb3_add192_i113_0_reg_390_fifo.DATA_WIDTH = 32;
defparam rnode_389to390_bb3_add192_i113_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb3_add192_i113_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb3_add192_i113_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add192_i113_stall_in = 1'b0;
assign rnode_389to390_bb3_add192_i113_0_stall_in_0_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb3_add192_i113_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb3_add192_i113_0_NO_SHIFT_REG = rnode_389to390_bb3_add192_i113_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb3_add192_i113_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb3_add192_i113_1_NO_SHIFT_REG = rnode_389to390_bb3_add192_i113_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb3_add192_i113_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb3_add192_i113_2_NO_SHIFT_REG = rnode_389to390_bb3_add192_i113_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb3_add192_i113_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb3_add192_i113_3_NO_SHIFT_REG = rnode_389to390_bb3_add192_i113_0_reg_390_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb3__26_i49_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to390_bb3__26_i49_0_stall_in_NO_SHIFT_REG;
 logic rnode_389to390_bb3__26_i49_0_NO_SHIFT_REG;
 logic rnode_389to390_bb3__26_i49_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to390_bb3__26_i49_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3__26_i49_0_valid_out_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3__26_i49_0_stall_in_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb3__26_i49_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb3__26_i49_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb3__26_i49_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb3__26_i49_0_stall_in_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb3__26_i49_0_valid_out_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb3__26_i49_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb3__26_i49),
	.data_out(rnode_389to390_bb3__26_i49_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb3__26_i49_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb3__26_i49_0_reg_390_fifo.DATA_WIDTH = 1;
defparam rnode_389to390_bb3__26_i49_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb3__26_i49_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb3__26_i49_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__26_i49_stall_in = 1'b0;
assign rnode_389to390_bb3__26_i49_0_NO_SHIFT_REG = rnode_389to390_bb3__26_i49_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb3__26_i49_0_stall_in_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb3__26_i49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_1_i_stall_local;
wire [31:0] local_bb3_reduction_1_i;

assign local_bb3_reduction_1_i = ((local_bb3_lnot_ext314_i & 32'h1) & (local_bb3_lor_ext_i & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb3_var__u82_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb3_var__u82_0_stall_in_NO_SHIFT_REG;
 logic rnode_390to391_bb3_var__u82_0_NO_SHIFT_REG;
 logic rnode_390to391_bb3_var__u82_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic rnode_390to391_bb3_var__u82_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_var__u82_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_var__u82_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_var__u82_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb3_var__u82_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb3_var__u82_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb3_var__u82_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb3_var__u82_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb3_var__u82_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in(rnode_389to390_bb3_var__u82_0_NO_SHIFT_REG),
	.data_out(rnode_390to391_bb3_var__u82_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb3_var__u82_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb3_var__u82_0_reg_391_fifo.DATA_WIDTH = 1;
defparam rnode_390to391_bb3_var__u82_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb3_var__u82_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb3_var__u82_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb3_var__u82_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_var__u82_0_NO_SHIFT_REG = rnode_390to391_bb3_var__u82_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb3_var__u82_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_var__u82_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and193_i114_valid_out;
wire local_bb3_and193_i114_stall_in;
wire local_bb3_and193_i114_inputs_ready;
wire local_bb3_and193_i114_stall_local;
wire [31:0] local_bb3_and193_i114;

assign local_bb3_and193_i114_inputs_ready = rnode_389to390_bb3_add192_i113_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_and193_i114 = (rnode_389to390_bb3_add192_i113_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb3_and193_i114_valid_out = 1'b1;
assign rnode_389to390_bb3_add192_i113_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and195_i115_valid_out;
wire local_bb3_and195_i115_stall_in;
wire local_bb3_and195_i115_inputs_ready;
wire local_bb3_and195_i115_stall_local;
wire [31:0] local_bb3_and195_i115;

assign local_bb3_and195_i115_inputs_ready = rnode_389to390_bb3_add192_i113_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_and195_i115 = (rnode_389to390_bb3_add192_i113_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb3_and195_i115_valid_out = 1'b1;
assign rnode_389to390_bb3_add192_i113_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and198_i116_valid_out;
wire local_bb3_and198_i116_stall_in;
wire local_bb3_and198_i116_inputs_ready;
wire local_bb3_and198_i116_stall_local;
wire [31:0] local_bb3_and198_i116;

assign local_bb3_and198_i116_inputs_ready = rnode_389to390_bb3_add192_i113_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_and198_i116 = (rnode_389to390_bb3_add192_i113_2_NO_SHIFT_REG & 32'h1);
assign local_bb3_and198_i116_valid_out = 1'b1;
assign rnode_389to390_bb3_add192_i113_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_and201_i117_stall_local;
wire [31:0] local_bb3_and201_i117;

assign local_bb3_and201_i117 = (rnode_389to390_bb3_add192_i113_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_390to392_bb3__26_i49_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to392_bb3__26_i49_0_stall_in_NO_SHIFT_REG;
 logic rnode_390to392_bb3__26_i49_0_NO_SHIFT_REG;
 logic rnode_390to392_bb3__26_i49_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_390to392_bb3__26_i49_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb3__26_i49_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb3__26_i49_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb3__26_i49_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_390to392_bb3__26_i49_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to392_bb3__26_i49_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to392_bb3__26_i49_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_390to392_bb3__26_i49_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_390to392_bb3__26_i49_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_389to390_bb3__26_i49_0_NO_SHIFT_REG),
	.data_out(rnode_390to392_bb3__26_i49_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_390to392_bb3__26_i49_0_reg_392_fifo.DEPTH = 2;
defparam rnode_390to392_bb3__26_i49_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_390to392_bb3__26_i49_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to392_bb3__26_i49_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_390to392_bb3__26_i49_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb3__26_i49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb3__26_i49_0_NO_SHIFT_REG = rnode_390to392_bb3__26_i49_0_reg_392_NO_SHIFT_REG;
assign rnode_390to392_bb3__26_i49_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb3__26_i49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_2_i_stall_local;
wire [31:0] local_bb3_reduction_2_i;

assign local_bb3_reduction_2_i = ((local_bb3_reduction_0_i & 32'h1) & (local_bb3_reduction_1_i & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb3_var__u82_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb3_var__u82_0_stall_in_NO_SHIFT_REG;
 logic rnode_391to392_bb3_var__u82_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3_var__u82_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_391to392_bb3_var__u82_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_var__u82_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_var__u82_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_var__u82_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb3_var__u82_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb3_var__u82_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb3_var__u82_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb3_var__u82_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb3_var__u82_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_390to391_bb3_var__u82_0_NO_SHIFT_REG),
	.data_out(rnode_391to392_bb3_var__u82_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb3_var__u82_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb3_var__u82_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_391to392_bb3_var__u82_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb3_var__u82_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb3_var__u82_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb3_var__u82_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_var__u82_0_NO_SHIFT_REG = rnode_391to392_bb3_var__u82_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb3_var__u82_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_var__u82_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb3_and193_i114_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and193_i114_0_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and193_i114_1_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and193_i114_2_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and193_i114_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_valid_out_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_stall_in_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and193_i114_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb3_and193_i114_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb3_and193_i114_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb3_and193_i114_0_stall_in_0_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb3_and193_i114_0_valid_out_0_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb3_and193_i114_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb3_and193_i114 & 32'hFFFFFFF)),
	.data_out(rnode_390to391_bb3_and193_i114_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb3_and193_i114_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb3_and193_i114_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb3_and193_i114_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb3_and193_i114_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb3_and193_i114_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and193_i114_stall_in = 1'b0;
assign rnode_390to391_bb3_and193_i114_0_stall_in_0_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and193_i114_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb3_and193_i114_0_NO_SHIFT_REG = rnode_390to391_bb3_and193_i114_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb3_and193_i114_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb3_and193_i114_1_NO_SHIFT_REG = rnode_390to391_bb3_and193_i114_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb3_and193_i114_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb3_and193_i114_2_NO_SHIFT_REG = rnode_390to391_bb3_and193_i114_0_reg_391_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb3_and195_i115_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and195_i115_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and195_i115_0_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and195_i115_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and195_i115_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and195_i115_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and195_i115_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and195_i115_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb3_and195_i115_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb3_and195_i115_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb3_and195_i115_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb3_and195_i115_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb3_and195_i115_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb3_and195_i115 & 32'h1F)),
	.data_out(rnode_390to391_bb3_and195_i115_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb3_and195_i115_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb3_and195_i115_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb3_and195_i115_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb3_and195_i115_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb3_and195_i115_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and195_i115_stall_in = 1'b0;
assign rnode_390to391_bb3_and195_i115_0_NO_SHIFT_REG = rnode_390to391_bb3_and195_i115_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb3_and195_i115_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and195_i115_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb3_and198_i116_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and198_i116_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and198_i116_0_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and198_i116_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3_and198_i116_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and198_i116_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and198_i116_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3_and198_i116_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb3_and198_i116_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb3_and198_i116_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb3_and198_i116_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb3_and198_i116_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb3_and198_i116_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb3_and198_i116 & 32'h1)),
	.data_out(rnode_390to391_bb3_and198_i116_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb3_and198_i116_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb3_and198_i116_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb3_and198_i116_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb3_and198_i116_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb3_and198_i116_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and198_i116_stall_in = 1'b0;
assign rnode_390to391_bb3_and198_i116_0_NO_SHIFT_REG = rnode_390to391_bb3_and198_i116_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb3_and198_i116_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and198_i116_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i_i118_stall_local;
wire [31:0] local_bb3_shr_i_i118;

assign local_bb3_shr_i_i118 = ((local_bb3_and201_i117 & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3__26_i49_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_2_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_valid_out_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_stall_in_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3__26_i49_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3__26_i49_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3__26_i49_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3__26_i49_0_stall_in_0_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3__26_i49_0_valid_out_0_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3__26_i49_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_390to392_bb3__26_i49_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb3__26_i49_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3__26_i49_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3__26_i49_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb3__26_i49_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3__26_i49_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3__26_i49_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb3__26_i49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__26_i49_0_stall_in_0_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__26_i49_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3__26_i49_0_NO_SHIFT_REG = rnode_392to393_bb3__26_i49_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3__26_i49_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3__26_i49_1_NO_SHIFT_REG = rnode_392to393_bb3__26_i49_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3__26_i49_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3__26_i49_2_NO_SHIFT_REG = rnode_392to393_bb3__26_i49_0_reg_393_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_add320_i_stall_local;
wire [31:0] local_bb3_add320_i;

assign local_bb3_add320_i = ((local_bb3_reduction_2_i & 32'h1) + local_bb3_or295_i);

// This section implements an unregistered operation.
// 
wire local_bb3_shr216_i139_stall_local;
wire [31:0] local_bb3_shr216_i139;

assign local_bb3_shr216_i139 = ((rnode_390to391_bb3_and193_i114_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__pre_i137_stall_local;
wire [31:0] local_bb3__pre_i137;

assign local_bb3__pre_i137 = ((rnode_390to391_bb3_and195_i115_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i_i119_stall_local;
wire [31:0] local_bb3_or_i_i119;

assign local_bb3_or_i_i119 = ((local_bb3_shr_i_i118 & 32'h3FFFFFF) | (local_bb3_and201_i117 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_cond292_i176_stall_local;
wire [31:0] local_bb3_cond292_i176;

assign local_bb3_cond292_i176 = (rnode_392to393_bb3__26_i49_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u90_stall_local;
wire [31:0] local_bb3_var__u90;

assign local_bb3_var__u90[31:1] = 31'h0;
assign local_bb3_var__u90[0] = rnode_392to393_bb3__26_i49_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u91_stall_local;
wire [31:0] local_bb3_var__u91;

assign local_bb3_var__u91 = local_bb3_add320_i;

// This section implements an unregistered operation.
// 
wire local_bb3_or219_i140_stall_local;
wire [31:0] local_bb3_or219_i140;

assign local_bb3_or219_i140 = ((local_bb3_shr216_i139 & 32'h7FFFFFF) | (rnode_390to391_bb3_and198_i116_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_tobool213_i138_stall_local;
wire local_bb3_tobool213_i138;

assign local_bb3_tobool213_i138 = ((local_bb3__pre_i137 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_shr1_i_i120_stall_local;
wire [31:0] local_bb3_shr1_i_i120;

assign local_bb3_shr1_i_i120 = ((local_bb3_or_i_i119 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext_i186_stall_local;
wire [31:0] local_bb3_lnot_ext_i186;

assign local_bb3_lnot_ext_i186 = ((local_bb3_var__u90 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3___valid_out;
wire local_bb3___stall_in;
wire local_bb3___inputs_ready;
wire local_bb3___stall_local;
wire [31:0] local_bb3__;

assign local_bb3___inputs_ready = (rnode_387to388_bb3_c0_ene7_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG & rnode_386to388_bb3_and269_i_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb3_resultSign_0_i_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb3_or2662_i_0_valid_out_1_NO_SHIFT_REG & rnode_387to388_bb3__26_i_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb3__26_i_0_valid_out_1_NO_SHIFT_REG & rnode_387to388_bb3__47_i_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb3_or2662_i_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb3__26_i_0_valid_out_2_NO_SHIFT_REG & rnode_387to388_bb3_or2662_i_0_valid_out_2_NO_SHIFT_REG & rnode_387to388_bb3_shr271_i_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb3__47_i_0_valid_out_1_NO_SHIFT_REG & rnode_387to388_bb3_cmp296_i_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb3_cmp299_i_0_valid_out_NO_SHIFT_REG);
assign local_bb3__ = (rnode_387to388_bb3_c0_ene7_0_NO_SHIFT_REG ? local_bb3_var__u91 : rnode_387to388_bb3_c0_ene6_0_NO_SHIFT_REG);
assign local_bb3___valid_out = 1'b1;
assign rnode_387to388_bb3_c0_ene7_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to388_bb3_and269_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_resultSign_0_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_or2662_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__26_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__26_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__47_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_or2662_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__26_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_or2662_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_shr271_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3__47_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_cmp296_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb3_cmp299_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__40_demorgan_i141_stall_local;
wire local_bb3__40_demorgan_i141;

assign local_bb3__40_demorgan_i141 = (rnode_389to391_bb3_cmp37_i36_0_NO_SHIFT_REG | local_bb3_tobool213_i138);

// This section implements an unregistered operation.
// 
wire local_bb3__42_i143_stall_local;
wire local_bb3__42_i143;

assign local_bb3__42_i143 = (local_bb3_tobool213_i138 & local_bb3_not_cmp37_i142);

// This section implements an unregistered operation.
// 
wire local_bb3_or2_i_i121_stall_local;
wire [31:0] local_bb3_or2_i_i121;

assign local_bb3_or2_i_i121 = ((local_bb3_shr1_i_i120 & 32'h1FFFFFF) | (local_bb3_or_i_i119 & 32'h7FFFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb3___0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb3___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3___0_NO_SHIFT_REG;
 logic rnode_388to389_bb3___0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb3___0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3___0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3___0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb3___0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb3___0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb3___0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb3___0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb3___0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb3___0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb3__),
	.data_out(rnode_388to389_bb3___0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb3___0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb3___0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb3___0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb3___0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb3___0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3___stall_in = 1'b0;
assign rnode_388to389_bb3___0_NO_SHIFT_REG = rnode_388to389_bb3___0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb3___0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb3___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__43_i144_stall_local;
wire [31:0] local_bb3__43_i144;

assign local_bb3__43_i144 = (local_bb3__42_i143 ? 32'h0 : (local_bb3__pre_i137 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_shr3_i_i122_stall_local;
wire [31:0] local_bb3_shr3_i_i122;

assign local_bb3_shr3_i_i122 = ((local_bb3_or2_i_i121 & 32'h7FFFFFF) >> 32'h4);

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_389to393_bb3___0_valid_out_NO_SHIFT_REG;
 logic rnode_389to393_bb3___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_389to393_bb3___0_NO_SHIFT_REG;
 logic rnode_389to393_bb3___0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to393_bb3___0_reg_393_NO_SHIFT_REG;
 logic rnode_389to393_bb3___0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_389to393_bb3___0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_389to393_bb3___0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_389to393_bb3___0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to393_bb3___0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to393_bb3___0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_389to393_bb3___0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_389to393_bb3___0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_388to389_bb3___0_NO_SHIFT_REG),
	.data_out(rnode_389to393_bb3___0_reg_393_NO_SHIFT_REG)
);

defparam rnode_389to393_bb3___0_reg_393_fifo.DEPTH = 4;
defparam rnode_389to393_bb3___0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_389to393_bb3___0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to393_bb3___0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_389to393_bb3___0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb3___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_389to393_bb3___0_NO_SHIFT_REG = rnode_389to393_bb3___0_reg_393_NO_SHIFT_REG;
assign rnode_389to393_bb3___0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_389to393_bb3___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_or4_i_i123_stall_local;
wire [31:0] local_bb3_or4_i_i123;

assign local_bb3_or4_i_i123 = ((local_bb3_shr3_i_i122 & 32'h7FFFFF) | (local_bb3_or2_i_i121 & 32'h7FFFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb3___0_valid_out_NO_SHIFT_REG;
 logic rnode_393to394_bb3___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb3___0_NO_SHIFT_REG;
 logic rnode_393to394_bb3___0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb3___0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb3___0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb3___0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb3___0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb3___0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb3___0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb3___0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb3___0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb3___0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in(rnode_389to393_bb3___0_NO_SHIFT_REG),
	.data_out(rnode_393to394_bb3___0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb3___0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb3___0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb3___0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb3___0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb3___0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to393_bb3___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb3___0_NO_SHIFT_REG = rnode_393to394_bb3___0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb3___0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb3___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_shr5_i_i124_stall_local;
wire [31:0] local_bb3_shr5_i_i124;

assign local_bb3_shr5_i_i124 = ((local_bb3_or4_i_i123 & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi1_stall_local;
wire [95:0] local_bb3_c0_exi1;

assign local_bb3_c0_exi1[31:0] = 32'bx;
assign local_bb3_c0_exi1[63:32] = rnode_393to394_bb3___0_NO_SHIFT_REG;
assign local_bb3_c0_exi1[95:64] = 32'bx;

// This section implements an unregistered operation.
// 
wire local_bb3_or6_i_i125_stall_local;
wire [31:0] local_bb3_or6_i_i125;

assign local_bb3_or6_i_i125 = ((local_bb3_shr5_i_i124 & 32'h7FFFF) | (local_bb3_or4_i_i123 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_shr7_i_i126_stall_local;
wire [31:0] local_bb3_shr7_i_i126;

assign local_bb3_shr7_i_i126 = ((local_bb3_or6_i_i125 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb3_or6_masked_i_i127_stall_local;
wire [31:0] local_bb3_or6_masked_i_i127;

assign local_bb3_or6_masked_i_i127 = ((local_bb3_or6_i_i125 & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_neg_i_i128_stall_local;
wire [31:0] local_bb3_neg_i_i128;

assign local_bb3_neg_i_i128 = ((local_bb3_or6_masked_i_i127 & 32'h7FFFFFF) | (local_bb3_shr7_i_i126 & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb3_and_i_i129_stall_local;
wire [31:0] local_bb3_and_i_i129;

assign local_bb3_and_i_i129 = ((local_bb3_neg_i_i128 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3__and_i_i129_valid_out;
wire local_bb3__and_i_i129_stall_in;
wire local_bb3__and_i_i129_inputs_ready;
wire local_bb3__and_i_i129_stall_local;
wire [31:0] local_bb3__and_i_i129;

thirtysix_six_comp local_bb3__and_i_i129_popcnt_instance (
	.data((local_bb3_and_i_i129 & 32'h7FFFFFF)),
	.sum(local_bb3__and_i_i129)
);


assign local_bb3__and_i_i129_inputs_ready = rnode_389to390_bb3_add192_i113_0_valid_out_3_NO_SHIFT_REG;
assign local_bb3__and_i_i129_valid_out = 1'b1;
assign rnode_389to390_bb3_add192_i113_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb3__and_i_i129_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3__and_i_i129_0_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3__and_i_i129_1_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3__and_i_i129_2_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb3__and_i_i129_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_valid_out_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_stall_in_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb3__and_i_i129_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb3__and_i_i129_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb3__and_i_i129_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb3__and_i_i129_0_stall_in_0_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb3__and_i_i129_0_valid_out_0_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb3__and_i_i129_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb3__and_i_i129 & 32'h3F)),
	.data_out(rnode_390to391_bb3__and_i_i129_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb3__and_i_i129_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb3__and_i_i129_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb3__and_i_i129_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb3__and_i_i129_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb3__and_i_i129_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__and_i_i129_stall_in = 1'b0;
assign rnode_390to391_bb3__and_i_i129_0_stall_in_0_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3__and_i_i129_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb3__and_i_i129_0_NO_SHIFT_REG = rnode_390to391_bb3__and_i_i129_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb3__and_i_i129_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb3__and_i_i129_1_NO_SHIFT_REG = rnode_390to391_bb3__and_i_i129_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb3__and_i_i129_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb3__and_i_i129_2_NO_SHIFT_REG = rnode_390to391_bb3__and_i_i129_0_reg_391_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_and9_i_i130_stall_local;
wire [31:0] local_bb3_and9_i_i130;

assign local_bb3_and9_i_i130 = ((rnode_390to391_bb3__and_i_i129_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb3_and203_i131_stall_local;
wire [31:0] local_bb3_and203_i131;

assign local_bb3_and203_i131 = ((rnode_390to391_bb3__and_i_i129_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb3_and206_i133_stall_local;
wire [31:0] local_bb3_and206_i133;

assign local_bb3_and206_i133 = ((rnode_390to391_bb3__and_i_i129_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb3_sub239_i152_stall_local;
wire [31:0] local_bb3_sub239_i152;

assign local_bb3_sub239_i152 = (32'h0 - (local_bb3_and9_i_i130 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb3_shl204_i132_stall_local;
wire [31:0] local_bb3_shl204_i132;

assign local_bb3_shl204_i132 = ((rnode_390to391_bb3_and193_i114_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb3_and203_i131 & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb3_cond244_i153_stall_local;
wire [31:0] local_bb3_cond244_i153;

assign local_bb3_cond244_i153 = (rnode_389to391_bb3_cmp37_i36_2_NO_SHIFT_REG ? local_bb3_sub239_i152 : (local_bb3__43_i144 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and205_i134_stall_local;
wire [31:0] local_bb3_and205_i134;

assign local_bb3_and205_i134 = (local_bb3_shl204_i132 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_add245_i154_stall_local;
wire [31:0] local_bb3_add245_i154;

assign local_bb3_add245_i154 = (local_bb3_cond244_i153 + (rnode_389to391_bb3_and17_i25_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb3_fold_i156_stall_local;
wire [31:0] local_bb3_fold_i156;

assign local_bb3_fold_i156 = (local_bb3_cond244_i153 + (rnode_389to391_bb3_shr16_i24_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb3_shl207_i135_stall_local;
wire [31:0] local_bb3_shl207_i135;

assign local_bb3_shl207_i135 = ((local_bb3_and205_i134 & 32'h7FFFFFF) << (local_bb3_and206_i133 & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb3_and250_i157_stall_local;
wire [31:0] local_bb3_and250_i157;

assign local_bb3_and250_i157 = (local_bb3_fold_i156 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and269_i168_stall_local;
wire [31:0] local_bb3_and269_i168;

assign local_bb3_and269_i168 = (local_bb3_fold_i156 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and208_i136_stall_local;
wire [31:0] local_bb3_and208_i136;

assign local_bb3_and208_i136 = (local_bb3_shl207_i135 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3__44_i145_stall_local;
wire [31:0] local_bb3__44_i145;

assign local_bb3__44_i145 = (local_bb3__40_demorgan_i141 ? (local_bb3_and208_i136 & 32'h7FFFFFF) : (local_bb3_or219_i140 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb3_and250_i157_valid_out;
wire local_bb3_and250_i157_stall_in;
wire local_bb3_and269_i168_valid_out;
wire local_bb3_and269_i168_stall_in;
wire local_bb3_add245_i154_valid_out;
wire local_bb3_add245_i154_stall_in;
wire local_bb3__45_i146_valid_out;
wire local_bb3__45_i146_stall_in;
wire local_bb3_not_cmp37_i142_valid_out_1;
wire local_bb3_not_cmp37_i142_stall_in_1;
wire local_bb3__45_i146_inputs_ready;
wire local_bb3__45_i146_stall_local;
wire [31:0] local_bb3__45_i146;

assign local_bb3__45_i146_inputs_ready = (rnode_389to391_bb3_shr16_i24_0_valid_out_NO_SHIFT_REG & rnode_389to391_bb3_and17_i25_0_valid_out_NO_SHIFT_REG & rnode_389to391_bb3_cmp37_i36_0_valid_out_2_NO_SHIFT_REG & rnode_389to391_bb3_cmp37_i36_0_valid_out_0_NO_SHIFT_REG & rnode_390to391_bb3_and193_i114_0_valid_out_2_NO_SHIFT_REG & rnode_389to391_bb3_cmp37_i36_0_valid_out_1_NO_SHIFT_REG & rnode_390to391_bb3_and195_i115_0_valid_out_NO_SHIFT_REG & rnode_390to391_bb3_and193_i114_0_valid_out_1_NO_SHIFT_REG & rnode_390to391_bb3_and198_i116_0_valid_out_NO_SHIFT_REG & rnode_390to391_bb3_and193_i114_0_valid_out_0_NO_SHIFT_REG & rnode_390to391_bb3__and_i_i129_0_valid_out_1_NO_SHIFT_REG & rnode_390to391_bb3__and_i_i129_0_valid_out_2_NO_SHIFT_REG & rnode_390to391_bb3__and_i_i129_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3__45_i146 = (local_bb3__42_i143 ? (rnode_390to391_bb3_and193_i114_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb3__44_i145 & 32'h7FFFFFF));
assign local_bb3_and250_i157_valid_out = 1'b1;
assign local_bb3_and269_i168_valid_out = 1'b1;
assign local_bb3_add245_i154_valid_out = 1'b1;
assign local_bb3__45_i146_valid_out = 1'b1;
assign local_bb3_not_cmp37_i142_valid_out_1 = 1'b1;
assign rnode_389to391_bb3_shr16_i24_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_and17_i25_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_cmp37_i36_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_cmp37_i36_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and193_i114_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb3_cmp37_i36_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and195_i115_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and193_i114_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and198_i116_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3_and193_i114_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3__and_i_i129_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3__and_i_i129_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb3__and_i_i129_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb3_and250_i157_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and250_i157_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3_and250_i157_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and250_i157_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3_and250_i157_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and250_i157_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and250_i157_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_and250_i157_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb3_and250_i157_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb3_and250_i157_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb3_and250_i157_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb3_and250_i157_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb3_and250_i157_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb3_and250_i157 & 32'hFF)),
	.data_out(rnode_391to392_bb3_and250_i157_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb3_and250_i157_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb3_and250_i157_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb3_and250_i157_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb3_and250_i157_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb3_and250_i157_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and250_i157_stall_in = 1'b0;
assign rnode_391to392_bb3_and250_i157_0_NO_SHIFT_REG = rnode_391to392_bb3_and250_i157_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb3_and250_i157_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_and250_i157_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_391to393_bb3_and269_i168_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to393_bb3_and269_i168_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to393_bb3_and269_i168_0_NO_SHIFT_REG;
 logic rnode_391to393_bb3_and269_i168_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to393_bb3_and269_i168_0_reg_393_NO_SHIFT_REG;
 logic rnode_391to393_bb3_and269_i168_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_391to393_bb3_and269_i168_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_391to393_bb3_and269_i168_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_391to393_bb3_and269_i168_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to393_bb3_and269_i168_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to393_bb3_and269_i168_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_391to393_bb3_and269_i168_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_391to393_bb3_and269_i168_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in((local_bb3_and269_i168 & 32'hFF800000)),
	.data_out(rnode_391to393_bb3_and269_i168_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_391to393_bb3_and269_i168_0_reg_393_fifo.DEPTH = 2;
defparam rnode_391to393_bb3_and269_i168_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_391to393_bb3_and269_i168_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to393_bb3_and269_i168_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_391to393_bb3_and269_i168_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_and269_i168_stall_in = 1'b0;
assign rnode_391to393_bb3_and269_i168_0_NO_SHIFT_REG = rnode_391to393_bb3_and269_i168_0_reg_393_NO_SHIFT_REG;
assign rnode_391to393_bb3_and269_i168_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_391to393_bb3_and269_i168_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb3_add245_i154_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3_add245_i154_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3_add245_i154_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3_add245_i154_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_391to392_bb3_add245_i154_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3_add245_i154_1_NO_SHIFT_REG;
 logic rnode_391to392_bb3_add245_i154_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3_add245_i154_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_add245_i154_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_add245_i154_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_add245_i154_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb3_add245_i154_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb3_add245_i154_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb3_add245_i154_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb3_add245_i154_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb3_add245_i154_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(local_bb3_add245_i154),
	.data_out(rnode_391to392_bb3_add245_i154_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb3_add245_i154_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb3_add245_i154_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb3_add245_i154_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb3_add245_i154_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb3_add245_i154_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add245_i154_stall_in = 1'b0;
assign rnode_391to392_bb3_add245_i154_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_add245_i154_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb3_add245_i154_0_NO_SHIFT_REG = rnode_391to392_bb3_add245_i154_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb3_add245_i154_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb3_add245_i154_1_NO_SHIFT_REG = rnode_391to392_bb3_add245_i154_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb3__45_i146_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3__45_i146_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3__45_i146_1_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3__45_i146_2_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb3__45_i146_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3__45_i146_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb3__45_i146_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb3__45_i146_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb3__45_i146_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb3__45_i146_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb3__45_i146_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb3__45_i146 & 32'hFFFFFFF)),
	.data_out(rnode_391to392_bb3__45_i146_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb3__45_i146_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb3__45_i146_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb3__45_i146_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb3__45_i146_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb3__45_i146_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__45_i146_stall_in = 1'b0;
assign rnode_391to392_bb3__45_i146_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3__45_i146_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb3__45_i146_0_NO_SHIFT_REG = rnode_391to392_bb3__45_i146_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb3__45_i146_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb3__45_i146_1_NO_SHIFT_REG = rnode_391to392_bb3__45_i146_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb3__45_i146_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb3__45_i146_2_NO_SHIFT_REG = rnode_391to392_bb3__45_i146_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb3_not_cmp37_i142_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb3_not_cmp37_i142_0_stall_in_NO_SHIFT_REG;
 logic rnode_391to392_bb3_not_cmp37_i142_0_NO_SHIFT_REG;
 logic rnode_391to392_bb3_not_cmp37_i142_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_391to392_bb3_not_cmp37_i142_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_not_cmp37_i142_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_not_cmp37_i142_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb3_not_cmp37_i142_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb3_not_cmp37_i142_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb3_not_cmp37_i142_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb3_not_cmp37_i142_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb3_not_cmp37_i142_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb3_not_cmp37_i142_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(local_bb3_not_cmp37_i142),
	.data_out(rnode_391to392_bb3_not_cmp37_i142_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb3_not_cmp37_i142_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb3_not_cmp37_i142_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_391to392_bb3_not_cmp37_i142_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb3_not_cmp37_i142_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb3_not_cmp37_i142_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_not_cmp37_i142_stall_in_1 = 1'b0;
assign rnode_391to392_bb3_not_cmp37_i142_0_NO_SHIFT_REG = rnode_391to392_bb3_not_cmp37_i142_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb3_not_cmp37_i142_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_not_cmp37_i142_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_notrhs_i159_stall_local;
wire local_bb3_notrhs_i159;

assign local_bb3_notrhs_i159 = ((rnode_391to392_bb3_and250_i157_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_shl273_i169_stall_local;
wire [31:0] local_bb3_shl273_i169;

assign local_bb3_shl273_i169 = ((rnode_391to393_bb3_and269_i168_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb3_and247_i155_stall_local;
wire [31:0] local_bb3_and247_i155;

assign local_bb3_and247_i155 = (rnode_391to392_bb3_add245_i154_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp258_i162_stall_local;
wire local_bb3_cmp258_i162;

assign local_bb3_cmp258_i162 = ($signed(rnode_391to392_bb3_add245_i154_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb3_and225_i147_stall_local;
wire [31:0] local_bb3_and225_i147;

assign local_bb3_and225_i147 = ((rnode_391to392_bb3__45_i146_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and270_i165_stall_local;
wire [31:0] local_bb3_and270_i165;

assign local_bb3_and270_i165 = ((rnode_391to392_bb3__45_i146_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb3_shr271_i166_valid_out;
wire local_bb3_shr271_i166_stall_in;
wire local_bb3_shr271_i166_inputs_ready;
wire local_bb3_shr271_i166_stall_local;
wire [31:0] local_bb3_shr271_i166;

assign local_bb3_shr271_i166_inputs_ready = rnode_391to392_bb3__45_i146_0_valid_out_2_NO_SHIFT_REG;
assign local_bb3_shr271_i166 = ((rnode_391to392_bb3__45_i146_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb3_shr271_i166_valid_out = 1'b1;
assign rnode_391to392_bb3__45_i146_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_notlhs_i158_stall_local;
wire local_bb3_notlhs_i158;

assign local_bb3_notlhs_i158 = ((local_bb3_and247_i155 & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp226_i148_stall_local;
wire local_bb3_cmp226_i148;

assign local_bb3_cmp226_i148 = ((local_bb3_and225_i147 & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp296_i180_stall_local;
wire local_bb3_cmp296_i180;

assign local_bb3_cmp296_i180 = ((local_bb3_and270_i165 & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp296_i180_valid_out;
wire local_bb3_cmp296_i180_stall_in;
wire local_bb3_cmp299_i181_valid_out;
wire local_bb3_cmp299_i181_stall_in;
wire local_bb3_cmp299_i181_inputs_ready;
wire local_bb3_cmp299_i181_stall_local;
wire local_bb3_cmp299_i181;

assign local_bb3_cmp299_i181_inputs_ready = rnode_391to392_bb3__45_i146_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_cmp299_i181 = ((local_bb3_and270_i165 & 32'h7) == 32'h4);
assign local_bb3_cmp296_i180_valid_out = 1'b1;
assign local_bb3_cmp299_i181_valid_out = 1'b1;
assign rnode_391to392_bb3__45_i146_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3_shr271_i166_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb3_shr271_i166_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb3_shr271_i166_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_shr271_i166_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb3_shr271_i166_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_shr271_i166_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_shr271_i166_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_shr271_i166_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3_shr271_i166_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3_shr271_i166_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3_shr271_i166_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3_shr271_i166_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3_shr271_i166_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in((local_bb3_shr271_i166 & 32'h1FFFFFF)),
	.data_out(rnode_392to393_bb3_shr271_i166_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3_shr271_i166_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3_shr271_i166_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_392to393_bb3_shr271_i166_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3_shr271_i166_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3_shr271_i166_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_shr271_i166_stall_in = 1'b0;
assign rnode_392to393_bb3_shr271_i166_0_NO_SHIFT_REG = rnode_392to393_bb3_shr271_i166_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_shr271_i166_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_shr271_i166_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_not__46_i160_stall_local;
wire local_bb3_not__46_i160;

assign local_bb3_not__46_i160 = (local_bb3_notrhs_i159 | local_bb3_notlhs_i158);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp226_not_i149_stall_local;
wire local_bb3_cmp226_not_i149;

assign local_bb3_cmp226_not_i149 = (local_bb3_cmp226_i148 ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3_cmp296_i180_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp296_i180_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp296_i180_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp296_i180_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp296_i180_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp296_i180_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp296_i180_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp296_i180_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3_cmp296_i180_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3_cmp296_i180_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3_cmp296_i180_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3_cmp296_i180_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3_cmp296_i180_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb3_cmp296_i180),
	.data_out(rnode_392to393_bb3_cmp296_i180_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3_cmp296_i180_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3_cmp296_i180_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb3_cmp296_i180_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3_cmp296_i180_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3_cmp296_i180_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp296_i180_stall_in = 1'b0;
assign rnode_392to393_bb3_cmp296_i180_0_NO_SHIFT_REG = rnode_392to393_bb3_cmp296_i180_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_cmp296_i180_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_cmp296_i180_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3_cmp299_i181_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp299_i181_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp299_i181_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp299_i181_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp299_i181_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp299_i181_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp299_i181_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_cmp299_i181_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3_cmp299_i181_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3_cmp299_i181_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3_cmp299_i181_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3_cmp299_i181_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3_cmp299_i181_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb3_cmp299_i181),
	.data_out(rnode_392to393_bb3_cmp299_i181_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3_cmp299_i181_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3_cmp299_i181_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb3_cmp299_i181_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3_cmp299_i181_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3_cmp299_i181_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp299_i181_stall_in = 1'b0;
assign rnode_392to393_bb3_cmp299_i181_0_NO_SHIFT_REG = rnode_392to393_bb3_cmp299_i181_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_cmp299_i181_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_cmp299_i181_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_and272_i167_stall_local;
wire [31:0] local_bb3_and272_i167;

assign local_bb3_and272_i167 = ((rnode_392to393_bb3_shr271_i166_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3__47_i161_stall_local;
wire local_bb3__47_i161;

assign local_bb3__47_i161 = (local_bb3_cmp226_i148 | local_bb3_not__46_i160);

// This section implements an unregistered operation.
// 
wire local_bb3_brmerge12_i150_stall_local;
wire local_bb3_brmerge12_i150;

assign local_bb3_brmerge12_i150 = (local_bb3_cmp226_not_i149 | rnode_391to392_bb3_not_cmp37_i142_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot262__i163_stall_local;
wire local_bb3_lnot262__i163;

assign local_bb3_lnot262__i163 = (local_bb3_cmp258_i162 & local_bb3_cmp226_not_i149);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp29649_i184_stall_local;
wire [31:0] local_bb3_cmp29649_i184;

assign local_bb3_cmp29649_i184[31:1] = 31'h0;
assign local_bb3_cmp29649_i184[0] = rnode_392to393_bb3_cmp296_i180_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_conv300_i182_stall_local;
wire [31:0] local_bb3_conv300_i182;

assign local_bb3_conv300_i182[31:1] = 31'h0;
assign local_bb3_conv300_i182[0] = rnode_392to393_bb3_cmp299_i181_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or274_i170_stall_local;
wire [31:0] local_bb3_or274_i170;

assign local_bb3_or274_i170 = ((local_bb3_and272_i167 & 32'h7FFFFF) | (local_bb3_shl273_i169 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb3_resultSign_0_i151_stall_local;
wire [31:0] local_bb3_resultSign_0_i151;

assign local_bb3_resultSign_0_i151 = (local_bb3_brmerge12_i150 ? (rnode_391to392_bb3_and35_i34_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_resultSign_0_i151_valid_out;
wire local_bb3_resultSign_0_i151_stall_in;
wire local_bb3__47_i161_valid_out;
wire local_bb3__47_i161_stall_in;
wire local_bb3_or2662_i164_valid_out;
wire local_bb3_or2662_i164_stall_in;
wire local_bb3_or2662_i164_inputs_ready;
wire local_bb3_or2662_i164_stall_local;
wire local_bb3_or2662_i164;

assign local_bb3_or2662_i164_inputs_ready = (rnode_391to392_bb3_and35_i34_0_valid_out_NO_SHIFT_REG & rnode_391to392_bb3_not_cmp37_i142_0_valid_out_NO_SHIFT_REG & rnode_391to392_bb3_add245_i154_0_valid_out_0_NO_SHIFT_REG & rnode_391to392_bb3_and250_i157_0_valid_out_NO_SHIFT_REG & rnode_391to392_bb3__45_i146_0_valid_out_0_NO_SHIFT_REG & rnode_391to392_bb3_add245_i154_0_valid_out_1_NO_SHIFT_REG & rnode_391to392_bb3_var__u82_0_valid_out_NO_SHIFT_REG);
assign local_bb3_or2662_i164 = (rnode_391to392_bb3_var__u82_0_NO_SHIFT_REG | local_bb3_lnot262__i163);
assign local_bb3_resultSign_0_i151_valid_out = 1'b1;
assign local_bb3__47_i161_valid_out = 1'b1;
assign local_bb3_or2662_i164_valid_out = 1'b1;
assign rnode_391to392_bb3_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_not_cmp37_i142_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_add245_i154_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_and250_i157_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3__45_i146_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_add245_i154_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb3_var__u82_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3_resultSign_0_i151_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb3_resultSign_0_i151_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb3_resultSign_0_i151_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_resultSign_0_i151_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb3_resultSign_0_i151_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_resultSign_0_i151_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_resultSign_0_i151_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_resultSign_0_i151_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3_resultSign_0_i151_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3_resultSign_0_i151_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3_resultSign_0_i151_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3_resultSign_0_i151_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3_resultSign_0_i151_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in((local_bb3_resultSign_0_i151 & 32'h80000000)),
	.data_out(rnode_392to393_bb3_resultSign_0_i151_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3_resultSign_0_i151_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3_resultSign_0_i151_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_392to393_bb3_resultSign_0_i151_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3_resultSign_0_i151_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3_resultSign_0_i151_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_resultSign_0_i151_stall_in = 1'b0;
assign rnode_392to393_bb3_resultSign_0_i151_0_NO_SHIFT_REG = rnode_392to393_bb3_resultSign_0_i151_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_resultSign_0_i151_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_resultSign_0_i151_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3__47_i161_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_valid_out_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_stall_in_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3__47_i161_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3__47_i161_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3__47_i161_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3__47_i161_0_stall_in_0_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3__47_i161_0_valid_out_0_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3__47_i161_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb3__47_i161),
	.data_out(rnode_392to393_bb3__47_i161_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3__47_i161_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3__47_i161_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb3__47_i161_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3__47_i161_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3__47_i161_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__47_i161_stall_in = 1'b0;
assign rnode_392to393_bb3__47_i161_0_stall_in_0_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__47_i161_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3__47_i161_0_NO_SHIFT_REG = rnode_392to393_bb3__47_i161_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3__47_i161_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3__47_i161_1_NO_SHIFT_REG = rnode_392to393_bb3__47_i161_0_reg_393_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb3_or2662_i164_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_1_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_2_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_valid_out_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_stall_in_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb3_or2662_i164_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb3_or2662_i164_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb3_or2662_i164_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb3_or2662_i164_0_stall_in_0_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb3_or2662_i164_0_valid_out_0_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb3_or2662_i164_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb3_or2662_i164),
	.data_out(rnode_392to393_bb3_or2662_i164_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb3_or2662_i164_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb3_or2662_i164_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb3_or2662_i164_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb3_or2662_i164_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb3_or2662_i164_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_or2662_i164_stall_in = 1'b0;
assign rnode_392to393_bb3_or2662_i164_0_stall_in_0_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_or2662_i164_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3_or2662_i164_0_NO_SHIFT_REG = rnode_392to393_bb3_or2662_i164_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_or2662_i164_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3_or2662_i164_1_NO_SHIFT_REG = rnode_392to393_bb3_or2662_i164_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb3_or2662_i164_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb3_or2662_i164_2_NO_SHIFT_REG = rnode_392to393_bb3_or2662_i164_0_reg_393_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or275_i171_stall_local;
wire [31:0] local_bb3_or275_i171;

assign local_bb3_or275_i171 = ((local_bb3_or274_i170 & 32'h7FFFFFFF) | (rnode_392to393_bb3_resultSign_0_i151_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb3_var__u92_stall_local;
wire [31:0] local_bb3_var__u92;

assign local_bb3_var__u92[31:1] = 31'h0;
assign local_bb3_var__u92[0] = rnode_392to393_bb3__47_i161_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_or2804_i172_stall_local;
wire local_bb3_or2804_i172;

assign local_bb3_or2804_i172 = (rnode_392to393_bb3__47_i161_0_NO_SHIFT_REG | rnode_392to393_bb3_or2662_i164_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_or2875_i174_stall_local;
wire local_bb3_or2875_i174;

assign local_bb3_or2875_i174 = (rnode_392to393_bb3_or2662_i164_1_NO_SHIFT_REG | rnode_392to393_bb3__26_i49_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u93_stall_local;
wire [31:0] local_bb3_var__u93;

assign local_bb3_var__u93[31:1] = 31'h0;
assign local_bb3_var__u93[0] = rnode_392to393_bb3_or2662_i164_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext314_i188_stall_local;
wire [31:0] local_bb3_lnot_ext314_i188;

assign local_bb3_lnot_ext314_i188 = ((local_bb3_var__u92 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_cond282_i173_stall_local;
wire [31:0] local_bb3_cond282_i173;

assign local_bb3_cond282_i173 = (local_bb3_or2804_i172 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cond289_i175_stall_local;
wire [31:0] local_bb3_cond289_i175;

assign local_bb3_cond289_i175 = (local_bb3_or2875_i174 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot_ext310_i187_stall_local;
wire [31:0] local_bb3_lnot_ext310_i187;

assign local_bb3_lnot_ext310_i187 = ((local_bb3_var__u93 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb3_and293_i177_stall_local;
wire [31:0] local_bb3_and293_i177;

assign local_bb3_and293_i177 = ((local_bb3_cond282_i173 | 32'h80000000) & local_bb3_or275_i171);

// This section implements an unregistered operation.
// 
wire local_bb3_or294_i178_stall_local;
wire [31:0] local_bb3_or294_i178;

assign local_bb3_or294_i178 = ((local_bb3_cond289_i175 & 32'h7F800000) | (local_bb3_cond292_i176 & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_0_i189_stall_local;
wire [31:0] local_bb3_reduction_0_i189;

assign local_bb3_reduction_0_i189 = ((local_bb3_lnot_ext310_i187 & 32'h1) & (local_bb3_lnot_ext_i186 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_and302_i183_stall_local;
wire [31:0] local_bb3_and302_i183;

assign local_bb3_and302_i183 = ((local_bb3_conv300_i182 & 32'h1) & local_bb3_and293_i177);

// This section implements an unregistered operation.
// 
wire local_bb3_or295_i179_stall_local;
wire [31:0] local_bb3_or295_i179;

assign local_bb3_or295_i179 = ((local_bb3_or294_i178 & 32'h7FC00000) | local_bb3_and293_i177);

// This section implements an unregistered operation.
// 
wire local_bb3_lor_ext_i185_stall_local;
wire [31:0] local_bb3_lor_ext_i185;

assign local_bb3_lor_ext_i185 = ((local_bb3_cmp29649_i184 & 32'h1) | (local_bb3_and302_i183 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_1_i190_stall_local;
wire [31:0] local_bb3_reduction_1_i190;

assign local_bb3_reduction_1_i190 = ((local_bb3_lnot_ext314_i188 & 32'h1) & (local_bb3_lor_ext_i185 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_reduction_2_i191_stall_local;
wire [31:0] local_bb3_reduction_2_i191;

assign local_bb3_reduction_2_i191 = ((local_bb3_reduction_0_i189 & 32'h1) & (local_bb3_reduction_1_i190 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb3_add320_i192_stall_local;
wire [31:0] local_bb3_add320_i192;

assign local_bb3_add320_i192 = ((local_bb3_reduction_2_i191 & 32'h1) + local_bb3_or295_i179);

// This section implements an unregistered operation.
// 
wire local_bb3_var__u94_stall_local;
wire [31:0] local_bb3_var__u94;

assign local_bb3_var__u94 = local_bb3_add320_i192;

// This section implements an unregistered operation.
// 
wire local_bb3__32_valid_out;
wire local_bb3__32_stall_in;
wire local_bb3__32_inputs_ready;
wire local_bb3__32_stall_local;
wire [31:0] local_bb3__32;

assign local_bb3__32_inputs_ready = (rnode_392to393_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG & rnode_391to393_bb3_and269_i168_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb3_resultSign_0_i151_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb3_or2662_i164_0_valid_out_1_NO_SHIFT_REG & rnode_392to393_bb3__26_i49_0_valid_out_0_NO_SHIFT_REG & rnode_392to393_bb3__26_i49_0_valid_out_1_NO_SHIFT_REG & rnode_392to393_bb3__47_i161_0_valid_out_0_NO_SHIFT_REG & rnode_392to393_bb3_or2662_i164_0_valid_out_0_NO_SHIFT_REG & rnode_392to393_bb3__26_i49_0_valid_out_2_NO_SHIFT_REG & rnode_392to393_bb3_or2662_i164_0_valid_out_2_NO_SHIFT_REG & rnode_392to393_bb3_shr271_i166_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb3__47_i161_0_valid_out_1_NO_SHIFT_REG & rnode_392to393_bb3_cmp296_i180_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb3_cmp299_i181_0_valid_out_NO_SHIFT_REG);
assign local_bb3__32 = (rnode_392to393_bb3_c0_ene7_0_NO_SHIFT_REG ? local_bb3_var__u94 : rnode_392to393_bb3_c0_ene5_0_NO_SHIFT_REG);
assign local_bb3__32_valid_out = 1'b1;
assign rnode_392to393_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to393_bb3_and269_i168_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_resultSign_0_i151_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_or2662_i164_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__26_i49_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__26_i49_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__47_i161_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_or2662_i164_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__26_i49_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_or2662_i164_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_shr271_i166_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3__47_i161_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_cmp296_i180_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb3_cmp299_i181_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb3__32_0_valid_out_NO_SHIFT_REG;
 logic rnode_393to394_bb3__32_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb3__32_0_NO_SHIFT_REG;
 logic rnode_393to394_bb3__32_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb3__32_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb3__32_0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb3__32_0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb3__32_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb3__32_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb3__32_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb3__32_0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb3__32_0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb3__32_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in(local_bb3__32),
	.data_out(rnode_393to394_bb3__32_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb3__32_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb3__32_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb3__32_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb3__32_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb3__32_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__32_stall_in = 1'b0;
assign rnode_393to394_bb3__32_0_NO_SHIFT_REG = rnode_393to394_bb3__32_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb3__32_0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb3__32_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi2_valid_out;
wire local_bb3_c0_exi2_stall_in;
wire local_bb3_c0_exi2_inputs_ready;
wire local_bb3_c0_exi2_stall_local;
wire [95:0] local_bb3_c0_exi2;

assign local_bb3_c0_exi2_inputs_ready = (rnode_393to394_bb3___0_valid_out_NO_SHIFT_REG & rnode_393to394_bb3__32_0_valid_out_NO_SHIFT_REG);
assign local_bb3_c0_exi2[63:0] = local_bb3_c0_exi1[63:0];
assign local_bb3_c0_exi2[95:64] = rnode_393to394_bb3__32_0_NO_SHIFT_REG;
assign local_bb3_c0_exi2_valid_out = 1'b1;
assign rnode_393to394_bb3___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb3__32_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb3_c0_exit_c0_exi2_inputs_ready;
 reg local_bb3_c0_exit_c0_exi2_valid_out_0_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi2_stall_in_0;
 reg local_bb3_c0_exit_c0_exi2_valid_out_1_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi2_stall_in_1;
 reg [95:0] local_bb3_c0_exit_c0_exi2_NO_SHIFT_REG;
wire [95:0] local_bb3_c0_exit_c0_exi2_in;
wire local_bb3_c0_exit_c0_exi2_valid;
wire local_bb3_c0_exit_c0_exi2_causedstall;

acl_stall_free_sink local_bb3_c0_exit_c0_exi2_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb3_c0_exi2),
	.data_out(local_bb3_c0_exit_c0_exi2_in),
	.input_accepted(local_bb3_c0_enter_c0_eni7_input_accepted),
	.valid_out(local_bb3_c0_exit_c0_exi2_valid),
	.stall_in(~(local_bb3_c0_exit_c0_exi2_output_regs_ready)),
	.stall_entry(local_bb3_c0_exit_c0_exi2_entry_stall),
	.valid_in(local_bb3_c0_exit_c0_exi2_valid_in),
	.IIphases(local_bb3_c0_exit_c0_exi2_phases),
	.inc_pipelined_thread(local_bb3_c0_enter_c0_eni7_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb3_c0_enter_c0_eni7_dec_pipelined_thread)
);

defparam local_bb3_c0_exit_c0_exi2_instance.DATA_WIDTH = 96;
defparam local_bb3_c0_exit_c0_exi2_instance.PIPELINE_DEPTH = 68;
defparam local_bb3_c0_exit_c0_exi2_instance.SHARINGII = 1;
defparam local_bb3_c0_exit_c0_exi2_instance.SCHEDULEII = 1;
defparam local_bb3_c0_exit_c0_exi2_instance.ALWAYS_THROTTLE = 0;

assign local_bb3_c0_exit_c0_exi2_inputs_ready = 1'b1;
assign local_bb3_c0_exit_c0_exi2_output_regs_ready = ((~(local_bb3_c0_exit_c0_exi2_valid_out_0_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi2_stall_in_0)) & (~(local_bb3_c0_exit_c0_exi2_valid_out_1_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi2_stall_in_1)));
assign local_bb3_c0_exit_c0_exi2_valid_in = SFC_1_VALID_393_394_0_NO_SHIFT_REG;
assign local_bb3_c0_exi2_stall_in = 1'b0;
assign SFC_1_VALID_393_394_0_stall_in = 1'b0;
assign local_bb3_c0_exit_c0_exi2_causedstall = (1'b1 && (1'b0 && !(~(local_bb3_c0_exit_c0_exi2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_c0_exit_c0_exi2_NO_SHIFT_REG <= 'x;
		local_bb3_c0_exit_c0_exi2_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi2_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_c0_exit_c0_exi2_output_regs_ready)
		begin
			local_bb3_c0_exit_c0_exi2_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi2_in;
			local_bb3_c0_exit_c0_exi2_valid_out_0_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi2_valid;
			local_bb3_c0_exit_c0_exi2_valid_out_1_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi2_valid;
		end
		else
		begin
			if (~(local_bb3_c0_exit_c0_exi2_stall_in_0))
			begin
				local_bb3_c0_exit_c0_exi2_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi2_stall_in_1))
			begin
				local_bb3_c0_exit_c0_exi2_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe1_stall_local;
wire [31:0] local_bb3_c0_exe1;

assign local_bb3_c0_exe1 = local_bb3_c0_exit_c0_exi2_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe2_valid_out;
wire local_bb3_c0_exe2_stall_in;
wire local_bb3_c0_exe1_valid_out;
wire local_bb3_c0_exe1_stall_in;
wire local_bb3_c0_exe2_inputs_ready;
wire local_bb3_c0_exe2_stall_local;
wire [31:0] local_bb3_c0_exe2;

assign local_bb3_c0_exe2_inputs_ready = (local_bb3_c0_exit_c0_exi2_valid_out_1_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi2_valid_out_0_NO_SHIFT_REG);
assign local_bb3_c0_exe2 = local_bb3_c0_exit_c0_exi2_NO_SHIFT_REG[95:64];
assign local_bb3_c0_exe2_stall_local = (local_bb3_c0_exe2_stall_in | local_bb3_c0_exe1_stall_in);
assign local_bb3_c0_exe2_valid_out = local_bb3_c0_exe2_inputs_ready;
assign local_bb3_c0_exe1_valid_out = local_bb3_c0_exe2_inputs_ready;
assign local_bb3_c0_exit_c0_exi2_stall_in_1 = (local_bb3_c0_exe2_stall_local | ~(local_bb3_c0_exe2_inputs_ready));
assign local_bb3_c0_exit_c0_exi2_stall_in_0 = (local_bb3_c0_exe2_stall_local | ~(local_bb3_c0_exe2_inputs_ready));

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_idxprom_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_ld__0_reg_NO_SHIFT_REG;
 reg lvb_cmp_0_reg_NO_SHIFT_REG;
 reg lvb_var__u8_0_reg_NO_SHIFT_REG;
 reg [63:0] lvb_indvars_iv29_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_sub25_add24_0_reg_NO_SHIFT_REG;
 reg [63:0] lvb_arrayidx43_0_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb3_indvars_iv_next_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe1_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe2_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb3_c0_exe2_valid_out & local_bb3_c0_exe1_valid_out & local_bb3_var__u11_valid_out & rnode_397to399_bb3_indvars_iv_next_0_valid_out_NO_SHIFT_REG & rcnode_398to399_rc0_idxprom_0_valid_out_0_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb3_c0_exe2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_var__u11_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_397to399_bb3_indvars_iv_next_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_398to399_rc0_idxprom_0_stall_in_0_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_idxprom_0 = lvb_idxprom_0_reg_NO_SHIFT_REG;
assign lvb_idxprom_1 = lvb_idxprom_0_reg_NO_SHIFT_REG;
assign lvb_ld__0 = lvb_ld__0_reg_NO_SHIFT_REG;
assign lvb_ld__1 = lvb_ld__0_reg_NO_SHIFT_REG;
assign lvb_cmp_0 = lvb_cmp_0_reg_NO_SHIFT_REG;
assign lvb_cmp_1 = lvb_cmp_0_reg_NO_SHIFT_REG;
assign lvb_var__u8_0 = lvb_var__u8_0_reg_NO_SHIFT_REG;
assign lvb_var__u8_1 = lvb_var__u8_0_reg_NO_SHIFT_REG;
assign lvb_indvars_iv29_0 = lvb_indvars_iv29_0_reg_NO_SHIFT_REG;
assign lvb_indvars_iv29_1 = lvb_indvars_iv29_0_reg_NO_SHIFT_REG;
assign lvb_sub25_add24_0 = lvb_sub25_add24_0_reg_NO_SHIFT_REG;
assign lvb_sub25_add24_1 = lvb_sub25_add24_0_reg_NO_SHIFT_REG;
assign lvb_arrayidx43_0 = lvb_arrayidx43_0_reg_NO_SHIFT_REG;
assign lvb_arrayidx43_1 = lvb_arrayidx43_0_reg_NO_SHIFT_REG;
assign lvb_bb3_indvars_iv_next_0 = lvb_bb3_indvars_iv_next_0_reg_NO_SHIFT_REG;
assign lvb_bb3_indvars_iv_next_1 = lvb_bb3_indvars_iv_next_0_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe1_0 = lvb_bb3_c0_exe1_0_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe1_1 = lvb_bb3_c0_exe1_0_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe2_0 = lvb_bb3_c0_exe2_0_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe2_1 = lvb_bb3_c0_exe2_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0_0 = lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0_1 = lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1_0 = lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1_1 = lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
assign lvb_input_acl_hw_wg_id_0 = lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG;
assign lvb_input_acl_hw_wg_id_1 = lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_idxprom_0_reg_NO_SHIFT_REG <= 'x;
		lvb_ld__0_reg_NO_SHIFT_REG <= 'x;
		lvb_cmp_0_reg_NO_SHIFT_REG <= 'x;
		lvb_var__u8_0_reg_NO_SHIFT_REG <= 'x;
		lvb_indvars_iv29_0_reg_NO_SHIFT_REG <= 'x;
		lvb_sub25_add24_0_reg_NO_SHIFT_REG <= 'x;
		lvb_arrayidx43_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_indvars_iv_next_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe1_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe2_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_idxprom_0_reg_NO_SHIFT_REG <= (rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[63:0] & 64'hFFFFFFFF);
			lvb_ld__0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[352:321];
			lvb_cmp_0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[64];
			lvb_var__u8_0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[353];
			lvb_indvars_iv29_0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[128:65];
			lvb_sub25_add24_0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[256:225];
			lvb_arrayidx43_0_reg_NO_SHIFT_REG <= (rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[320:257] & 64'hFFFFFFFFFFFFFFFC);
			lvb_bb3_indvars_iv_next_0_reg_NO_SHIFT_REG <= rnode_397to399_bb3_indvars_iv_next_0_NO_SHIFT_REG;
			lvb_bb3_c0_exe1_0_reg_NO_SHIFT_REG <= local_bb3_c0_exe1;
			lvb_bb3_c0_exe2_0_reg_NO_SHIFT_REG <= local_bb3_c0_exe2;
			lvb_input_global_id_0_0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[160:129];
			lvb_input_global_id_1_0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[192:161];
			lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG <= rcnode_398to399_rc0_idxprom_0_NO_SHIFT_REG[224:193];
			branch_compare_result_NO_SHIFT_REG <= local_bb3_var__u11;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_4
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_r,
		input [31:0] 		input_wii_sub25,
		input [31:0] 		input_wii_sub29,
		input [31:0] 		input_wii_mul50,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u95,
		input 		valid_in,
		output 		stall_out,
		input [63:0] 		input_idxprom,
		input [31:0] 		input_ld_,
		input 		input_cmp,
		input 		input_var__u96,
		input [63:0] 		input_indvars_iv29,
		input [31:0] 		input_c0_exe1,
		input [31:0] 		input_c0_exe2,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		input [31:0] 		input_acl_hw_wg_id,
		output 		valid_out_0,
		input 		stall_in_0,
		output [63:0] 		lvb_idxprom_0,
		output [31:0] 		lvb_ld__0,
		output 		lvb_cmp_0,
		output 		lvb_var__u96_0,
		output [31:0] 		lvb_c0_exe1_0,
		output [31:0] 		lvb_c0_exe2_0,
		output [63:0] 		lvb_bb4_indvars_iv_next30_0,
		output [31:0] 		lvb_input_global_id_0_0,
		output [31:0] 		lvb_input_global_id_1_0,
		output [31:0] 		lvb_input_acl_hw_wg_id_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [63:0] 		lvb_idxprom_1,
		output [31:0] 		lvb_ld__1,
		output 		lvb_cmp_1,
		output 		lvb_var__u96_1,
		output [31:0] 		lvb_c0_exe1_1,
		output [31:0] 		lvb_c0_exe2_1,
		output [63:0] 		lvb_bb4_indvars_iv_next30_1,
		output [31:0] 		lvb_input_global_id_0_1,
		output [31:0] 		lvb_input_global_id_1_1,
		output [31:0] 		lvb_input_acl_hw_wg_id_1,
		input [31:0] 		workgroup_size,
		input 		start
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_idxprom_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_ld__staging_reg_NO_SHIFT_REG;
 reg input_cmp_staging_reg_NO_SHIFT_REG;
 reg input_var__u96_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv29_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe2_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_idxprom_NO_SHIFT_REG;
 reg [31:0] local_lvm_ld__NO_SHIFT_REG;
 reg local_lvm_cmp_NO_SHIFT_REG;
 reg local_lvm_var__u96_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv29_NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe1_NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe2_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_idxprom_staging_reg_NO_SHIFT_REG <= 'x;
		input_ld__staging_reg_NO_SHIFT_REG <= 'x;
		input_cmp_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u96_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv29_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe2_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_idxprom_staging_reg_NO_SHIFT_REG <= input_idxprom;
				input_ld__staging_reg_NO_SHIFT_REG <= input_ld_;
				input_cmp_staging_reg_NO_SHIFT_REG <= input_cmp;
				input_var__u96_staging_reg_NO_SHIFT_REG <= input_var__u96;
				input_indvars_iv29_staging_reg_NO_SHIFT_REG <= input_indvars_iv29;
				input_c0_exe1_staging_reg_NO_SHIFT_REG <= input_c0_exe1;
				input_c0_exe2_staging_reg_NO_SHIFT_REG <= input_c0_exe2;
				input_global_id_0_staging_reg_NO_SHIFT_REG <= input_global_id_0;
				input_global_id_1_staging_reg_NO_SHIFT_REG <= input_global_id_1;
				input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_staging_reg_NO_SHIFT_REG;
					local_lvm_ld__NO_SHIFT_REG <= input_ld__staging_reg_NO_SHIFT_REG;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u96_NO_SHIFT_REG <= input_var__u96_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1_NO_SHIFT_REG <= input_c0_exe1_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe2_NO_SHIFT_REG <= input_c0_exe2_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom;
					local_lvm_ld__NO_SHIFT_REG <= input_ld_;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp;
					local_lvm_var__u96_NO_SHIFT_REG <= input_var__u96;
					local_lvm_indvars_iv29_NO_SHIFT_REG <= input_indvars_iv29;
					local_lvm_c0_exe1_NO_SHIFT_REG <= input_c0_exe1;
					local_lvm_c0_exe2_NO_SHIFT_REG <= input_c0_exe2;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_indvars_iv_next30_stall_local;
wire [63:0] local_bb4_indvars_iv_next30;
wire [257:0] rci_rcnode_1to3_rc1_idxprom_0_reg_1;

assign local_bb4_indvars_iv_next30 = (local_lvm_indvars_iv29_NO_SHIFT_REG + 64'h1);
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[63:0] = (local_lvm_idxprom_NO_SHIFT_REG & 64'hFFFFFFFF);
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[95:64] = local_lvm_ld__NO_SHIFT_REG;
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[96] = local_lvm_cmp_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[97] = local_lvm_var__u96_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[129:98] = local_lvm_c0_exe1_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[161:130] = local_lvm_c0_exe2_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[193:162] = local_lvm_input_global_id_0_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[225:194] = local_lvm_input_global_id_1_NO_SHIFT_REG;
assign rci_rcnode_1to3_rc1_idxprom_0_reg_1[257:226] = local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rcnode_1to3_rc1_idxprom_0_valid_out_0_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_stall_in_0_NO_SHIFT_REG;
 logic [257:0] rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_valid_out_1_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_stall_in_1_NO_SHIFT_REG;
 logic [257:0] rcnode_1to3_rc1_idxprom_1_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [257:0] rcnode_1to3_rc1_idxprom_0_reg_3_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_valid_out_0_reg_3_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_stall_in_0_reg_3_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_stall_out_reg_3_IP_NO_SHIFT_REG;
 logic rcnode_1to3_rc1_idxprom_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rcnode_1to3_rc1_idxprom_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to3_rc1_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to3_rc1_idxprom_0_stall_in_0_reg_3_NO_SHIFT_REG),
	.valid_out(rcnode_1to3_rc1_idxprom_0_valid_out_0_reg_3_NO_SHIFT_REG),
	.stall_out(rcnode_1to3_rc1_idxprom_0_stall_out_reg_3_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to3_rc1_idxprom_0_reg_1),
	.data_out(rcnode_1to3_rc1_idxprom_0_reg_3_NO_SHIFT_REG)
);

defparam rcnode_1to3_rc1_idxprom_0_reg_3_fifo.DEPTH = 3;
defparam rcnode_1to3_rc1_idxprom_0_reg_3_fifo.DATA_WIDTH = 258;
defparam rcnode_1to3_rc1_idxprom_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to3_rc1_idxprom_0_reg_3_fifo.IMPL = "ll_reg";

assign rcnode_1to3_rc1_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign rcnode_1to3_rc1_idxprom_0_stall_out_reg_3_NO_SHIFT_REG = (~(rcnode_1to3_rc1_idxprom_0_reg_3_inputs_ready_NO_SHIFT_REG) | rcnode_1to3_rc1_idxprom_0_stall_out_reg_3_IP_NO_SHIFT_REG);
assign merge_node_stall_in_1 = rcnode_1to3_rc1_idxprom_0_stall_out_reg_3_NO_SHIFT_REG;
assign rcnode_1to3_rc1_idxprom_0_stall_in_0_reg_3_NO_SHIFT_REG = (rcnode_1to3_rc1_idxprom_0_stall_in_0_NO_SHIFT_REG | rcnode_1to3_rc1_idxprom_0_stall_in_1_NO_SHIFT_REG);
assign rcnode_1to3_rc1_idxprom_0_valid_out_0_NO_SHIFT_REG = rcnode_1to3_rc1_idxprom_0_valid_out_0_reg_3_NO_SHIFT_REG;
assign rcnode_1to3_rc1_idxprom_0_valid_out_1_NO_SHIFT_REG = rcnode_1to3_rc1_idxprom_0_valid_out_0_reg_3_NO_SHIFT_REG;
assign rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG = rcnode_1to3_rc1_idxprom_0_reg_3_NO_SHIFT_REG;
assign rcnode_1to3_rc1_idxprom_1_NO_SHIFT_REG = rcnode_1to3_rc1_idxprom_0_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_indvars_iv_next30_valid_out_1;
wire local_bb4_indvars_iv_next30_stall_in_1;
wire local_bb4_var__valid_out;
wire local_bb4_var__stall_in;
wire local_bb4_var__inputs_ready;
wire local_bb4_var__stall_local;
wire [31:0] local_bb4_var_;
 reg local_bb4_indvars_iv_next30_consumed_1_NO_SHIFT_REG;
 reg local_bb4_var__consumed_0_NO_SHIFT_REG;

assign local_bb4_var__inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb4_var_ = local_bb4_indvars_iv_next30[31:0];
assign local_bb4_var__stall_local = ((local_bb4_indvars_iv_next30_stall_in_1 & ~(local_bb4_indvars_iv_next30_consumed_1_NO_SHIFT_REG)) | (local_bb4_var__stall_in & ~(local_bb4_var__consumed_0_NO_SHIFT_REG)));
assign local_bb4_indvars_iv_next30_valid_out_1 = (local_bb4_var__inputs_ready & ~(local_bb4_indvars_iv_next30_consumed_1_NO_SHIFT_REG));
assign local_bb4_var__valid_out = (local_bb4_var__inputs_ready & ~(local_bb4_var__consumed_0_NO_SHIFT_REG));
assign merge_node_stall_in_0 = (|local_bb4_var__stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_indvars_iv_next30_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_var__consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb4_indvars_iv_next30_consumed_1_NO_SHIFT_REG <= (local_bb4_var__inputs_ready & (local_bb4_indvars_iv_next30_consumed_1_NO_SHIFT_REG | ~(local_bb4_indvars_iv_next30_stall_in_1)) & local_bb4_var__stall_local);
		local_bb4_var__consumed_0_NO_SHIFT_REG <= (local_bb4_var__inputs_ready & (local_bb4_var__consumed_0_NO_SHIFT_REG | ~(local_bb4_var__stall_in)) & local_bb4_var__stall_local);
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb4_indvars_iv_next30_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb4_indvars_iv_next30_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_1to3_bb4_indvars_iv_next30_0_NO_SHIFT_REG;
 logic rnode_1to3_bb4_indvars_iv_next30_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to3_bb4_indvars_iv_next30_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb4_indvars_iv_next30_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb4_indvars_iv_next30_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb4_indvars_iv_next30_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb4_indvars_iv_next30_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb4_indvars_iv_next30_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb4_indvars_iv_next30_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb4_indvars_iv_next30_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb4_indvars_iv_next30_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb4_indvars_iv_next30),
	.data_out(rnode_1to3_bb4_indvars_iv_next30_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb4_indvars_iv_next30_0_reg_3_fifo.DEPTH = 3;
defparam rnode_1to3_bb4_indvars_iv_next30_0_reg_3_fifo.DATA_WIDTH = 64;
defparam rnode_1to3_bb4_indvars_iv_next30_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to3_bb4_indvars_iv_next30_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_1to3_bb4_indvars_iv_next30_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb4_indvars_iv_next30_valid_out_1;
assign local_bb4_indvars_iv_next30_stall_in_1 = rnode_1to3_bb4_indvars_iv_next30_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb4_indvars_iv_next30_0_NO_SHIFT_REG = rnode_1to3_bb4_indvars_iv_next30_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb4_indvars_iv_next30_0_stall_in_reg_3_NO_SHIFT_REG = rnode_1to3_bb4_indvars_iv_next30_0_stall_in_NO_SHIFT_REG;
assign rnode_1to3_bb4_indvars_iv_next30_0_valid_out_NO_SHIFT_REG = rnode_1to3_bb4_indvars_iv_next30_0_valid_out_reg_3_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_var__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_var__0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_var__0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_var__0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_var__0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_var__0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_var__0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_var__0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_var__0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_var__0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_var__0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_var__0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_var_),
	.data_out(rnode_1to2_bb4_var__0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_var__0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_var__0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_var__0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_var__0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb4_var__0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb4_var__valid_out;
assign local_bb4_var__stall_in = rnode_1to2_bb4_var__0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_var__0_NO_SHIFT_REG = rnode_1to2_bb4_var__0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_var__0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb4_var__0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb4_var__0_valid_out_NO_SHIFT_REG = rnode_1to2_bb4_var__0_valid_out_reg_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp16_valid_out;
wire local_bb4_cmp16_stall_in;
wire local_bb4_cmp16_inputs_ready;
wire local_bb4_cmp16_stall_local;
wire local_bb4_cmp16;

assign local_bb4_cmp16_inputs_ready = rnode_1to2_bb4_var__0_valid_out_NO_SHIFT_REG;
assign local_bb4_cmp16 = ($signed(rnode_1to2_bb4_var__0_NO_SHIFT_REG) > $signed(input_r));
assign local_bb4_cmp16_valid_out = local_bb4_cmp16_inputs_ready;
assign local_bb4_cmp16_stall_local = local_bb4_cmp16_stall_in;
assign rnode_1to2_bb4_var__0_stall_in_NO_SHIFT_REG = (|local_bb4_cmp16_stall_local);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb4_cmp16_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb4_cmp16_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb4_cmp16_0_NO_SHIFT_REG;
 logic rnode_2to3_bb4_cmp16_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb4_cmp16_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb4_cmp16_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb4_cmp16_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb4_cmp16_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb4_cmp16_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb4_cmp16_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb4_cmp16_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb4_cmp16_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb4_cmp16_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb4_cmp16),
	.data_out(rnode_2to3_bb4_cmp16_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb4_cmp16_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb4_cmp16_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb4_cmp16_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb4_cmp16_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_2to3_bb4_cmp16_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb4_cmp16_valid_out;
assign local_bb4_cmp16_stall_in = rnode_2to3_bb4_cmp16_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb4_cmp16_0_NO_SHIFT_REG = rnode_2to3_bb4_cmp16_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb4_cmp16_0_stall_in_reg_3_NO_SHIFT_REG = rnode_2to3_bb4_cmp16_0_stall_in_NO_SHIFT_REG;
assign rnode_2to3_bb4_cmp16_0_valid_out_NO_SHIFT_REG = rnode_2to3_bb4_cmp16_0_valid_out_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u97_valid_out;
wire local_bb4_var__u97_stall_in;
wire local_bb4_var__u97_inputs_ready;
wire local_bb4_var__u97_stall_local;
wire local_bb4_var__u97;

assign local_bb4_var__u97_inputs_ready = (rnode_2to3_bb4_cmp16_0_valid_out_NO_SHIFT_REG & rcnode_1to3_rc1_idxprom_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_var__u97 = (rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[97] | rnode_2to3_bb4_cmp16_0_NO_SHIFT_REG);
assign local_bb4_var__u97_valid_out = local_bb4_var__u97_inputs_ready;
assign local_bb4_var__u97_stall_local = local_bb4_var__u97_stall_in;
assign rnode_2to3_bb4_cmp16_0_stall_in_NO_SHIFT_REG = (local_bb4_var__u97_stall_local | ~(local_bb4_var__u97_inputs_ready));
assign rcnode_1to3_rc1_idxprom_0_stall_in_1_NO_SHIFT_REG = (local_bb4_var__u97_stall_local | ~(local_bb4_var__u97_inputs_ready));

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_idxprom_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_ld__0_reg_NO_SHIFT_REG;
 reg lvb_cmp_0_reg_NO_SHIFT_REG;
 reg lvb_var__u96_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_c0_exe1_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_c0_exe2_0_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb4_indvars_iv_next30_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb4_var__u97_valid_out & rnode_1to3_bb4_indvars_iv_next30_0_valid_out_NO_SHIFT_REG & rcnode_1to3_rc1_idxprom_0_valid_out_0_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb4_var__u97_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to3_bb4_indvars_iv_next30_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_1to3_rc1_idxprom_0_stall_in_0_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_idxprom_0 = lvb_idxprom_0_reg_NO_SHIFT_REG;
assign lvb_idxprom_1 = lvb_idxprom_0_reg_NO_SHIFT_REG;
assign lvb_ld__0 = lvb_ld__0_reg_NO_SHIFT_REG;
assign lvb_ld__1 = lvb_ld__0_reg_NO_SHIFT_REG;
assign lvb_cmp_0 = lvb_cmp_0_reg_NO_SHIFT_REG;
assign lvb_cmp_1 = lvb_cmp_0_reg_NO_SHIFT_REG;
assign lvb_var__u96_0 = lvb_var__u96_0_reg_NO_SHIFT_REG;
assign lvb_var__u96_1 = lvb_var__u96_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1_0 = lvb_c0_exe1_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1_1 = lvb_c0_exe1_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe2_0 = lvb_c0_exe2_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe2_1 = lvb_c0_exe2_0_reg_NO_SHIFT_REG;
assign lvb_bb4_indvars_iv_next30_0 = lvb_bb4_indvars_iv_next30_0_reg_NO_SHIFT_REG;
assign lvb_bb4_indvars_iv_next30_1 = lvb_bb4_indvars_iv_next30_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0_0 = lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0_1 = lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1_0 = lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1_1 = lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
assign lvb_input_acl_hw_wg_id_0 = lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG;
assign lvb_input_acl_hw_wg_id_1 = lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_idxprom_0_reg_NO_SHIFT_REG <= 'x;
		lvb_ld__0_reg_NO_SHIFT_REG <= 'x;
		lvb_cmp_0_reg_NO_SHIFT_REG <= 'x;
		lvb_var__u96_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe1_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe2_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_indvars_iv_next30_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_idxprom_0_reg_NO_SHIFT_REG <= (rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[63:0] & 64'hFFFFFFFF);
			lvb_ld__0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[95:64];
			lvb_cmp_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[96];
			lvb_var__u96_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[97];
			lvb_c0_exe1_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[129:98];
			lvb_c0_exe2_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[161:130];
			lvb_bb4_indvars_iv_next30_0_reg_NO_SHIFT_REG <= rnode_1to3_bb4_indvars_iv_next30_0_NO_SHIFT_REG;
			lvb_input_global_id_0_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[193:162];
			lvb_input_global_id_1_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[225:194];
			lvb_input_acl_hw_wg_id_0_reg_NO_SHIFT_REG <= rcnode_1to3_rc1_idxprom_0_NO_SHIFT_REG[257:226];
			branch_compare_result_NO_SHIFT_REG <= local_bb4_var__u97;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_5
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_out,
		input 		valid_in,
		output 		stall_out,
		input [63:0] 		input_idxprom,
		input 		input_cmp,
		input 		input_var_,
		input [31:0] 		input_c0_exe1,
		input [31:0] 		input_c0_exe2,
		input [31:0] 		input_acl_hw_wg_id,
		output 		valid_out,
		input 		stall_in,
		output [31:0] 		lvb_input_acl_hw_wg_id,
		input [31:0] 		workgroup_size,
		input 		start,
		input [511:0] 		avm_local_bb5_st_c0_exe112_readdata,
		input 		avm_local_bb5_st_c0_exe112_readdatavalid,
		input 		avm_local_bb5_st_c0_exe112_waitrequest,
		output [32:0] 		avm_local_bb5_st_c0_exe112_address,
		output 		avm_local_bb5_st_c0_exe112_read,
		output 		avm_local_bb5_st_c0_exe112_write,
		input 		avm_local_bb5_st_c0_exe112_writeack,
		output [511:0] 		avm_local_bb5_st_c0_exe112_writedata,
		output [63:0] 		avm_local_bb5_st_c0_exe112_byteenable,
		output [4:0] 		avm_local_bb5_st_c0_exe112_burstcount,
		output 		local_bb5_st_c0_exe112_active,
		input 		clock2x
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_idxprom_staging_reg_NO_SHIFT_REG;
 reg input_cmp_staging_reg_NO_SHIFT_REG;
 reg input_var__staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe2_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_idxprom_NO_SHIFT_REG;
 reg local_lvm_cmp_NO_SHIFT_REG;
 reg local_lvm_var__NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe1_NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe2_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_idxprom_staging_reg_NO_SHIFT_REG <= 'x;
		input_cmp_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe2_staging_reg_NO_SHIFT_REG <= 'x;
		input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_idxprom_staging_reg_NO_SHIFT_REG <= input_idxprom;
				input_cmp_staging_reg_NO_SHIFT_REG <= input_cmp;
				input_var__staging_reg_NO_SHIFT_REG <= input_var_;
				input_c0_exe1_staging_reg_NO_SHIFT_REG <= input_c0_exe1;
				input_c0_exe2_staging_reg_NO_SHIFT_REG <= input_c0_exe2;
				input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG <= input_acl_hw_wg_id;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom_staging_reg_NO_SHIFT_REG;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp_staging_reg_NO_SHIFT_REG;
					local_lvm_var__NO_SHIFT_REG <= input_var__staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1_NO_SHIFT_REG <= input_c0_exe1_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe2_NO_SHIFT_REG <= input_c0_exe2_staging_reg_NO_SHIFT_REG;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_idxprom_NO_SHIFT_REG <= input_idxprom;
					local_lvm_cmp_NO_SHIFT_REG <= input_cmp;
					local_lvm_var__NO_SHIFT_REG <= input_var_;
					local_lvm_c0_exe1_NO_SHIFT_REG <= input_c0_exe1;
					local_lvm_c0_exe2_NO_SHIFT_REG <= input_c0_exe2;
					local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG <= input_acl_hw_wg_id;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5_c0_eni11_stall_local;
wire [127:0] local_bb5_c0_eni11;

assign local_bb5_c0_eni11[7:0] = 8'bx;
assign local_bb5_c0_eni11[8] = local_lvm_var__NO_SHIFT_REG;
assign local_bb5_c0_eni11[127:9] = 119'bx;

// Register node:
//  * latency = 23
//  * capacity = 23
 logic rnode_1to24_input_acl_hw_wg_id_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to24_input_acl_hw_wg_id_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to24_input_acl_hw_wg_id_0_NO_SHIFT_REG;
 logic rnode_1to24_input_acl_hw_wg_id_0_reg_24_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to24_input_acl_hw_wg_id_0_reg_24_NO_SHIFT_REG;
 logic rnode_1to24_input_acl_hw_wg_id_0_valid_out_reg_24_NO_SHIFT_REG;
 logic rnode_1to24_input_acl_hw_wg_id_0_stall_in_reg_24_NO_SHIFT_REG;
 logic rnode_1to24_input_acl_hw_wg_id_0_stall_out_reg_24_NO_SHIFT_REG;
wire [127:0] rci_rcnode_1to19_rc5_input_out_0_reg_1;

acl_data_fifo rnode_1to24_input_acl_hw_wg_id_0_reg_24_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to24_input_acl_hw_wg_id_0_reg_24_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to24_input_acl_hw_wg_id_0_stall_in_reg_24_NO_SHIFT_REG),
	.valid_out(rnode_1to24_input_acl_hw_wg_id_0_valid_out_reg_24_NO_SHIFT_REG),
	.stall_out(rnode_1to24_input_acl_hw_wg_id_0_stall_out_reg_24_NO_SHIFT_REG),
	.data_in(local_lvm_input_acl_hw_wg_id_NO_SHIFT_REG),
	.data_out(rnode_1to24_input_acl_hw_wg_id_0_reg_24_NO_SHIFT_REG)
);

defparam rnode_1to24_input_acl_hw_wg_id_0_reg_24_fifo.DEPTH = 24;
defparam rnode_1to24_input_acl_hw_wg_id_0_reg_24_fifo.DATA_WIDTH = 32;
defparam rnode_1to24_input_acl_hw_wg_id_0_reg_24_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to24_input_acl_hw_wg_id_0_reg_24_fifo.IMPL = "ram";

assign rnode_1to24_input_acl_hw_wg_id_0_reg_24_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_4_NO_SHIFT_REG;
assign merge_node_stall_in_4 = rnode_1to24_input_acl_hw_wg_id_0_stall_out_reg_24_NO_SHIFT_REG;
assign rnode_1to24_input_acl_hw_wg_id_0_NO_SHIFT_REG = rnode_1to24_input_acl_hw_wg_id_0_reg_24_NO_SHIFT_REG;
assign rnode_1to24_input_acl_hw_wg_id_0_stall_in_reg_24_NO_SHIFT_REG = rnode_1to24_input_acl_hw_wg_id_0_stall_in_NO_SHIFT_REG;
assign rnode_1to24_input_acl_hw_wg_id_0_valid_out_NO_SHIFT_REG = rnode_1to24_input_acl_hw_wg_id_0_valid_out_reg_24_NO_SHIFT_REG;
assign rci_rcnode_1to19_rc5_input_out_0_reg_1[63:0] = (input_out & 64'hFFFFFFFFFFFFFC00);
assign rci_rcnode_1to19_rc5_input_out_0_reg_1[127:64] = (local_lvm_idxprom_NO_SHIFT_REG & 64'hFFFFFFFF);

// Register node:
//  * latency = 18
//  * capacity = 18
 logic rcnode_1to19_rc5_input_out_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to19_rc5_input_out_0_stall_in_NO_SHIFT_REG;
 logic [127:0] rcnode_1to19_rc5_input_out_0_NO_SHIFT_REG;
 logic rcnode_1to19_rc5_input_out_0_reg_19_inputs_ready_NO_SHIFT_REG;
 logic [127:0] rcnode_1to19_rc5_input_out_0_reg_19_NO_SHIFT_REG;
 logic rcnode_1to19_rc5_input_out_0_valid_out_reg_19_NO_SHIFT_REG;
 logic rcnode_1to19_rc5_input_out_0_stall_in_reg_19_NO_SHIFT_REG;
 logic rcnode_1to19_rc5_input_out_0_stall_out_reg_19_IP_NO_SHIFT_REG;
 logic rcnode_1to19_rc5_input_out_0_stall_out_reg_19_NO_SHIFT_REG;

acl_data_fifo rcnode_1to19_rc5_input_out_0_reg_19_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to19_rc5_input_out_0_reg_19_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to19_rc5_input_out_0_stall_in_reg_19_NO_SHIFT_REG),
	.valid_out(rcnode_1to19_rc5_input_out_0_valid_out_reg_19_NO_SHIFT_REG),
	.stall_out(rcnode_1to19_rc5_input_out_0_stall_out_reg_19_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to19_rc5_input_out_0_reg_1),
	.data_out(rcnode_1to19_rc5_input_out_0_reg_19_NO_SHIFT_REG)
);

defparam rcnode_1to19_rc5_input_out_0_reg_19_fifo.DEPTH = 19;
defparam rcnode_1to19_rc5_input_out_0_reg_19_fifo.DATA_WIDTH = 128;
defparam rcnode_1to19_rc5_input_out_0_reg_19_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to19_rc5_input_out_0_reg_19_fifo.IMPL = "ram";

assign rcnode_1to19_rc5_input_out_0_reg_19_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign rcnode_1to19_rc5_input_out_0_stall_out_reg_19_NO_SHIFT_REG = (~(rcnode_1to19_rc5_input_out_0_reg_19_inputs_ready_NO_SHIFT_REG) | rcnode_1to19_rc5_input_out_0_stall_out_reg_19_IP_NO_SHIFT_REG);
assign merge_node_stall_in_5 = rcnode_1to19_rc5_input_out_0_stall_out_reg_19_NO_SHIFT_REG;
assign rcnode_1to19_rc5_input_out_0_NO_SHIFT_REG = rcnode_1to19_rc5_input_out_0_reg_19_NO_SHIFT_REG;
assign rcnode_1to19_rc5_input_out_0_stall_in_reg_19_NO_SHIFT_REG = rcnode_1to19_rc5_input_out_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to19_rc5_input_out_0_valid_out_NO_SHIFT_REG = rcnode_1to19_rc5_input_out_0_valid_out_reg_19_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb5_c0_eni22_stall_local;
wire [127:0] local_bb5_c0_eni22;

assign local_bb5_c0_eni22[31:0] = local_bb5_c0_eni11[31:0];
assign local_bb5_c0_eni22[63:32] = local_lvm_c0_exe2_NO_SHIFT_REG;
assign local_bb5_c0_eni22[127:64] = local_bb5_c0_eni11[127:64];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_24to25_input_acl_hw_wg_id_0_valid_out_NO_SHIFT_REG;
 logic rnode_24to25_input_acl_hw_wg_id_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_24to25_input_acl_hw_wg_id_0_NO_SHIFT_REG;
 logic rnode_24to25_input_acl_hw_wg_id_0_reg_25_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_24to25_input_acl_hw_wg_id_0_reg_25_NO_SHIFT_REG;
 logic rnode_24to25_input_acl_hw_wg_id_0_valid_out_reg_25_NO_SHIFT_REG;
 logic rnode_24to25_input_acl_hw_wg_id_0_stall_in_reg_25_NO_SHIFT_REG;
 logic rnode_24to25_input_acl_hw_wg_id_0_stall_out_reg_25_NO_SHIFT_REG;
wire [127:0] rci_rcnode_19to20_rc0_input_out_0_reg_19;

acl_data_fifo rnode_24to25_input_acl_hw_wg_id_0_reg_25_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_24to25_input_acl_hw_wg_id_0_reg_25_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_24to25_input_acl_hw_wg_id_0_stall_in_reg_25_NO_SHIFT_REG),
	.valid_out(rnode_24to25_input_acl_hw_wg_id_0_valid_out_reg_25_NO_SHIFT_REG),
	.stall_out(rnode_24to25_input_acl_hw_wg_id_0_stall_out_reg_25_NO_SHIFT_REG),
	.data_in(rnode_1to24_input_acl_hw_wg_id_0_NO_SHIFT_REG),
	.data_out(rnode_24to25_input_acl_hw_wg_id_0_reg_25_NO_SHIFT_REG)
);

defparam rnode_24to25_input_acl_hw_wg_id_0_reg_25_fifo.DEPTH = 1;
defparam rnode_24to25_input_acl_hw_wg_id_0_reg_25_fifo.DATA_WIDTH = 32;
defparam rnode_24to25_input_acl_hw_wg_id_0_reg_25_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_24to25_input_acl_hw_wg_id_0_reg_25_fifo.IMPL = "ll_reg";

assign rnode_24to25_input_acl_hw_wg_id_0_reg_25_inputs_ready_NO_SHIFT_REG = rnode_1to24_input_acl_hw_wg_id_0_valid_out_NO_SHIFT_REG;
assign rnode_1to24_input_acl_hw_wg_id_0_stall_in_NO_SHIFT_REG = rnode_24to25_input_acl_hw_wg_id_0_stall_out_reg_25_NO_SHIFT_REG;
assign rnode_24to25_input_acl_hw_wg_id_0_NO_SHIFT_REG = rnode_24to25_input_acl_hw_wg_id_0_reg_25_NO_SHIFT_REG;
assign rnode_24to25_input_acl_hw_wg_id_0_stall_in_reg_25_NO_SHIFT_REG = rnode_24to25_input_acl_hw_wg_id_0_stall_in_NO_SHIFT_REG;
assign rnode_24to25_input_acl_hw_wg_id_0_valid_out_NO_SHIFT_REG = rnode_24to25_input_acl_hw_wg_id_0_valid_out_reg_25_NO_SHIFT_REG;
assign rci_rcnode_19to20_rc0_input_out_0_reg_19[63:0] = (input_out & 64'hFFFFFFFFFFFFFC00);
assign rci_rcnode_19to20_rc0_input_out_0_reg_19[127:64] = (rcnode_1to19_rc5_input_out_0_NO_SHIFT_REG[127:64] & 64'hFFFFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_19to20_rc0_input_out_0_valid_out_NO_SHIFT_REG;
 logic rcnode_19to20_rc0_input_out_0_stall_in_NO_SHIFT_REG;
 logic [127:0] rcnode_19to20_rc0_input_out_0_NO_SHIFT_REG;
 logic rcnode_19to20_rc0_input_out_0_reg_20_inputs_ready_NO_SHIFT_REG;
 logic [127:0] rcnode_19to20_rc0_input_out_0_reg_20_NO_SHIFT_REG;
 logic rcnode_19to20_rc0_input_out_0_valid_out_reg_20_NO_SHIFT_REG;
 logic rcnode_19to20_rc0_input_out_0_stall_in_reg_20_NO_SHIFT_REG;
 logic rcnode_19to20_rc0_input_out_0_stall_out_reg_20_IP_NO_SHIFT_REG;
 logic rcnode_19to20_rc0_input_out_0_stall_out_reg_20_NO_SHIFT_REG;

acl_data_fifo rcnode_19to20_rc0_input_out_0_reg_20_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_19to20_rc0_input_out_0_reg_20_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_19to20_rc0_input_out_0_stall_in_reg_20_NO_SHIFT_REG),
	.valid_out(rcnode_19to20_rc0_input_out_0_valid_out_reg_20_NO_SHIFT_REG),
	.stall_out(rcnode_19to20_rc0_input_out_0_stall_out_reg_20_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_19to20_rc0_input_out_0_reg_19),
	.data_out(rcnode_19to20_rc0_input_out_0_reg_20_NO_SHIFT_REG)
);

defparam rcnode_19to20_rc0_input_out_0_reg_20_fifo.DEPTH = 1;
defparam rcnode_19to20_rc0_input_out_0_reg_20_fifo.DATA_WIDTH = 128;
defparam rcnode_19to20_rc0_input_out_0_reg_20_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_19to20_rc0_input_out_0_reg_20_fifo.IMPL = "ll_reg";

assign rcnode_19to20_rc0_input_out_0_reg_20_inputs_ready_NO_SHIFT_REG = rcnode_1to19_rc5_input_out_0_valid_out_NO_SHIFT_REG;
assign rcnode_19to20_rc0_input_out_0_stall_out_reg_20_NO_SHIFT_REG = (~(rcnode_19to20_rc0_input_out_0_reg_20_inputs_ready_NO_SHIFT_REG) | rcnode_19to20_rc0_input_out_0_stall_out_reg_20_IP_NO_SHIFT_REG);
assign rcnode_1to19_rc5_input_out_0_stall_in_NO_SHIFT_REG = rcnode_19to20_rc0_input_out_0_stall_out_reg_20_NO_SHIFT_REG;
assign rcnode_19to20_rc0_input_out_0_NO_SHIFT_REG = rcnode_19to20_rc0_input_out_0_reg_20_NO_SHIFT_REG;
assign rcnode_19to20_rc0_input_out_0_stall_in_reg_20_NO_SHIFT_REG = rcnode_19to20_rc0_input_out_0_stall_in_NO_SHIFT_REG;
assign rcnode_19to20_rc0_input_out_0_valid_out_NO_SHIFT_REG = rcnode_19to20_rc0_input_out_0_valid_out_reg_20_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb5_c0_eni33_stall_local;
wire [127:0] local_bb5_c0_eni33;

assign local_bb5_c0_eni33[63:0] = local_bb5_c0_eni22[63:0];
assign local_bb5_c0_eni33[95:64] = local_lvm_c0_exe1_NO_SHIFT_REG;
assign local_bb5_c0_eni33[127:96] = local_bb5_c0_eni22[127:96];

// This section implements an unregistered operation.
// 
wire local_bb5_arrayidx15_valid_out;
wire local_bb5_arrayidx15_stall_in;
wire local_bb5_arrayidx15_inputs_ready;
wire local_bb5_arrayidx15_stall_local;
wire [63:0] local_bb5_arrayidx15;

assign local_bb5_arrayidx15_inputs_ready = rcnode_19to20_rc0_input_out_0_valid_out_NO_SHIFT_REG;
assign local_bb5_arrayidx15 = ((input_out & 64'hFFFFFFFFFFFFFC00) + ((rcnode_19to20_rc0_input_out_0_NO_SHIFT_REG[127:64] & 64'hFFFFFFFF) << 6'h2));
assign local_bb5_arrayidx15_valid_out = local_bb5_arrayidx15_inputs_ready;
assign local_bb5_arrayidx15_stall_local = local_bb5_arrayidx15_stall_in;
assign rcnode_19to20_rc0_input_out_0_stall_in_NO_SHIFT_REG = (|local_bb5_arrayidx15_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb5_c0_eni44_valid_out;
wire local_bb5_c0_eni44_stall_in;
wire local_bb5_c0_eni44_inputs_ready;
wire local_bb5_c0_eni44_stall_local;
wire [127:0] local_bb5_c0_eni44;

assign local_bb5_c0_eni44_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_3_NO_SHIFT_REG);
assign local_bb5_c0_eni44[95:0] = local_bb5_c0_eni33[95:0];
assign local_bb5_c0_eni44[96] = local_lvm_cmp_NO_SHIFT_REG;
assign local_bb5_c0_eni44[127:97] = local_bb5_c0_eni33[127:97];
assign local_bb5_c0_eni44_valid_out = local_bb5_c0_eni44_inputs_ready;
assign local_bb5_c0_eni44_stall_local = local_bb5_c0_eni44_stall_in;
assign merge_node_stall_in_0 = (local_bb5_c0_eni44_stall_local | ~(local_bb5_c0_eni44_inputs_ready));
assign merge_node_stall_in_1 = (local_bb5_c0_eni44_stall_local | ~(local_bb5_c0_eni44_inputs_ready));
assign merge_node_stall_in_2 = (local_bb5_c0_eni44_stall_local | ~(local_bb5_c0_eni44_inputs_ready));
assign merge_node_stall_in_3 = (local_bb5_c0_eni44_stall_local | ~(local_bb5_c0_eni44_inputs_ready));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_20to21_bb5_arrayidx15_0_valid_out_NO_SHIFT_REG;
 logic rnode_20to21_bb5_arrayidx15_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb5_arrayidx15_0_NO_SHIFT_REG;
 logic rnode_20to21_bb5_arrayidx15_0_reg_21_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb5_arrayidx15_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb5_arrayidx15_0_valid_out_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb5_arrayidx15_0_stall_in_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb5_arrayidx15_0_stall_out_reg_21_NO_SHIFT_REG;

acl_data_fifo rnode_20to21_bb5_arrayidx15_0_reg_21_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_20to21_bb5_arrayidx15_0_reg_21_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_20to21_bb5_arrayidx15_0_stall_in_reg_21_NO_SHIFT_REG),
	.valid_out(rnode_20to21_bb5_arrayidx15_0_valid_out_reg_21_NO_SHIFT_REG),
	.stall_out(rnode_20to21_bb5_arrayidx15_0_stall_out_reg_21_NO_SHIFT_REG),
	.data_in((local_bb5_arrayidx15 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_20to21_bb5_arrayidx15_0_reg_21_NO_SHIFT_REG)
);

defparam rnode_20to21_bb5_arrayidx15_0_reg_21_fifo.DEPTH = 2;
defparam rnode_20to21_bb5_arrayidx15_0_reg_21_fifo.DATA_WIDTH = 64;
defparam rnode_20to21_bb5_arrayidx15_0_reg_21_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_20to21_bb5_arrayidx15_0_reg_21_fifo.IMPL = "ll_reg";

assign rnode_20to21_bb5_arrayidx15_0_reg_21_inputs_ready_NO_SHIFT_REG = local_bb5_arrayidx15_valid_out;
assign local_bb5_arrayidx15_stall_in = rnode_20to21_bb5_arrayidx15_0_stall_out_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb5_arrayidx15_0_NO_SHIFT_REG = rnode_20to21_bb5_arrayidx15_0_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb5_arrayidx15_0_stall_in_reg_21_NO_SHIFT_REG = rnode_20to21_bb5_arrayidx15_0_stall_in_NO_SHIFT_REG;
assign rnode_20to21_bb5_arrayidx15_0_valid_out_NO_SHIFT_REG = rnode_20to21_bb5_arrayidx15_0_valid_out_reg_21_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb5_c0_enter5_c0_eni44_inputs_ready;
 reg local_bb5_c0_enter5_c0_eni44_valid_out_0_NO_SHIFT_REG;
wire local_bb5_c0_enter5_c0_eni44_stall_in_0;
 reg local_bb5_c0_enter5_c0_eni44_valid_out_1_NO_SHIFT_REG;
wire local_bb5_c0_enter5_c0_eni44_stall_in_1;
 reg local_bb5_c0_enter5_c0_eni44_valid_out_2_NO_SHIFT_REG;
wire local_bb5_c0_enter5_c0_eni44_stall_in_2;
 reg local_bb5_c0_enter5_c0_eni44_valid_out_3_NO_SHIFT_REG;
wire local_bb5_c0_enter5_c0_eni44_stall_in_3;
 reg local_bb5_c0_enter5_c0_eni44_valid_out_4_NO_SHIFT_REG;
wire local_bb5_c0_enter5_c0_eni44_stall_in_4;
wire local_bb5_c0_enter5_c0_eni44_output_regs_ready;
 reg [127:0] local_bb5_c0_enter5_c0_eni44_NO_SHIFT_REG;
wire local_bb5_c0_enter5_c0_eni44_input_accepted;
 reg local_bb5_c0_enter5_c0_eni44_valid_bit_NO_SHIFT_REG;
wire local_bb5_c0_exit11_c0_exi110_entry_stall;
wire local_bb5_c0_exit11_c0_exi110_output_regs_ready;
wire [15:0] local_bb5_c0_exit11_c0_exi110_valid_bits;
wire local_bb5_c0_exit11_c0_exi110_valid_in;
wire local_bb5_c0_exit11_c0_exi110_phases;
wire local_bb5_c0_enter5_c0_eni44_inc_pipelined_thread;
wire local_bb5_c0_enter5_c0_eni44_dec_pipelined_thread;
wire local_bb5_c0_enter5_c0_eni44_causedstall;

assign local_bb5_c0_enter5_c0_eni44_inputs_ready = local_bb5_c0_eni44_valid_out;
assign local_bb5_c0_enter5_c0_eni44_output_regs_ready = 1'b1;
assign local_bb5_c0_enter5_c0_eni44_input_accepted = (local_bb5_c0_enter5_c0_eni44_inputs_ready && !(local_bb5_c0_exit11_c0_exi110_entry_stall));
assign local_bb5_c0_enter5_c0_eni44_inc_pipelined_thread = 1'b1;
assign local_bb5_c0_enter5_c0_eni44_dec_pipelined_thread = ~(1'b0);
assign local_bb5_c0_eni44_stall_in = ((~(local_bb5_c0_enter5_c0_eni44_inputs_ready) | local_bb5_c0_exit11_c0_exi110_entry_stall) | ~(1'b1));
assign local_bb5_c0_enter5_c0_eni44_causedstall = (1'b1 && ((~(local_bb5_c0_enter5_c0_eni44_inputs_ready) | local_bb5_c0_exit11_c0_exi110_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_c0_enter5_c0_eni44_valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb5_c0_enter5_c0_eni44_valid_bit_NO_SHIFT_REG <= local_bb5_c0_enter5_c0_eni44_input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_c0_enter5_c0_eni44_NO_SHIFT_REG <= 'x;
		local_bb5_c0_enter5_c0_eni44_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb5_c0_enter5_c0_eni44_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb5_c0_enter5_c0_eni44_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb5_c0_enter5_c0_eni44_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb5_c0_enter5_c0_eni44_valid_out_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_c0_enter5_c0_eni44_output_regs_ready)
		begin
			local_bb5_c0_enter5_c0_eni44_NO_SHIFT_REG <= local_bb5_c0_eni44;
			local_bb5_c0_enter5_c0_eni44_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb5_c0_enter5_c0_eni44_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb5_c0_enter5_c0_eni44_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb5_c0_enter5_c0_eni44_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb5_c0_enter5_c0_eni44_valid_out_4_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb5_c0_enter5_c0_eni44_stall_in_0))
			begin
				local_bb5_c0_enter5_c0_eni44_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb5_c0_enter5_c0_eni44_stall_in_1))
			begin
				local_bb5_c0_enter5_c0_eni44_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb5_c0_enter5_c0_eni44_stall_in_2))
			begin
				local_bb5_c0_enter5_c0_eni44_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb5_c0_enter5_c0_eni44_stall_in_3))
			begin
				local_bb5_c0_enter5_c0_eni44_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb5_c0_enter5_c0_eni44_stall_in_4))
			begin
				local_bb5_c0_enter5_c0_eni44_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5_c0_ene16_stall_local;
wire local_bb5_c0_ene16;

assign local_bb5_c0_ene16 = local_bb5_c0_enter5_c0_eni44_NO_SHIFT_REG[8];

// This section implements an unregistered operation.
// 
wire local_bb5_c0_ene27_stall_local;
wire [31:0] local_bb5_c0_ene27;

assign local_bb5_c0_ene27 = local_bb5_c0_enter5_c0_eni44_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb5_c0_ene38_stall_local;
wire [31:0] local_bb5_c0_ene38;

assign local_bb5_c0_ene38 = local_bb5_c0_enter5_c0_eni44_NO_SHIFT_REG[95:64];

// This section implements an unregistered operation.
// 
wire local_bb5_c0_ene49_valid_out;
wire local_bb5_c0_ene49_stall_in;
wire local_bb5_c0_ene49_inputs_ready;
wire local_bb5_c0_ene49_stall_local;
wire local_bb5_c0_ene49;

assign local_bb5_c0_ene49_inputs_ready = local_bb5_c0_enter5_c0_eni44_valid_out_3_NO_SHIFT_REG;
assign local_bb5_c0_ene49 = local_bb5_c0_enter5_c0_eni44_NO_SHIFT_REG[96];
assign local_bb5_c0_ene49_valid_out = 1'b1;
assign local_bb5_c0_enter5_c0_eni44_stall_in_3 = 1'b0;

// This section implements an unregistered operation.
// 
wire SFC_2_VALID_2_2_0_valid_out;
wire SFC_2_VALID_2_2_0_stall_in;
wire SFC_2_VALID_2_2_0_inputs_ready;
wire SFC_2_VALID_2_2_0_stall_local;
wire SFC_2_VALID_2_2_0;

assign SFC_2_VALID_2_2_0_inputs_ready = local_bb5_c0_enter5_c0_eni44_valid_out_4_NO_SHIFT_REG;
assign SFC_2_VALID_2_2_0 = local_bb5_c0_enter5_c0_eni44_valid_bit_NO_SHIFT_REG;
assign SFC_2_VALID_2_2_0_valid_out = 1'b1;
assign local_bb5_c0_enter5_c0_eni44_stall_in_4 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb5_select34_stall_local;
wire [31:0] local_bb5_select34;

assign local_bb5_select34 = (local_bb5_c0_ene16 ? 32'h0 : local_bb5_c0_ene27);

// This section implements an unregistered operation.
// 
wire local_bb5_select34_valid_out;
wire local_bb5_select34_stall_in;
wire local_bb5_select37_valid_out;
wire local_bb5_select37_stall_in;
wire local_bb5_select37_inputs_ready;
wire local_bb5_select37_stall_local;
wire [31:0] local_bb5_select37;

assign local_bb5_select37_inputs_ready = (local_bb5_c0_enter5_c0_eni44_valid_out_0_NO_SHIFT_REG & local_bb5_c0_enter5_c0_eni44_valid_out_1_NO_SHIFT_REG & local_bb5_c0_enter5_c0_eni44_valid_out_2_NO_SHIFT_REG);
assign local_bb5_select37 = (local_bb5_c0_ene16 ? 32'h0 : local_bb5_c0_ene38);
assign local_bb5_select34_valid_out = 1'b1;
assign local_bb5_select37_valid_out = 1'b1;
assign local_bb5_c0_enter5_c0_eni44_stall_in_0 = 1'b0;
assign local_bb5_c0_enter5_c0_eni44_stall_in_1 = 1'b0;
assign local_bb5_c0_enter5_c0_eni44_stall_in_2 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb5_c0_ene49_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb5_c0_ene49_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb5_c0_ene49_0_NO_SHIFT_REG;
 logic rnode_2to3_bb5_c0_ene49_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb5_c0_ene49_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb5_c0_ene49_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb5_c0_ene49_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb5_c0_ene49_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb5_c0_ene49_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb5_c0_ene49_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb5_c0_ene49_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb5_c0_ene49_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb5_c0_ene49_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb5_c0_ene49),
	.data_out(rnode_2to3_bb5_c0_ene49_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb5_c0_ene49_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb5_c0_ene49_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb5_c0_ene49_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb5_c0_ene49_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb5_c0_ene49_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb5_c0_ene49_stall_in = 1'b0;
assign rnode_2to3_bb5_c0_ene49_0_NO_SHIFT_REG = rnode_2to3_bb5_c0_ene49_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb5_c0_ene49_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb5_c0_ene49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_2_3_0_inputs_ready;
 reg SFC_2_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_2_3_0_stall_in;
wire SFC_2_VALID_2_3_0_output_regs_ready;
 reg SFC_2_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_2_3_0_causedstall;

assign SFC_2_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_2_2_0_stall_in = 1'b0;
assign SFC_2_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_2_3_0_output_regs_ready)
		begin
			SFC_2_VALID_2_3_0_NO_SHIFT_REG <= SFC_2_VALID_2_2_0;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb5_div60_inputs_ready;
 reg local_bb5_div60_valid_out_NO_SHIFT_REG;
wire local_bb5_div60_stall_in;
wire local_bb5_div60_output_regs_ready;
wire [31:0] local_bb5_div60;
 reg local_bb5_div60_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb5_div60_valid_pipe_12_NO_SHIFT_REG;
wire local_bb5_div60_causedstall;

acl_fp_div_s5 fp_module_local_bb5_div60 (
	.clock(clock),
	.dataa(local_bb5_select34),
	.datab(local_bb5_select37),
	.enable(local_bb5_div60_output_regs_ready),
	.result(local_bb5_div60)
);


assign local_bb5_div60_inputs_ready = 1'b1;
assign local_bb5_div60_output_regs_ready = 1'b1;
assign local_bb5_select34_stall_in = 1'b0;
assign local_bb5_select37_stall_in = 1'b0;
assign local_bb5_div60_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_div60_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb5_div60_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_div60_output_regs_ready)
		begin
			local_bb5_div60_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb5_div60_valid_pipe_1_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_0_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_2_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_1_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_3_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_2_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_4_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_3_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_5_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_4_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_6_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_5_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_7_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_6_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_8_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_7_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_9_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_8_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_10_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_9_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_11_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_10_NO_SHIFT_REG;
			local_bb5_div60_valid_pipe_12_NO_SHIFT_REG <= local_bb5_div60_valid_pipe_11_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_div60_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_div60_output_regs_ready)
		begin
			local_bb5_div60_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb5_div60_stall_in))
			begin
				local_bb5_div60_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb5_c0_ene49_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb5_c0_ene49_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb5_c0_ene49_0_NO_SHIFT_REG;
 logic rnode_3to15_bb5_c0_ene49_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb5_c0_ene49_0_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb5_c0_ene49_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb5_c0_ene49_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb5_c0_ene49_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb5_c0_ene49_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb5_c0_ene49_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb5_c0_ene49_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb5_c0_ene49_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb5_c0_ene49_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(rnode_2to3_bb5_c0_ene49_0_NO_SHIFT_REG),
	.data_out(rnode_3to15_bb5_c0_ene49_0_reg_15_NO_SHIFT_REG)
);

defparam rnode_3to15_bb5_c0_ene49_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb5_c0_ene49_0_reg_15_fifo.DATA_WIDTH = 1;
defparam rnode_3to15_bb5_c0_ene49_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb5_c0_ene49_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb5_c0_ene49_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb5_c0_ene49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb5_c0_ene49_0_NO_SHIFT_REG = rnode_3to15_bb5_c0_ene49_0_reg_15_NO_SHIFT_REG;
assign rnode_3to15_bb5_c0_ene49_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb5_c0_ene49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_3_4_0_inputs_ready;
 reg SFC_2_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_3_4_0_stall_in;
wire SFC_2_VALID_3_4_0_output_regs_ready;
 reg SFC_2_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_3_4_0_causedstall;

assign SFC_2_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_stall_in = 1'b0;
assign SFC_2_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_3_4_0_output_regs_ready)
		begin
			SFC_2_VALID_3_4_0_NO_SHIFT_REG <= SFC_2_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb5_c0_ene49_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb5_c0_ene49_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb5_c0_ene49_0_NO_SHIFT_REG;
 logic rnode_15to16_bb5_c0_ene49_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb5_c0_ene49_0_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb5_c0_ene49_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb5_c0_ene49_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb5_c0_ene49_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb5_c0_ene49_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb5_c0_ene49_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb5_c0_ene49_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb5_c0_ene49_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb5_c0_ene49_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(rnode_3to15_bb5_c0_ene49_0_NO_SHIFT_REG),
	.data_out(rnode_15to16_bb5_c0_ene49_0_reg_16_NO_SHIFT_REG)
);

defparam rnode_15to16_bb5_c0_ene49_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb5_c0_ene49_0_reg_16_fifo.DATA_WIDTH = 1;
defparam rnode_15to16_bb5_c0_ene49_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb5_c0_ene49_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb5_c0_ene49_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb5_c0_ene49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb5_c0_ene49_0_NO_SHIFT_REG = rnode_15to16_bb5_c0_ene49_0_reg_16_NO_SHIFT_REG;
assign rnode_15to16_bb5_c0_ene49_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb5_c0_ene49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_4_5_0_inputs_ready;
 reg SFC_2_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_4_5_0_stall_in;
wire SFC_2_VALID_4_5_0_output_regs_ready;
 reg SFC_2_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_4_5_0_causedstall;

assign SFC_2_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_stall_in = 1'b0;
assign SFC_2_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_4_5_0_output_regs_ready)
		begin
			SFC_2_VALID_4_5_0_NO_SHIFT_REG <= SFC_2_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5__39_stall_local;
wire [31:0] local_bb5__39;

assign local_bb5__39 = (rnode_15to16_bb5_c0_ene49_0_NO_SHIFT_REG ? 32'h0 : local_bb5_div60);

// This section implements a registered operation.
// 
wire SFC_2_VALID_5_6_0_inputs_ready;
 reg SFC_2_VALID_5_6_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_5_6_0_stall_in;
wire SFC_2_VALID_5_6_0_output_regs_ready;
 reg SFC_2_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_5_6_0_causedstall;

assign SFC_2_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_stall_in = 1'b0;
assign SFC_2_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_5_6_0_output_regs_ready)
		begin
			SFC_2_VALID_5_6_0_NO_SHIFT_REG <= SFC_2_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5_c0_exi110_valid_out;
wire local_bb5_c0_exi110_stall_in;
wire local_bb5_c0_exi110_inputs_ready;
wire local_bb5_c0_exi110_stall_local;
wire [63:0] local_bb5_c0_exi110;

assign local_bb5_c0_exi110_inputs_ready = (local_bb5_div60_valid_out_NO_SHIFT_REG & rnode_15to16_bb5_c0_ene49_0_valid_out_NO_SHIFT_REG);
assign local_bb5_c0_exi110[31:0] = 32'bx;
assign local_bb5_c0_exi110[63:32] = local_bb5__39;
assign local_bb5_c0_exi110_valid_out = 1'b1;
assign local_bb5_div60_stall_in = 1'b0;
assign rnode_15to16_bb5_c0_ene49_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_2_VALID_6_7_0_inputs_ready;
 reg SFC_2_VALID_6_7_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_6_7_0_stall_in;
wire SFC_2_VALID_6_7_0_output_regs_ready;
 reg SFC_2_VALID_6_7_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_6_7_0_causedstall;

assign SFC_2_VALID_6_7_0_inputs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_stall_in = 1'b0;
assign SFC_2_VALID_6_7_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_6_7_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_6_7_0_output_regs_ready)
		begin
			SFC_2_VALID_6_7_0_NO_SHIFT_REG <= SFC_2_VALID_5_6_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_7_8_0_inputs_ready;
 reg SFC_2_VALID_7_8_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_7_8_0_stall_in;
wire SFC_2_VALID_7_8_0_output_regs_ready;
 reg SFC_2_VALID_7_8_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_7_8_0_causedstall;

assign SFC_2_VALID_7_8_0_inputs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_stall_in = 1'b0;
assign SFC_2_VALID_7_8_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_7_8_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_7_8_0_output_regs_ready)
		begin
			SFC_2_VALID_7_8_0_NO_SHIFT_REG <= SFC_2_VALID_6_7_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_8_9_0_inputs_ready;
 reg SFC_2_VALID_8_9_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in;
wire SFC_2_VALID_8_9_0_output_regs_ready;
 reg SFC_2_VALID_8_9_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_8_9_0_causedstall;

assign SFC_2_VALID_8_9_0_inputs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_stall_in = 1'b0;
assign SFC_2_VALID_8_9_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_8_9_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_8_9_0_output_regs_ready)
		begin
			SFC_2_VALID_8_9_0_NO_SHIFT_REG <= SFC_2_VALID_7_8_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_9_10_0_inputs_ready;
 reg SFC_2_VALID_9_10_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in;
wire SFC_2_VALID_9_10_0_output_regs_ready;
 reg SFC_2_VALID_9_10_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_9_10_0_causedstall;

assign SFC_2_VALID_9_10_0_inputs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in = 1'b0;
assign SFC_2_VALID_9_10_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_9_10_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_9_10_0_output_regs_ready)
		begin
			SFC_2_VALID_9_10_0_NO_SHIFT_REG <= SFC_2_VALID_8_9_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_10_11_0_inputs_ready;
 reg SFC_2_VALID_10_11_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_10_11_0_stall_in;
wire SFC_2_VALID_10_11_0_output_regs_ready;
 reg SFC_2_VALID_10_11_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_10_11_0_causedstall;

assign SFC_2_VALID_10_11_0_inputs_ready = 1'b1;
assign SFC_2_VALID_10_11_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in = 1'b0;
assign SFC_2_VALID_10_11_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_10_11_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_10_11_0_output_regs_ready)
		begin
			SFC_2_VALID_10_11_0_NO_SHIFT_REG <= SFC_2_VALID_9_10_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_11_12_0_inputs_ready;
 reg SFC_2_VALID_11_12_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_11_12_0_stall_in;
wire SFC_2_VALID_11_12_0_output_regs_ready;
 reg SFC_2_VALID_11_12_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_11_12_0_causedstall;

assign SFC_2_VALID_11_12_0_inputs_ready = 1'b1;
assign SFC_2_VALID_11_12_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_10_11_0_stall_in = 1'b0;
assign SFC_2_VALID_11_12_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_11_12_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_11_12_0_output_regs_ready)
		begin
			SFC_2_VALID_11_12_0_NO_SHIFT_REG <= SFC_2_VALID_10_11_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_12_13_0_inputs_ready;
 reg SFC_2_VALID_12_13_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_12_13_0_stall_in;
wire SFC_2_VALID_12_13_0_output_regs_ready;
 reg SFC_2_VALID_12_13_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_12_13_0_causedstall;

assign SFC_2_VALID_12_13_0_inputs_ready = 1'b1;
assign SFC_2_VALID_12_13_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_11_12_0_stall_in = 1'b0;
assign SFC_2_VALID_12_13_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_12_13_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_12_13_0_output_regs_ready)
		begin
			SFC_2_VALID_12_13_0_NO_SHIFT_REG <= SFC_2_VALID_11_12_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_13_14_0_inputs_ready;
 reg SFC_2_VALID_13_14_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_13_14_0_stall_in;
wire SFC_2_VALID_13_14_0_output_regs_ready;
 reg SFC_2_VALID_13_14_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_13_14_0_causedstall;

assign SFC_2_VALID_13_14_0_inputs_ready = 1'b1;
assign SFC_2_VALID_13_14_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_12_13_0_stall_in = 1'b0;
assign SFC_2_VALID_13_14_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_13_14_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_13_14_0_output_regs_ready)
		begin
			SFC_2_VALID_13_14_0_NO_SHIFT_REG <= SFC_2_VALID_12_13_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_14_15_0_inputs_ready;
 reg SFC_2_VALID_14_15_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_14_15_0_stall_in;
wire SFC_2_VALID_14_15_0_output_regs_ready;
 reg SFC_2_VALID_14_15_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_14_15_0_causedstall;

assign SFC_2_VALID_14_15_0_inputs_ready = 1'b1;
assign SFC_2_VALID_14_15_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_13_14_0_stall_in = 1'b0;
assign SFC_2_VALID_14_15_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_14_15_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_14_15_0_output_regs_ready)
		begin
			SFC_2_VALID_14_15_0_NO_SHIFT_REG <= SFC_2_VALID_13_14_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_15_16_0_inputs_ready;
 reg SFC_2_VALID_15_16_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_15_16_0_stall_in;
wire SFC_2_VALID_15_16_0_output_regs_ready;
 reg SFC_2_VALID_15_16_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_15_16_0_causedstall;

assign SFC_2_VALID_15_16_0_inputs_ready = 1'b1;
assign SFC_2_VALID_15_16_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_14_15_0_stall_in = 1'b0;
assign SFC_2_VALID_15_16_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_15_16_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_15_16_0_output_regs_ready)
		begin
			SFC_2_VALID_15_16_0_NO_SHIFT_REG <= SFC_2_VALID_14_15_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb5_c0_exit11_c0_exi110_inputs_ready;
 reg local_bb5_c0_exit11_c0_exi110_valid_out_NO_SHIFT_REG;
wire local_bb5_c0_exit11_c0_exi110_stall_in;
 reg [63:0] local_bb5_c0_exit11_c0_exi110_NO_SHIFT_REG;
wire [63:0] local_bb5_c0_exit11_c0_exi110_in;
wire local_bb5_c0_exit11_c0_exi110_valid;
wire local_bb5_c0_exit11_c0_exi110_causedstall;

acl_stall_free_sink local_bb5_c0_exit11_c0_exi110_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb5_c0_exi110),
	.data_out(local_bb5_c0_exit11_c0_exi110_in),
	.input_accepted(local_bb5_c0_enter5_c0_eni44_input_accepted),
	.valid_out(local_bb5_c0_exit11_c0_exi110_valid),
	.stall_in(~(local_bb5_c0_exit11_c0_exi110_output_regs_ready)),
	.stall_entry(local_bb5_c0_exit11_c0_exi110_entry_stall),
	.valid_in(local_bb5_c0_exit11_c0_exi110_valid_in),
	.IIphases(local_bb5_c0_exit11_c0_exi110_phases),
	.inc_pipelined_thread(local_bb5_c0_enter5_c0_eni44_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb5_c0_enter5_c0_eni44_dec_pipelined_thread)
);

defparam local_bb5_c0_exit11_c0_exi110_instance.DATA_WIDTH = 64;
defparam local_bb5_c0_exit11_c0_exi110_instance.PIPELINE_DEPTH = 20;
defparam local_bb5_c0_exit11_c0_exi110_instance.SHARINGII = 1;
defparam local_bb5_c0_exit11_c0_exi110_instance.SCHEDULEII = 1;
defparam local_bb5_c0_exit11_c0_exi110_instance.ALWAYS_THROTTLE = 0;

assign local_bb5_c0_exit11_c0_exi110_inputs_ready = 1'b1;
assign local_bb5_c0_exit11_c0_exi110_output_regs_ready = (&(~(local_bb5_c0_exit11_c0_exi110_valid_out_NO_SHIFT_REG) | ~(local_bb5_c0_exit11_c0_exi110_stall_in)));
assign local_bb5_c0_exit11_c0_exi110_valid_in = SFC_2_VALID_15_16_0_NO_SHIFT_REG;
assign local_bb5_c0_exi110_stall_in = 1'b0;
assign SFC_2_VALID_15_16_0_stall_in = 1'b0;
assign local_bb5_c0_exit11_c0_exi110_causedstall = (1'b1 && (1'b0 && !(~(local_bb5_c0_exit11_c0_exi110_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_c0_exit11_c0_exi110_NO_SHIFT_REG <= 'x;
		local_bb5_c0_exit11_c0_exi110_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_c0_exit11_c0_exi110_output_regs_ready)
		begin
			local_bb5_c0_exit11_c0_exi110_NO_SHIFT_REG <= local_bb5_c0_exit11_c0_exi110_in;
			local_bb5_c0_exit11_c0_exi110_valid_out_NO_SHIFT_REG <= local_bb5_c0_exit11_c0_exi110_valid;
		end
		else
		begin
			if (~(local_bb5_c0_exit11_c0_exi110_stall_in))
			begin
				local_bb5_c0_exit11_c0_exi110_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5_c0_exe112_valid_out;
wire local_bb5_c0_exe112_stall_in;
wire local_bb5_c0_exe112_inputs_ready;
wire local_bb5_c0_exe112_stall_local;
wire [31:0] local_bb5_c0_exe112;

assign local_bb5_c0_exe112_inputs_ready = local_bb5_c0_exit11_c0_exi110_valid_out_NO_SHIFT_REG;
assign local_bb5_c0_exe112 = local_bb5_c0_exit11_c0_exi110_NO_SHIFT_REG[63:32];
assign local_bb5_c0_exe112_valid_out = local_bb5_c0_exe112_inputs_ready;
assign local_bb5_c0_exe112_stall_local = local_bb5_c0_exe112_stall_in;
assign local_bb5_c0_exit11_c0_exi110_stall_in = (|local_bb5_c0_exe112_stall_local);

// This section implements a registered operation.
// 
wire local_bb5_st_c0_exe112_inputs_ready;
 reg local_bb5_st_c0_exe112_valid_out_NO_SHIFT_REG;
wire local_bb5_st_c0_exe112_stall_in;
wire local_bb5_st_c0_exe112_output_regs_ready;
wire local_bb5_st_c0_exe112_fu_stall_out;
wire local_bb5_st_c0_exe112_fu_valid_out;
wire local_bb5_st_c0_exe112_causedstall;

lsu_top lsu_local_bb5_st_c0_exe112 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb5_st_c0_exe112_fu_stall_out),
	.i_valid(local_bb5_st_c0_exe112_inputs_ready),
	.i_address((rnode_20to21_bb5_arrayidx15_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(local_bb5_c0_exe112),
	.i_cmpdata(),
	.i_predicate(1'b0),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb5_st_c0_exe112_output_regs_ready)),
	.o_valid(local_bb5_st_c0_exe112_fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb5_st_c0_exe112_active),
	.avm_address(avm_local_bb5_st_c0_exe112_address),
	.avm_read(avm_local_bb5_st_c0_exe112_read),
	.avm_readdata(avm_local_bb5_st_c0_exe112_readdata),
	.avm_write(avm_local_bb5_st_c0_exe112_write),
	.avm_writeack(avm_local_bb5_st_c0_exe112_writeack),
	.avm_burstcount(avm_local_bb5_st_c0_exe112_burstcount),
	.avm_writedata(avm_local_bb5_st_c0_exe112_writedata),
	.avm_byteenable(avm_local_bb5_st_c0_exe112_byteenable),
	.avm_waitrequest(avm_local_bb5_st_c0_exe112_waitrequest),
	.avm_readdatavalid(avm_local_bb5_st_c0_exe112_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb5_st_c0_exe112.AWIDTH = 33;
defparam lsu_local_bb5_st_c0_exe112.WIDTH_BYTES = 4;
defparam lsu_local_bb5_st_c0_exe112.MWIDTH_BYTES = 64;
defparam lsu_local_bb5_st_c0_exe112.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb5_st_c0_exe112.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb5_st_c0_exe112.READ = 0;
defparam lsu_local_bb5_st_c0_exe112.ATOMIC = 0;
defparam lsu_local_bb5_st_c0_exe112.WIDTH = 32;
defparam lsu_local_bb5_st_c0_exe112.MWIDTH = 512;
defparam lsu_local_bb5_st_c0_exe112.ATOMIC_WIDTH = 3;
defparam lsu_local_bb5_st_c0_exe112.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb5_st_c0_exe112.KERNEL_SIDE_MEM_LATENCY = 4;
defparam lsu_local_bb5_st_c0_exe112.MEMORY_SIDE_MEM_LATENCY = 8;
defparam lsu_local_bb5_st_c0_exe112.USE_WRITE_ACK = 0;
defparam lsu_local_bb5_st_c0_exe112.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb5_st_c0_exe112.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb5_st_c0_exe112.NUMBER_BANKS = 1;
defparam lsu_local_bb5_st_c0_exe112.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb5_st_c0_exe112.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb5_st_c0_exe112.USEINPUTFIFO = 0;
defparam lsu_local_bb5_st_c0_exe112.USECACHING = 0;
defparam lsu_local_bb5_st_c0_exe112.USEOUTPUTFIFO = 1;
defparam lsu_local_bb5_st_c0_exe112.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb5_st_c0_exe112.HIGH_FMAX = 1;
defparam lsu_local_bb5_st_c0_exe112.ADDRSPACE = 1;
defparam lsu_local_bb5_st_c0_exe112.STYLE = "BURST-COALESCED";
defparam lsu_local_bb5_st_c0_exe112.USE_BYTE_EN = 0;

assign local_bb5_st_c0_exe112_inputs_ready = (local_bb5_c0_exe112_valid_out & rnode_20to21_bb5_arrayidx15_0_valid_out_NO_SHIFT_REG);
assign local_bb5_st_c0_exe112_output_regs_ready = (&(~(local_bb5_st_c0_exe112_valid_out_NO_SHIFT_REG) | ~(local_bb5_st_c0_exe112_stall_in)));
assign local_bb5_c0_exe112_stall_in = (local_bb5_st_c0_exe112_fu_stall_out | ~(local_bb5_st_c0_exe112_inputs_ready));
assign rnode_20to21_bb5_arrayidx15_0_stall_in_NO_SHIFT_REG = (local_bb5_st_c0_exe112_fu_stall_out | ~(local_bb5_st_c0_exe112_inputs_ready));
assign local_bb5_st_c0_exe112_causedstall = (local_bb5_st_c0_exe112_inputs_ready && (local_bb5_st_c0_exe112_fu_stall_out && !(~(local_bb5_st_c0_exe112_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_st_c0_exe112_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_st_c0_exe112_output_regs_ready)
		begin
			local_bb5_st_c0_exe112_valid_out_NO_SHIFT_REG <= local_bb5_st_c0_exe112_fu_valid_out;
		end
		else
		begin
			if (~(local_bb5_st_c0_exe112_stall_in))
			begin
				local_bb5_st_c0_exe112_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_25to25_bb5_st_c0_exe112_valid_out;
wire rstag_25to25_bb5_st_c0_exe112_stall_in;
wire rstag_25to25_bb5_st_c0_exe112_inputs_ready;
wire rstag_25to25_bb5_st_c0_exe112_stall_local;
 reg rstag_25to25_bb5_st_c0_exe112_staging_valid_NO_SHIFT_REG;
wire rstag_25to25_bb5_st_c0_exe112_combined_valid;

assign rstag_25to25_bb5_st_c0_exe112_inputs_ready = local_bb5_st_c0_exe112_valid_out_NO_SHIFT_REG;
assign rstag_25to25_bb5_st_c0_exe112_combined_valid = (rstag_25to25_bb5_st_c0_exe112_staging_valid_NO_SHIFT_REG | rstag_25to25_bb5_st_c0_exe112_inputs_ready);
assign rstag_25to25_bb5_st_c0_exe112_valid_out = rstag_25to25_bb5_st_c0_exe112_combined_valid;
assign rstag_25to25_bb5_st_c0_exe112_stall_local = rstag_25to25_bb5_st_c0_exe112_stall_in;
assign local_bb5_st_c0_exe112_stall_in = (|rstag_25to25_bb5_st_c0_exe112_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_25to25_bb5_st_c0_exe112_staging_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (rstag_25to25_bb5_st_c0_exe112_stall_local)
		begin
			if (~(rstag_25to25_bb5_st_c0_exe112_staging_valid_NO_SHIFT_REG))
			begin
				rstag_25to25_bb5_st_c0_exe112_staging_valid_NO_SHIFT_REG <= rstag_25to25_bb5_st_c0_exe112_inputs_ready;
			end
		end
		else
		begin
			rstag_25to25_bb5_st_c0_exe112_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
wire branch_var__output_regs_ready;

assign branch_var__inputs_ready = (rnode_24to25_input_acl_hw_wg_id_0_valid_out_NO_SHIFT_REG & rstag_25to25_bb5_st_c0_exe112_valid_out);
assign branch_var__output_regs_ready = ~(stall_in);
assign rnode_24to25_input_acl_hw_wg_id_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_25to25_bb5_st_c0_exe112_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out = branch_var__inputs_ready;
assign lvb_input_acl_hw_wg_id = rnode_24to25_input_acl_hw_wg_id_0_NO_SHIFT_REG;

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_function
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		input [31:0] 		input_acl_hw_wg_id,
		output 		stall_out,
		input 		valid_in,
		output [31:0] 		output_0,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input [511:0] 		avm_local_bb1_ld__readdata,
		input 		avm_local_bb1_ld__readdatavalid,
		input 		avm_local_bb1_ld__waitrequest,
		output [32:0] 		avm_local_bb1_ld__address,
		output 		avm_local_bb1_ld__read,
		output 		avm_local_bb1_ld__write,
		input 		avm_local_bb1_ld__writeack,
		output [511:0] 		avm_local_bb1_ld__writedata,
		output [63:0] 		avm_local_bb1_ld__byteenable,
		output [4:0] 		avm_local_bb1_ld__burstcount,
		input [511:0] 		avm_local_bb3_ld__readdata,
		input 		avm_local_bb3_ld__readdatavalid,
		input 		avm_local_bb3_ld__waitrequest,
		output [32:0] 		avm_local_bb3_ld__address,
		output 		avm_local_bb3_ld__read,
		output 		avm_local_bb3_ld__write,
		input 		avm_local_bb3_ld__writeack,
		output [511:0] 		avm_local_bb3_ld__writedata,
		output [63:0] 		avm_local_bb3_ld__byteenable,
		output [4:0] 		avm_local_bb3_ld__burstcount,
		input [511:0] 		avm_local_bb3_ld__u12_readdata,
		input 		avm_local_bb3_ld__u12_readdatavalid,
		input 		avm_local_bb3_ld__u12_waitrequest,
		output [32:0] 		avm_local_bb3_ld__u12_address,
		output 		avm_local_bb3_ld__u12_read,
		output 		avm_local_bb3_ld__u12_write,
		input 		avm_local_bb3_ld__u12_writeack,
		output [511:0] 		avm_local_bb3_ld__u12_writedata,
		output [63:0] 		avm_local_bb3_ld__u12_byteenable,
		output [4:0] 		avm_local_bb3_ld__u12_burstcount,
		input [511:0] 		avm_local_bb3_ld__u13_readdata,
		input 		avm_local_bb3_ld__u13_readdatavalid,
		input 		avm_local_bb3_ld__u13_waitrequest,
		output [32:0] 		avm_local_bb3_ld__u13_address,
		output 		avm_local_bb3_ld__u13_read,
		output 		avm_local_bb3_ld__u13_write,
		input 		avm_local_bb3_ld__u13_writeack,
		output [511:0] 		avm_local_bb3_ld__u13_writedata,
		output [63:0] 		avm_local_bb3_ld__u13_byteenable,
		output [4:0] 		avm_local_bb3_ld__u13_burstcount,
		input [511:0] 		avm_local_bb5_st_c0_exe112_readdata,
		input 		avm_local_bb5_st_c0_exe112_readdatavalid,
		input 		avm_local_bb5_st_c0_exe112_waitrequest,
		output [32:0] 		avm_local_bb5_st_c0_exe112_address,
		output 		avm_local_bb5_st_c0_exe112_read,
		output 		avm_local_bb5_st_c0_exe112_write,
		input 		avm_local_bb5_st_c0_exe112_writeack,
		output [511:0] 		avm_local_bb5_st_c0_exe112_writedata,
		output [63:0] 		avm_local_bb5_st_c0_exe112_byteenable,
		output [4:0] 		avm_local_bb5_st_c0_exe112_burstcount,
		input 		start,
		input [31:0] 		input_r,
		input [31:0] 		input_global_size_0,
		input [31:0] 		input_global_size_1,
		input [31:0] 		input_e_d,
		input 		clock2x,
		input [63:0] 		input_in,
		input [63:0] 		input_gaussian,
		input [63:0] 		input_out,
		output reg 		has_a_write_pending,
		output reg 		has_a_lsu_active
	);


wire [31:0] cur_cycle;
wire bb_0_stall_out;
wire bb_0_valid_out;
wire bb_0_lvb_bb0_cmp1622;
wire [31:0] bb_0_lvb_bb0_sub25;
wire [31:0] bb_0_lvb_bb0_sub29;
wire [31:0] bb_0_lvb_bb0_mul50;
wire [63:0] bb_0_lvb_bb0_var_;
wire [63:0] bb_0_lvb_bb0_var__u0;
wire [31:0] bb_0_lvb_input_global_id_0;
wire [31:0] bb_0_lvb_input_global_id_1;
wire [31:0] bb_0_lvb_input_acl_hw_wg_id;
wire bb_1_stall_out;
wire bb_1_valid_out;
wire [63:0] bb_1_lvb_bb1_idxprom;
wire [31:0] bb_1_lvb_bb1_ld_;
wire bb_1_lvb_bb1_cmp;
wire bb_1_lvb_bb1_var_;
wire [31:0] bb_1_lvb_input_global_id_0;
wire [31:0] bb_1_lvb_input_global_id_1;
wire [31:0] bb_1_lvb_input_acl_hw_wg_id;
wire bb_1_local_bb1_ld__active;
wire bb_2_stall_out_0;
wire bb_2_stall_out_1;
wire bb_2_valid_out;
wire [63:0] bb_2_lvb_idxprom;
wire [31:0] bb_2_lvb_ld_;
wire bb_2_lvb_cmp;
wire bb_2_lvb_var__u5;
wire [63:0] bb_2_lvb_indvars_iv29;
wire [31:0] bb_2_lvb_t_024;
wire [31:0] bb_2_lvb_sum_023;
wire [31:0] bb_2_lvb_bb2_sub25_add24;
wire [63:0] bb_2_lvb_bb2_arrayidx43;
wire [31:0] bb_2_lvb_input_global_id_0;
wire [31:0] bb_2_lvb_input_global_id_1;
wire [31:0] bb_2_lvb_input_acl_hw_wg_id;
wire bb_3_stall_out_0;
wire bb_3_stall_out_1;
wire bb_3_valid_out_0;
wire [63:0] bb_3_lvb_idxprom_0;
wire [31:0] bb_3_lvb_ld__0;
wire bb_3_lvb_cmp_0;
wire bb_3_lvb_var__u8_0;
wire [63:0] bb_3_lvb_indvars_iv29_0;
wire [31:0] bb_3_lvb_sub25_add24_0;
wire [63:0] bb_3_lvb_arrayidx43_0;
wire [63:0] bb_3_lvb_bb3_indvars_iv_next_0;
wire [31:0] bb_3_lvb_bb3_c0_exe1_0;
wire [31:0] bb_3_lvb_bb3_c0_exe2_0;
wire [31:0] bb_3_lvb_input_global_id_0_0;
wire [31:0] bb_3_lvb_input_global_id_1_0;
wire [31:0] bb_3_lvb_input_acl_hw_wg_id_0;
wire bb_3_valid_out_1;
wire [63:0] bb_3_lvb_idxprom_1;
wire [31:0] bb_3_lvb_ld__1;
wire bb_3_lvb_cmp_1;
wire bb_3_lvb_var__u8_1;
wire [63:0] bb_3_lvb_indvars_iv29_1;
wire [31:0] bb_3_lvb_sub25_add24_1;
wire [63:0] bb_3_lvb_arrayidx43_1;
wire [63:0] bb_3_lvb_bb3_indvars_iv_next_1;
wire [31:0] bb_3_lvb_bb3_c0_exe1_1;
wire [31:0] bb_3_lvb_bb3_c0_exe2_1;
wire [31:0] bb_3_lvb_input_global_id_0_1;
wire [31:0] bb_3_lvb_input_global_id_1_1;
wire [31:0] bb_3_lvb_input_acl_hw_wg_id_1;
wire bb_3_local_bb3_ld__active;
wire bb_3_local_bb3_ld__u12_active;
wire bb_3_local_bb3_ld__u13_active;
wire bb_4_stall_out;
wire bb_4_valid_out_0;
wire [63:0] bb_4_lvb_idxprom_0;
wire [31:0] bb_4_lvb_ld__0;
wire bb_4_lvb_cmp_0;
wire bb_4_lvb_var__u96_0;
wire [31:0] bb_4_lvb_c0_exe1_0;
wire [31:0] bb_4_lvb_c0_exe2_0;
wire [63:0] bb_4_lvb_bb4_indvars_iv_next30_0;
wire [31:0] bb_4_lvb_input_global_id_0_0;
wire [31:0] bb_4_lvb_input_global_id_1_0;
wire [31:0] bb_4_lvb_input_acl_hw_wg_id_0;
wire bb_4_valid_out_1;
wire [63:0] bb_4_lvb_idxprom_1;
wire [31:0] bb_4_lvb_ld__1;
wire bb_4_lvb_cmp_1;
wire bb_4_lvb_var__u96_1;
wire [31:0] bb_4_lvb_c0_exe1_1;
wire [31:0] bb_4_lvb_c0_exe2_1;
wire [63:0] bb_4_lvb_bb4_indvars_iv_next30_1;
wire [31:0] bb_4_lvb_input_global_id_0_1;
wire [31:0] bb_4_lvb_input_global_id_1_1;
wire [31:0] bb_4_lvb_input_acl_hw_wg_id_1;
wire bb_5_stall_out;
wire bb_5_valid_out;
wire [31:0] bb_5_lvb_input_acl_hw_wg_id;
wire bb_5_local_bb5_st_c0_exe112_active;
wire loop_limiter_0_stall_out;
wire loop_limiter_0_valid_out;
wire loop_limiter_1_stall_out;
wire loop_limiter_1_valid_out;
wire writes_pending;
wire [4:0] lsus_active;

AOCbilateralFilterkernel_basic_block_0 AOCbilateralFilterkernel_basic_block_0 (
	.clock(clock),
	.resetn(resetn),
	.start(start),
	.input_r(input_r),
	.input_global_size_0(input_global_size_0),
	.input_global_size_1(input_global_size_1),
	.input_e_d(input_e_d),
	.valid_in(valid_in),
	.stall_out(bb_0_stall_out),
	.input_global_id_0(input_global_id_0),
	.input_global_id_1(input_global_id_1),
	.input_acl_hw_wg_id(input_acl_hw_wg_id),
	.valid_out(bb_0_valid_out),
	.stall_in(bb_1_stall_out),
	.lvb_bb0_cmp1622(bb_0_lvb_bb0_cmp1622),
	.lvb_bb0_sub25(bb_0_lvb_bb0_sub25),
	.lvb_bb0_sub29(bb_0_lvb_bb0_sub29),
	.lvb_bb0_mul50(bb_0_lvb_bb0_mul50),
	.lvb_bb0_var_(bb_0_lvb_bb0_var_),
	.lvb_bb0_var__u0(bb_0_lvb_bb0_var__u0),
	.lvb_input_global_id_0(bb_0_lvb_input_global_id_0),
	.lvb_input_global_id_1(bb_0_lvb_input_global_id_1),
	.lvb_input_acl_hw_wg_id(bb_0_lvb_input_acl_hw_wg_id),
	.workgroup_size(workgroup_size)
);


AOCbilateralFilterkernel_basic_block_1 AOCbilateralFilterkernel_basic_block_1 (
	.clock(clock),
	.resetn(resetn),
	.input_global_size_0(input_global_size_0),
	.input_in(input_in),
	.input_wii_cmp1622(bb_0_lvb_bb0_cmp1622),
	.input_wii_sub25(bb_0_lvb_bb0_sub25),
	.input_wii_sub29(bb_0_lvb_bb0_sub29),
	.input_wii_mul50(bb_0_lvb_bb0_mul50),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u3(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_0_valid_out),
	.stall_out(bb_1_stall_out),
	.input_global_id_0(bb_0_lvb_input_global_id_0),
	.input_global_id_1(bb_0_lvb_input_global_id_1),
	.input_acl_hw_wg_id(bb_0_lvb_input_acl_hw_wg_id),
	.valid_out(bb_1_valid_out),
	.stall_in(loop_limiter_0_stall_out),
	.lvb_bb1_idxprom(bb_1_lvb_bb1_idxprom),
	.lvb_bb1_ld_(bb_1_lvb_bb1_ld_),
	.lvb_bb1_cmp(bb_1_lvb_bb1_cmp),
	.lvb_bb1_var_(bb_1_lvb_bb1_var_),
	.lvb_input_global_id_0(bb_1_lvb_input_global_id_0),
	.lvb_input_global_id_1(bb_1_lvb_input_global_id_1),
	.lvb_input_acl_hw_wg_id(bb_1_lvb_input_acl_hw_wg_id),
	.workgroup_size(workgroup_size),
	.start(start),
	.avm_local_bb1_ld__readdata(avm_local_bb1_ld__readdata),
	.avm_local_bb1_ld__readdatavalid(avm_local_bb1_ld__readdatavalid),
	.avm_local_bb1_ld__waitrequest(avm_local_bb1_ld__waitrequest),
	.avm_local_bb1_ld__address(avm_local_bb1_ld__address),
	.avm_local_bb1_ld__read(avm_local_bb1_ld__read),
	.avm_local_bb1_ld__write(avm_local_bb1_ld__write),
	.avm_local_bb1_ld__writeack(avm_local_bb1_ld__writeack),
	.avm_local_bb1_ld__writedata(avm_local_bb1_ld__writedata),
	.avm_local_bb1_ld__byteenable(avm_local_bb1_ld__byteenable),
	.avm_local_bb1_ld__burstcount(avm_local_bb1_ld__burstcount),
	.local_bb1_ld__active(bb_1_local_bb1_ld__active),
	.clock2x(clock2x)
);


AOCbilateralFilterkernel_basic_block_2 AOCbilateralFilterkernel_basic_block_2 (
	.clock(clock),
	.resetn(resetn),
	.input_gaussian(input_gaussian),
	.input_wii_sub25(bb_0_lvb_bb0_sub25),
	.input_wii_sub29(bb_0_lvb_bb0_sub29),
	.input_wii_mul50(bb_0_lvb_bb0_mul50),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u4(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_4_valid_out_1),
	.stall_out_0(bb_2_stall_out_0),
	.input_idxprom_0(bb_4_lvb_idxprom_1),
	.input_ld__0(bb_4_lvb_ld__1),
	.input_cmp_0(bb_4_lvb_cmp_1),
	.input_var__u5_0(bb_4_lvb_var__u96_1),
	.input_indvars_iv29_0(bb_4_lvb_bb4_indvars_iv_next30_1),
	.input_t_024_0(bb_4_lvb_c0_exe2_1),
	.input_sum_023_0(bb_4_lvb_c0_exe1_1),
	.input_global_id_0_0(bb_4_lvb_input_global_id_0_1),
	.input_global_id_1_0(bb_4_lvb_input_global_id_1_1),
	.input_acl_hw_wg_id_0(bb_4_lvb_input_acl_hw_wg_id_1),
	.valid_in_1(loop_limiter_0_valid_out),
	.stall_out_1(bb_2_stall_out_1),
	.input_idxprom_1(bb_1_lvb_bb1_idxprom),
	.input_ld__1(bb_1_lvb_bb1_ld_),
	.input_cmp_1(bb_1_lvb_bb1_cmp),
	.input_var__u5_1(bb_1_lvb_bb1_var_),
	.input_indvars_iv29_1(bb_0_lvb_bb0_var_),
	.input_t_024_1(32'h0),
	.input_sum_023_1(32'h0),
	.input_global_id_0_1(bb_1_lvb_input_global_id_0),
	.input_global_id_1_1(bb_1_lvb_input_global_id_1),
	.input_acl_hw_wg_id_1(bb_1_lvb_input_acl_hw_wg_id),
	.valid_out(bb_2_valid_out),
	.stall_in(loop_limiter_1_stall_out),
	.lvb_idxprom(bb_2_lvb_idxprom),
	.lvb_ld_(bb_2_lvb_ld_),
	.lvb_cmp(bb_2_lvb_cmp),
	.lvb_var__u5(bb_2_lvb_var__u5),
	.lvb_indvars_iv29(bb_2_lvb_indvars_iv29),
	.lvb_t_024(bb_2_lvb_t_024),
	.lvb_sum_023(bb_2_lvb_sum_023),
	.lvb_bb2_sub25_add24(bb_2_lvb_bb2_sub25_add24),
	.lvb_bb2_arrayidx43(bb_2_lvb_bb2_arrayidx43),
	.lvb_input_global_id_0(bb_2_lvb_input_global_id_0),
	.lvb_input_global_id_1(bb_2_lvb_input_global_id_1),
	.lvb_input_acl_hw_wg_id(bb_2_lvb_input_acl_hw_wg_id),
	.workgroup_size(workgroup_size),
	.start(start)
);


AOCbilateralFilterkernel_basic_block_3 AOCbilateralFilterkernel_basic_block_3 (
	.clock(clock),
	.resetn(resetn),
	.input_gaussian(input_gaussian),
	.input_r(input_r),
	.input_global_size_0(input_global_size_0),
	.input_in(input_in),
	.input_wii_sub25(bb_0_lvb_bb0_sub25),
	.input_wii_sub29(bb_0_lvb_bb0_sub29),
	.input_wii_mul50(bb_0_lvb_bb0_mul50),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u7(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_3_valid_out_1),
	.stall_out_0(bb_3_stall_out_0),
	.input_idxprom_0(bb_3_lvb_idxprom_1),
	.input_ld__0(bb_3_lvb_ld__1),
	.input_cmp_0(bb_3_lvb_cmp_1),
	.input_var__u8_0(bb_3_lvb_var__u8_1),
	.input_indvars_iv29_0(bb_3_lvb_indvars_iv29_1),
	.input_sub25_add24_0(bb_3_lvb_sub25_add24_1),
	.input_arrayidx43_0(bb_3_lvb_arrayidx43_1),
	.input_indvars_iv_0(bb_3_lvb_bb3_indvars_iv_next_1),
	.input_t_119_0(bb_3_lvb_bb3_c0_exe2_1),
	.input_sum_118_0(bb_3_lvb_bb3_c0_exe1_1),
	.input_global_id_0_0(bb_3_lvb_input_global_id_0_1),
	.input_global_id_1_0(bb_3_lvb_input_global_id_1_1),
	.input_acl_hw_wg_id_0(bb_3_lvb_input_acl_hw_wg_id_1),
	.valid_in_1(loop_limiter_1_valid_out),
	.stall_out_1(bb_3_stall_out_1),
	.input_idxprom_1(bb_2_lvb_idxprom),
	.input_ld__1(bb_2_lvb_ld_),
	.input_cmp_1(bb_2_lvb_cmp),
	.input_var__u8_1(bb_2_lvb_var__u5),
	.input_indvars_iv29_1(bb_2_lvb_indvars_iv29),
	.input_sub25_add24_1(bb_2_lvb_bb2_sub25_add24),
	.input_arrayidx43_1(bb_2_lvb_bb2_arrayidx43),
	.input_indvars_iv_1(bb_0_lvb_bb0_var_),
	.input_t_119_1(bb_2_lvb_t_024),
	.input_sum_118_1(bb_2_lvb_sum_023),
	.input_global_id_0_1(bb_2_lvb_input_global_id_0),
	.input_global_id_1_1(bb_2_lvb_input_global_id_1),
	.input_acl_hw_wg_id_1(bb_2_lvb_input_acl_hw_wg_id),
	.valid_out_0(bb_3_valid_out_0),
	.stall_in_0(bb_4_stall_out),
	.lvb_idxprom_0(bb_3_lvb_idxprom_0),
	.lvb_ld__0(bb_3_lvb_ld__0),
	.lvb_cmp_0(bb_3_lvb_cmp_0),
	.lvb_var__u8_0(bb_3_lvb_var__u8_0),
	.lvb_indvars_iv29_0(bb_3_lvb_indvars_iv29_0),
	.lvb_sub25_add24_0(bb_3_lvb_sub25_add24_0),
	.lvb_arrayidx43_0(bb_3_lvb_arrayidx43_0),
	.lvb_bb3_indvars_iv_next_0(bb_3_lvb_bb3_indvars_iv_next_0),
	.lvb_bb3_c0_exe1_0(bb_3_lvb_bb3_c0_exe1_0),
	.lvb_bb3_c0_exe2_0(bb_3_lvb_bb3_c0_exe2_0),
	.lvb_input_global_id_0_0(bb_3_lvb_input_global_id_0_0),
	.lvb_input_global_id_1_0(bb_3_lvb_input_global_id_1_0),
	.lvb_input_acl_hw_wg_id_0(bb_3_lvb_input_acl_hw_wg_id_0),
	.valid_out_1(bb_3_valid_out_1),
	.stall_in_1(bb_3_stall_out_0),
	.lvb_idxprom_1(bb_3_lvb_idxprom_1),
	.lvb_ld__1(bb_3_lvb_ld__1),
	.lvb_cmp_1(bb_3_lvb_cmp_1),
	.lvb_var__u8_1(bb_3_lvb_var__u8_1),
	.lvb_indvars_iv29_1(bb_3_lvb_indvars_iv29_1),
	.lvb_sub25_add24_1(bb_3_lvb_sub25_add24_1),
	.lvb_arrayidx43_1(bb_3_lvb_arrayidx43_1),
	.lvb_bb3_indvars_iv_next_1(bb_3_lvb_bb3_indvars_iv_next_1),
	.lvb_bb3_c0_exe1_1(bb_3_lvb_bb3_c0_exe1_1),
	.lvb_bb3_c0_exe2_1(bb_3_lvb_bb3_c0_exe2_1),
	.lvb_input_global_id_0_1(bb_3_lvb_input_global_id_0_1),
	.lvb_input_global_id_1_1(bb_3_lvb_input_global_id_1_1),
	.lvb_input_acl_hw_wg_id_1(bb_3_lvb_input_acl_hw_wg_id_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.avm_local_bb3_ld__readdata(avm_local_bb3_ld__readdata),
	.avm_local_bb3_ld__readdatavalid(avm_local_bb3_ld__readdatavalid),
	.avm_local_bb3_ld__waitrequest(avm_local_bb3_ld__waitrequest),
	.avm_local_bb3_ld__address(avm_local_bb3_ld__address),
	.avm_local_bb3_ld__read(avm_local_bb3_ld__read),
	.avm_local_bb3_ld__write(avm_local_bb3_ld__write),
	.avm_local_bb3_ld__writeack(avm_local_bb3_ld__writeack),
	.avm_local_bb3_ld__writedata(avm_local_bb3_ld__writedata),
	.avm_local_bb3_ld__byteenable(avm_local_bb3_ld__byteenable),
	.avm_local_bb3_ld__burstcount(avm_local_bb3_ld__burstcount),
	.local_bb3_ld__active(bb_3_local_bb3_ld__active),
	.clock2x(clock2x),
	.avm_local_bb3_ld__u12_readdata(avm_local_bb3_ld__u12_readdata),
	.avm_local_bb3_ld__u12_readdatavalid(avm_local_bb3_ld__u12_readdatavalid),
	.avm_local_bb3_ld__u12_waitrequest(avm_local_bb3_ld__u12_waitrequest),
	.avm_local_bb3_ld__u12_address(avm_local_bb3_ld__u12_address),
	.avm_local_bb3_ld__u12_read(avm_local_bb3_ld__u12_read),
	.avm_local_bb3_ld__u12_write(avm_local_bb3_ld__u12_write),
	.avm_local_bb3_ld__u12_writeack(avm_local_bb3_ld__u12_writeack),
	.avm_local_bb3_ld__u12_writedata(avm_local_bb3_ld__u12_writedata),
	.avm_local_bb3_ld__u12_byteenable(avm_local_bb3_ld__u12_byteenable),
	.avm_local_bb3_ld__u12_burstcount(avm_local_bb3_ld__u12_burstcount),
	.local_bb3_ld__u12_active(bb_3_local_bb3_ld__u12_active),
	.avm_local_bb3_ld__u13_readdata(avm_local_bb3_ld__u13_readdata),
	.avm_local_bb3_ld__u13_readdatavalid(avm_local_bb3_ld__u13_readdatavalid),
	.avm_local_bb3_ld__u13_waitrequest(avm_local_bb3_ld__u13_waitrequest),
	.avm_local_bb3_ld__u13_address(avm_local_bb3_ld__u13_address),
	.avm_local_bb3_ld__u13_read(avm_local_bb3_ld__u13_read),
	.avm_local_bb3_ld__u13_write(avm_local_bb3_ld__u13_write),
	.avm_local_bb3_ld__u13_writeack(avm_local_bb3_ld__u13_writeack),
	.avm_local_bb3_ld__u13_writedata(avm_local_bb3_ld__u13_writedata),
	.avm_local_bb3_ld__u13_byteenable(avm_local_bb3_ld__u13_byteenable),
	.avm_local_bb3_ld__u13_burstcount(avm_local_bb3_ld__u13_burstcount),
	.local_bb3_ld__u13_active(bb_3_local_bb3_ld__u13_active)
);


AOCbilateralFilterkernel_basic_block_4 AOCbilateralFilterkernel_basic_block_4 (
	.clock(clock),
	.resetn(resetn),
	.input_r(input_r),
	.input_wii_sub25(bb_0_lvb_bb0_sub25),
	.input_wii_sub29(bb_0_lvb_bb0_sub29),
	.input_wii_mul50(bb_0_lvb_bb0_mul50),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u95(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_3_valid_out_0),
	.stall_out(bb_4_stall_out),
	.input_idxprom(bb_3_lvb_idxprom_0),
	.input_ld_(bb_3_lvb_ld__0),
	.input_cmp(bb_3_lvb_cmp_0),
	.input_var__u96(bb_3_lvb_var__u8_0),
	.input_indvars_iv29(bb_3_lvb_indvars_iv29_0),
	.input_c0_exe1(bb_3_lvb_bb3_c0_exe1_0),
	.input_c0_exe2(bb_3_lvb_bb3_c0_exe2_0),
	.input_global_id_0(bb_3_lvb_input_global_id_0_0),
	.input_global_id_1(bb_3_lvb_input_global_id_1_0),
	.input_acl_hw_wg_id(bb_3_lvb_input_acl_hw_wg_id_0),
	.valid_out_0(bb_4_valid_out_0),
	.stall_in_0(bb_5_stall_out),
	.lvb_idxprom_0(bb_4_lvb_idxprom_0),
	.lvb_ld__0(bb_4_lvb_ld__0),
	.lvb_cmp_0(bb_4_lvb_cmp_0),
	.lvb_var__u96_0(bb_4_lvb_var__u96_0),
	.lvb_c0_exe1_0(bb_4_lvb_c0_exe1_0),
	.lvb_c0_exe2_0(bb_4_lvb_c0_exe2_0),
	.lvb_bb4_indvars_iv_next30_0(bb_4_lvb_bb4_indvars_iv_next30_0),
	.lvb_input_global_id_0_0(bb_4_lvb_input_global_id_0_0),
	.lvb_input_global_id_1_0(bb_4_lvb_input_global_id_1_0),
	.lvb_input_acl_hw_wg_id_0(bb_4_lvb_input_acl_hw_wg_id_0),
	.valid_out_1(bb_4_valid_out_1),
	.stall_in_1(bb_2_stall_out_0),
	.lvb_idxprom_1(bb_4_lvb_idxprom_1),
	.lvb_ld__1(bb_4_lvb_ld__1),
	.lvb_cmp_1(bb_4_lvb_cmp_1),
	.lvb_var__u96_1(bb_4_lvb_var__u96_1),
	.lvb_c0_exe1_1(bb_4_lvb_c0_exe1_1),
	.lvb_c0_exe2_1(bb_4_lvb_c0_exe2_1),
	.lvb_bb4_indvars_iv_next30_1(bb_4_lvb_bb4_indvars_iv_next30_1),
	.lvb_input_global_id_0_1(bb_4_lvb_input_global_id_0_1),
	.lvb_input_global_id_1_1(bb_4_lvb_input_global_id_1_1),
	.lvb_input_acl_hw_wg_id_1(bb_4_lvb_input_acl_hw_wg_id_1),
	.workgroup_size(workgroup_size),
	.start(start)
);


AOCbilateralFilterkernel_basic_block_5 AOCbilateralFilterkernel_basic_block_5 (
	.clock(clock),
	.resetn(resetn),
	.input_out(input_out),
	.valid_in(bb_4_valid_out_0),
	.stall_out(bb_5_stall_out),
	.input_idxprom(bb_4_lvb_idxprom_0),
	.input_cmp(bb_4_lvb_cmp_0),
	.input_var_(bb_4_lvb_var__u96_0),
	.input_c0_exe1(bb_4_lvb_c0_exe1_0),
	.input_c0_exe2(bb_4_lvb_c0_exe2_0),
	.input_acl_hw_wg_id(bb_4_lvb_input_acl_hw_wg_id_0),
	.valid_out(bb_5_valid_out),
	.stall_in(stall_in),
	.lvb_input_acl_hw_wg_id(bb_5_lvb_input_acl_hw_wg_id),
	.workgroup_size(workgroup_size),
	.start(start),
	.avm_local_bb5_st_c0_exe112_readdata(avm_local_bb5_st_c0_exe112_readdata),
	.avm_local_bb5_st_c0_exe112_readdatavalid(avm_local_bb5_st_c0_exe112_readdatavalid),
	.avm_local_bb5_st_c0_exe112_waitrequest(avm_local_bb5_st_c0_exe112_waitrequest),
	.avm_local_bb5_st_c0_exe112_address(avm_local_bb5_st_c0_exe112_address),
	.avm_local_bb5_st_c0_exe112_read(avm_local_bb5_st_c0_exe112_read),
	.avm_local_bb5_st_c0_exe112_write(avm_local_bb5_st_c0_exe112_write),
	.avm_local_bb5_st_c0_exe112_writeack(avm_local_bb5_st_c0_exe112_writeack),
	.avm_local_bb5_st_c0_exe112_writedata(avm_local_bb5_st_c0_exe112_writedata),
	.avm_local_bb5_st_c0_exe112_byteenable(avm_local_bb5_st_c0_exe112_byteenable),
	.avm_local_bb5_st_c0_exe112_burstcount(avm_local_bb5_st_c0_exe112_burstcount),
	.local_bb5_st_c0_exe112_active(bb_5_local_bb5_st_c0_exe112_active),
	.clock2x(clock2x)
);


acl_loop_limiter loop_limiter_0 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_1_valid_out),
	.i_stall(bb_2_stall_out_1),
	.i_valid_exit(bb_4_valid_out_0),
	.i_stall_exit(bb_5_stall_out),
	.o_valid(loop_limiter_0_valid_out),
	.o_stall(loop_limiter_0_stall_out)
);

defparam loop_limiter_0.ENTRY_WIDTH = 1;
defparam loop_limiter_0.EXIT_WIDTH = 1;
defparam loop_limiter_0.THRESHOLD = 408;

acl_loop_limiter loop_limiter_1 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_2_valid_out),
	.i_stall(bb_3_stall_out_1),
	.i_valid_exit(bb_3_valid_out_0),
	.i_stall_exit(bb_4_stall_out),
	.o_valid(loop_limiter_1_valid_out),
	.o_stall(loop_limiter_1_stall_out)
);

defparam loop_limiter_1.ENTRY_WIDTH = 1;
defparam loop_limiter_1.EXIT_WIDTH = 1;
defparam loop_limiter_1.THRESHOLD = 400;

AOCbilateralFilterkernel_sys_cycle_time system_cycle_time_module (
	.clock(clock),
	.resetn(resetn),
	.cur_cycle(cur_cycle)
);


assign valid_out = bb_5_valid_out;
assign output_0 = bb_5_lvb_input_acl_hw_wg_id;
assign stall_out = bb_0_stall_out;
assign writes_pending = bb_5_local_bb5_st_c0_exe112_active;
assign lsus_active[0] = bb_1_local_bb1_ld__active;
assign lsus_active[1] = bb_3_local_bb3_ld__active;
assign lsus_active[2] = bb_3_local_bb3_ld__u12_active;
assign lsus_active[3] = bb_3_local_bb3_ld__u13_active;
assign lsus_active[4] = bb_5_local_bb5_st_c0_exe112_active;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		has_a_write_pending <= 1'b0;
		has_a_lsu_active <= 1'b0;
	end
	else
	begin
		has_a_write_pending <= (|writes_pending);
		has_a_lsu_active <= (|lsus_active);
	end
end

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_function_wrapper
	(
		input 		clock,
		input 		resetn,
		input 		clock2x,
		input 		local_router_hang,
		input 		avs_cra_read,
		input 		avs_cra_write,
		input [4:0] 		avs_cra_address,
		input [63:0] 		avs_cra_writedata,
		input [7:0] 		avs_cra_byteenable,
		output reg [63:0] 		avs_cra_readdata,
		output reg 		avs_cra_readdatavalid,
		output 		cra_irq,
		input [511:0] 		avm_local_bb1_ld__inst0_readdata,
		input 		avm_local_bb1_ld__inst0_readdatavalid,
		input 		avm_local_bb1_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb1_ld__inst0_address,
		output 		avm_local_bb1_ld__inst0_read,
		output 		avm_local_bb1_ld__inst0_write,
		input 		avm_local_bb1_ld__inst0_writeack,
		output [511:0] 		avm_local_bb1_ld__inst0_writedata,
		output [63:0] 		avm_local_bb1_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb1_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb3_ld__inst0_readdata,
		input 		avm_local_bb3_ld__inst0_readdatavalid,
		input 		avm_local_bb3_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb3_ld__inst0_address,
		output 		avm_local_bb3_ld__inst0_read,
		output 		avm_local_bb3_ld__inst0_write,
		input 		avm_local_bb3_ld__inst0_writeack,
		output [511:0] 		avm_local_bb3_ld__inst0_writedata,
		output [63:0] 		avm_local_bb3_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb3_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb3_ld__u12_inst0_readdata,
		input 		avm_local_bb3_ld__u12_inst0_readdatavalid,
		input 		avm_local_bb3_ld__u12_inst0_waitrequest,
		output [32:0] 		avm_local_bb3_ld__u12_inst0_address,
		output 		avm_local_bb3_ld__u12_inst0_read,
		output 		avm_local_bb3_ld__u12_inst0_write,
		input 		avm_local_bb3_ld__u12_inst0_writeack,
		output [511:0] 		avm_local_bb3_ld__u12_inst0_writedata,
		output [63:0] 		avm_local_bb3_ld__u12_inst0_byteenable,
		output [4:0] 		avm_local_bb3_ld__u12_inst0_burstcount,
		input [511:0] 		avm_local_bb3_ld__u13_inst0_readdata,
		input 		avm_local_bb3_ld__u13_inst0_readdatavalid,
		input 		avm_local_bb3_ld__u13_inst0_waitrequest,
		output [32:0] 		avm_local_bb3_ld__u13_inst0_address,
		output 		avm_local_bb3_ld__u13_inst0_read,
		output 		avm_local_bb3_ld__u13_inst0_write,
		input 		avm_local_bb3_ld__u13_inst0_writeack,
		output [511:0] 		avm_local_bb3_ld__u13_inst0_writedata,
		output [63:0] 		avm_local_bb3_ld__u13_inst0_byteenable,
		output [4:0] 		avm_local_bb3_ld__u13_inst0_burstcount,
		input [511:0] 		avm_local_bb5_st_c0_exe112_inst0_readdata,
		input 		avm_local_bb5_st_c0_exe112_inst0_readdatavalid,
		input 		avm_local_bb5_st_c0_exe112_inst0_waitrequest,
		output [32:0] 		avm_local_bb5_st_c0_exe112_inst0_address,
		output 		avm_local_bb5_st_c0_exe112_inst0_read,
		output 		avm_local_bb5_st_c0_exe112_inst0_write,
		input 		avm_local_bb5_st_c0_exe112_inst0_writeack,
		output [511:0] 		avm_local_bb5_st_c0_exe112_inst0_writedata,
		output [63:0] 		avm_local_bb5_st_c0_exe112_inst0_byteenable,
		output [4:0] 		avm_local_bb5_st_c0_exe112_inst0_burstcount
	);

// Responsible for interfacing a kernel with the outside world. It comprises a
// slave interface to specify the kernel arguments and retain kernel status. 

// This section of the wrapper implements the slave interface.
// twoXclock_consumer uses clock2x, even if nobody inside the kernel does. Keeps interface to acl_iface consistent for all kernels.
 reg start_NO_SHIFT_REG;
 reg started_NO_SHIFT_REG;
wire finish;
 reg [31:0] status_NO_SHIFT_REG;
wire has_a_write_pending;
wire has_a_lsu_active;
 reg [255:0] kernel_arguments_NO_SHIFT_REG;
 reg twoXclock_consumer_NO_SHIFT_REG /* synthesis  preserve  noprune  */;
 reg [31:0] workgroup_size_NO_SHIFT_REG;
 reg [31:0] global_size_NO_SHIFT_REG[2:0];
 reg [31:0] num_groups_NO_SHIFT_REG[2:0];
 reg [31:0] local_size_NO_SHIFT_REG[2:0];
 reg [31:0] work_dim_NO_SHIFT_REG;
 reg [31:0] global_offset_NO_SHIFT_REG[2:0];
 reg [63:0] profile_data_NO_SHIFT_REG;
 reg [31:0] profile_ctrl_NO_SHIFT_REG;
 reg [63:0] profile_start_cycle_NO_SHIFT_REG;
 reg [63:0] profile_stop_cycle_NO_SHIFT_REG;
wire dispatched_all_groups;
wire [31:0] group_id_tmp[2:0];
wire [31:0] global_id_base_out[2:0];
wire start_out;
wire [31:0] local_id[0:0][2:0];
wire [31:0] global_id[0:0][2:0];
wire [31:0] group_id[0:0][2:0];
wire iter_valid_in;
wire iter_stall_out;
wire stall_in;
wire stall_out;
wire valid_in;
wire valid_out;

always @(posedge clock2x or negedge resetn)
begin
	if (~(resetn))
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b1;
	end
end



// Work group dispatcher is responsible for issuing work-groups to id iterator(s)
acl_work_group_dispatcher group_dispatcher (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.num_groups(num_groups_NO_SHIFT_REG),
	.local_size(local_size_NO_SHIFT_REG),
	.stall_in(iter_stall_out),
	.valid_out(iter_valid_in),
	.group_id_out(group_id_tmp),
	.global_id_base_out(global_id_base_out),
	.start_out(start_out),
	.dispatched_all_groups(dispatched_all_groups)
);

defparam group_dispatcher.NUM_COPIES = 1;
defparam group_dispatcher.RUN_FOREVER = 0;


// This section of the wrapper implements an Avalon Slave Interface used to configure a kernel invocation.
// The few words words contain the status and the workgroup size registers.
// The remaining addressable space is reserved for kernel arguments.
 reg [63:0] cra_readdata_st1_NO_SHIFT_REG;
 reg [4:0] cra_addr_st1_NO_SHIFT_REG;
 reg cra_read_st1_NO_SHIFT_REG;
wire [63:0] bitenable;

assign bitenable[7:0] = (avs_cra_byteenable[0] ? 8'hFF : 8'h0);
assign bitenable[15:8] = (avs_cra_byteenable[1] ? 8'hFF : 8'h0);
assign bitenable[23:16] = (avs_cra_byteenable[2] ? 8'hFF : 8'h0);
assign bitenable[31:24] = (avs_cra_byteenable[3] ? 8'hFF : 8'h0);
assign bitenable[39:32] = (avs_cra_byteenable[4] ? 8'hFF : 8'h0);
assign bitenable[47:40] = (avs_cra_byteenable[5] ? 8'hFF : 8'h0);
assign bitenable[55:48] = (avs_cra_byteenable[6] ? 8'hFF : 8'h0);
assign bitenable[63:56] = (avs_cra_byteenable[7] ? 8'hFF : 8'h0);
assign cra_irq = (status_NO_SHIFT_REG[1] | status_NO_SHIFT_REG[3]);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		start_NO_SHIFT_REG <= 1'b0;
		started_NO_SHIFT_REG <= 1'b0;
		kernel_arguments_NO_SHIFT_REG <= 256'h0;
		status_NO_SHIFT_REG <= 32'h30000;
		profile_ctrl_NO_SHIFT_REG <= 32'h4;
		profile_start_cycle_NO_SHIFT_REG <= 64'h0;
		profile_stop_cycle_NO_SHIFT_REG <= 64'hFFFFFFFFFFFFFFFF;
		work_dim_NO_SHIFT_REG <= 32'h0;
		workgroup_size_NO_SHIFT_REG <= 32'h0;
		global_size_NO_SHIFT_REG[0] <= 32'h0;
		global_size_NO_SHIFT_REG[1] <= 32'h0;
		global_size_NO_SHIFT_REG[2] <= 32'h0;
		num_groups_NO_SHIFT_REG[0] <= 32'h0;
		num_groups_NO_SHIFT_REG[1] <= 32'h0;
		num_groups_NO_SHIFT_REG[2] <= 32'h0;
		local_size_NO_SHIFT_REG[0] <= 32'h0;
		local_size_NO_SHIFT_REG[1] <= 32'h0;
		local_size_NO_SHIFT_REG[2] <= 32'h0;
		global_offset_NO_SHIFT_REG[0] <= 32'h0;
		global_offset_NO_SHIFT_REG[1] <= 32'h0;
		global_offset_NO_SHIFT_REG[2] <= 32'h0;
	end
	else
	begin
		if (avs_cra_write)
		begin
			case (avs_cra_address)
				5'h0:
				begin
					status_NO_SHIFT_REG[31:16] <= 16'h3;
					status_NO_SHIFT_REG[15:0] <= ((status_NO_SHIFT_REG[15:0] & ~(bitenable[15:0])) | (avs_cra_writedata[15:0] & bitenable[15:0]));
				end

				5'h1:
				begin
					profile_ctrl_NO_SHIFT_REG <= ((profile_ctrl_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h3:
				begin
					profile_start_cycle_NO_SHIFT_REG[31:0] <= ((profile_start_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_start_cycle_NO_SHIFT_REG[63:32] <= ((profile_start_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h4:
				begin
					profile_stop_cycle_NO_SHIFT_REG[31:0] <= ((profile_stop_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_stop_cycle_NO_SHIFT_REG[63:32] <= ((profile_stop_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h5:
				begin
					work_dim_NO_SHIFT_REG <= ((work_dim_NO_SHIFT_REG & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					workgroup_size_NO_SHIFT_REG <= ((workgroup_size_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h6:
				begin
					global_size_NO_SHIFT_REG[0] <= ((global_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_size_NO_SHIFT_REG[1] <= ((global_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h7:
				begin
					global_size_NO_SHIFT_REG[2] <= ((global_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[0] <= ((num_groups_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h8:
				begin
					num_groups_NO_SHIFT_REG[1] <= ((num_groups_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[2] <= ((num_groups_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h9:
				begin
					local_size_NO_SHIFT_REG[0] <= ((local_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					local_size_NO_SHIFT_REG[1] <= ((local_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hA:
				begin
					local_size_NO_SHIFT_REG[2] <= ((local_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[0] <= ((global_offset_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hB:
				begin
					global_offset_NO_SHIFT_REG[1] <= ((global_offset_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[2] <= ((global_offset_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hC:
				begin
					kernel_arguments_NO_SHIFT_REG[31:0] <= ((kernel_arguments_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[63:32] <= ((kernel_arguments_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hD:
				begin
					kernel_arguments_NO_SHIFT_REG[95:64] <= ((kernel_arguments_NO_SHIFT_REG[95:64] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[127:96] <= ((kernel_arguments_NO_SHIFT_REG[127:96] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hE:
				begin
					kernel_arguments_NO_SHIFT_REG[159:128] <= ((kernel_arguments_NO_SHIFT_REG[159:128] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[191:160] <= ((kernel_arguments_NO_SHIFT_REG[191:160] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hF:
				begin
					kernel_arguments_NO_SHIFT_REG[223:192] <= ((kernel_arguments_NO_SHIFT_REG[223:192] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[255:224] <= ((kernel_arguments_NO_SHIFT_REG[255:224] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				default:
				begin
				end

			endcase
		end
		else
		begin
			if (status_NO_SHIFT_REG[0])
			begin
				start_NO_SHIFT_REG <= 1'b1;
			end
			if (start_NO_SHIFT_REG)
			begin
				status_NO_SHIFT_REG[0] <= 1'b0;
				started_NO_SHIFT_REG <= 1'b1;
			end
			if (started_NO_SHIFT_REG)
			begin
				start_NO_SHIFT_REG <= 1'b0;
			end
			if (finish)
			begin
				status_NO_SHIFT_REG[1] <= 1'b1;
				started_NO_SHIFT_REG <= 1'b0;
			end
		end
		status_NO_SHIFT_REG[11] <= 1'b0;
		status_NO_SHIFT_REG[12] <= (|has_a_lsu_active);
		status_NO_SHIFT_REG[13] <= (|has_a_write_pending);
		status_NO_SHIFT_REG[14] <= (|valid_in);
		status_NO_SHIFT_REG[15] <= started_NO_SHIFT_REG;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cra_read_st1_NO_SHIFT_REG <= 1'b0;
		cra_addr_st1_NO_SHIFT_REG <= 5'h0;
		cra_readdata_st1_NO_SHIFT_REG <= 64'h0;
	end
	else
	begin
		cra_read_st1_NO_SHIFT_REG <= avs_cra_read;
		cra_addr_st1_NO_SHIFT_REG <= avs_cra_address;
		case (avs_cra_address)
			5'h0:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= status_NO_SHIFT_REG;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			5'h1:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= 'x;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			5'h2:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			5'h3:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			5'h4:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			default:
			begin
				cra_readdata_st1_NO_SHIFT_REG <= status_NO_SHIFT_REG;
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		avs_cra_readdatavalid <= 1'b0;
		avs_cra_readdata <= 64'h0;
	end
	else
	begin
		avs_cra_readdatavalid <= cra_read_st1_NO_SHIFT_REG;
		case (cra_addr_st1_NO_SHIFT_REG)
			5'h2:
			begin
				avs_cra_readdata[63:0] <= profile_data_NO_SHIFT_REG;
			end

			default:
			begin
				avs_cra_readdata <= cra_readdata_st1_NO_SHIFT_REG;
			end

		endcase
	end
end


// Handshaking signals used to control data through the pipeline

// Determine when the kernel is finished.
acl_kernel_finish_detector kernel_finish_detector (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.wg_size(workgroup_size_NO_SHIFT_REG),
	.wg_dispatch_valid_out(iter_valid_in),
	.wg_dispatch_stall_in(iter_stall_out),
	.dispatched_all_groups(dispatched_all_groups),
	.kernel_copy_valid_out(valid_out),
	.kernel_copy_stall_in(stall_in),
	.pending_writes(has_a_write_pending),
	.finish(finish)
);

defparam kernel_finish_detector.TESSELLATION_SIZE = 0;
defparam kernel_finish_detector.NUM_COPIES = 1;
defparam kernel_finish_detector.WG_SIZE_W = 32;

assign stall_in = 1'b0;

// Creating ID iterator and kernel instance for every requested kernel copy

// ID iterator is responsible for iterating over all local ids for given work-groups
acl_id_iterator id_iter_inst0 (
	.clock(clock),
	.resetn(resetn),
	.start(start_out),
	.valid_in(iter_valid_in),
	.stall_out(iter_stall_out),
	.stall_in(stall_out),
	.valid_out(valid_in),
	.group_id_in(group_id_tmp),
	.global_id_base_in(global_id_base_out),
	.local_size(local_size_NO_SHIFT_REG),
	.global_size(global_size_NO_SHIFT_REG),
	.local_id(local_id[0]),
	.global_id(global_id[0]),
	.group_id(group_id[0])
);



// This section instantiates a kernel function block
AOCbilateralFilterkernel_function AOCbilateralFilterkernel_function_inst0 (
	.clock(clock),
	.resetn(resetn),
	.input_global_id_0(global_id[0][0]),
	.input_global_id_1(global_id[0][1]),
	.input_acl_hw_wg_id(),
	.stall_out(stall_out),
	.valid_in(valid_in),
	.output_0(),
	.valid_out(valid_out),
	.stall_in(stall_in),
	.workgroup_size(workgroup_size_NO_SHIFT_REG),
	.avm_local_bb1_ld__readdata(avm_local_bb1_ld__inst0_readdata),
	.avm_local_bb1_ld__readdatavalid(avm_local_bb1_ld__inst0_readdatavalid),
	.avm_local_bb1_ld__waitrequest(avm_local_bb1_ld__inst0_waitrequest),
	.avm_local_bb1_ld__address(avm_local_bb1_ld__inst0_address),
	.avm_local_bb1_ld__read(avm_local_bb1_ld__inst0_read),
	.avm_local_bb1_ld__write(avm_local_bb1_ld__inst0_write),
	.avm_local_bb1_ld__writeack(avm_local_bb1_ld__inst0_writeack),
	.avm_local_bb1_ld__writedata(avm_local_bb1_ld__inst0_writedata),
	.avm_local_bb1_ld__byteenable(avm_local_bb1_ld__inst0_byteenable),
	.avm_local_bb1_ld__burstcount(avm_local_bb1_ld__inst0_burstcount),
	.avm_local_bb3_ld__readdata(avm_local_bb3_ld__inst0_readdata),
	.avm_local_bb3_ld__readdatavalid(avm_local_bb3_ld__inst0_readdatavalid),
	.avm_local_bb3_ld__waitrequest(avm_local_bb3_ld__inst0_waitrequest),
	.avm_local_bb3_ld__address(avm_local_bb3_ld__inst0_address),
	.avm_local_bb3_ld__read(avm_local_bb3_ld__inst0_read),
	.avm_local_bb3_ld__write(avm_local_bb3_ld__inst0_write),
	.avm_local_bb3_ld__writeack(avm_local_bb3_ld__inst0_writeack),
	.avm_local_bb3_ld__writedata(avm_local_bb3_ld__inst0_writedata),
	.avm_local_bb3_ld__byteenable(avm_local_bb3_ld__inst0_byteenable),
	.avm_local_bb3_ld__burstcount(avm_local_bb3_ld__inst0_burstcount),
	.avm_local_bb3_ld__u12_readdata(avm_local_bb3_ld__u12_inst0_readdata),
	.avm_local_bb3_ld__u12_readdatavalid(avm_local_bb3_ld__u12_inst0_readdatavalid),
	.avm_local_bb3_ld__u12_waitrequest(avm_local_bb3_ld__u12_inst0_waitrequest),
	.avm_local_bb3_ld__u12_address(avm_local_bb3_ld__u12_inst0_address),
	.avm_local_bb3_ld__u12_read(avm_local_bb3_ld__u12_inst0_read),
	.avm_local_bb3_ld__u12_write(avm_local_bb3_ld__u12_inst0_write),
	.avm_local_bb3_ld__u12_writeack(avm_local_bb3_ld__u12_inst0_writeack),
	.avm_local_bb3_ld__u12_writedata(avm_local_bb3_ld__u12_inst0_writedata),
	.avm_local_bb3_ld__u12_byteenable(avm_local_bb3_ld__u12_inst0_byteenable),
	.avm_local_bb3_ld__u12_burstcount(avm_local_bb3_ld__u12_inst0_burstcount),
	.avm_local_bb3_ld__u13_readdata(avm_local_bb3_ld__u13_inst0_readdata),
	.avm_local_bb3_ld__u13_readdatavalid(avm_local_bb3_ld__u13_inst0_readdatavalid),
	.avm_local_bb3_ld__u13_waitrequest(avm_local_bb3_ld__u13_inst0_waitrequest),
	.avm_local_bb3_ld__u13_address(avm_local_bb3_ld__u13_inst0_address),
	.avm_local_bb3_ld__u13_read(avm_local_bb3_ld__u13_inst0_read),
	.avm_local_bb3_ld__u13_write(avm_local_bb3_ld__u13_inst0_write),
	.avm_local_bb3_ld__u13_writeack(avm_local_bb3_ld__u13_inst0_writeack),
	.avm_local_bb3_ld__u13_writedata(avm_local_bb3_ld__u13_inst0_writedata),
	.avm_local_bb3_ld__u13_byteenable(avm_local_bb3_ld__u13_inst0_byteenable),
	.avm_local_bb3_ld__u13_burstcount(avm_local_bb3_ld__u13_inst0_burstcount),
	.avm_local_bb5_st_c0_exe112_readdata(avm_local_bb5_st_c0_exe112_inst0_readdata),
	.avm_local_bb5_st_c0_exe112_readdatavalid(avm_local_bb5_st_c0_exe112_inst0_readdatavalid),
	.avm_local_bb5_st_c0_exe112_waitrequest(avm_local_bb5_st_c0_exe112_inst0_waitrequest),
	.avm_local_bb5_st_c0_exe112_address(avm_local_bb5_st_c0_exe112_inst0_address),
	.avm_local_bb5_st_c0_exe112_read(avm_local_bb5_st_c0_exe112_inst0_read),
	.avm_local_bb5_st_c0_exe112_write(avm_local_bb5_st_c0_exe112_inst0_write),
	.avm_local_bb5_st_c0_exe112_writeack(avm_local_bb5_st_c0_exe112_inst0_writeack),
	.avm_local_bb5_st_c0_exe112_writedata(avm_local_bb5_st_c0_exe112_inst0_writedata),
	.avm_local_bb5_st_c0_exe112_byteenable(avm_local_bb5_st_c0_exe112_inst0_byteenable),
	.avm_local_bb5_st_c0_exe112_burstcount(avm_local_bb5_st_c0_exe112_inst0_burstcount),
	.start(start_out),
	.input_r(kernel_arguments_NO_SHIFT_REG[255:224]),
	.input_global_size_0(global_size_NO_SHIFT_REG[0]),
	.input_global_size_1(global_size_NO_SHIFT_REG[1]),
	.input_e_d(kernel_arguments_NO_SHIFT_REG[223:192]),
	.clock2x(clock2x),
	.input_in(kernel_arguments_NO_SHIFT_REG[127:64]),
	.input_gaussian(kernel_arguments_NO_SHIFT_REG[191:128]),
	.input_out(kernel_arguments_NO_SHIFT_REG[63:0]),
	.has_a_write_pending(has_a_write_pending),
	.has_a_lsu_active(has_a_lsu_active)
);



endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_sys_cycle_time
	(
		input 		clock,
		input 		resetn,
		output [31:0] 		cur_cycle
	);


 reg [31:0] cur_count_NO_SHIFT_REG;

assign cur_cycle = cur_count_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cur_count_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		cur_count_NO_SHIFT_REG <= (cur_count_NO_SHIFT_REG + 32'h1);
	end
end

endmodule

