// (C) 1992-2015 Altera Corporation. All rights reserved.                         
// Your use of Altera Corporation's design tools, logic functions and other       
// software and tools, and its AMPP partner logic functions, and any output       
// files any of the foregoing (including device programming or simulation         
// files), and any associated documentation or information are expressly subject  
// to the terms and conditions of the Altera Program License Subscription         
// Agreement, Altera MegaCore Function License Agreement, or other applicable     
// license agreement, including, without limitation, that your use is for the     
// sole purpose of programming logic devices manufactured by Altera and sold by   
// Altera or its authorized distributors.  Please refer to the applicable         
// agreement for further details.                                                 
    

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_0
	(
		input 		clock,
		input 		resetn,
		input 		start,
		input [31:0] 		input_r,
		input [31:0] 		input_e_d,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out,
		input 		stall_in,
		output 		lvb_bb0_cmp1017,
		output [31:0] 		lvb_bb0_mul39,
		output [63:0] 		lvb_bb0_var_,
		output [63:0] 		lvb_bb0_var__u0,
		input [31:0] 		workgroup_size
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub_inputs_ready;
 reg local_bb0_sub_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub_valid_out_0_NO_SHIFT_REG;
wire local_bb0_sub_stall_in_0;
 reg local_bb0_sub_valid_out_1_NO_SHIFT_REG;
wire local_bb0_sub_stall_in_1;
wire local_bb0_sub_output_regs_ready;
 reg [31:0] local_bb0_sub_NO_SHIFT_REG;
wire local_bb0_sub_causedstall;

assign local_bb0_sub_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb0_sub_output_regs_ready = (~(local_bb0_sub_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_sub_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_sub_stall_in_0)) & (~(local_bb0_sub_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_sub_stall_in_1))));
assign merge_node_stall_in_0 = (~(local_bb0_sub_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub_output_regs_ready) | ~(local_bb0_sub_inputs_ready)));
assign local_bb0_sub_causedstall = (local_bb0_sub_inputs_ready && (~(local_bb0_sub_output_regs_ready) && !(~(local_bb0_sub_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub_NO_SHIFT_REG <= 'x;
		local_bb0_sub_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_sub_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub_NO_SHIFT_REG <= 'x;
			local_bb0_sub_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_sub_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub_output_regs_ready)
			begin
				local_bb0_sub_NO_SHIFT_REG <= (32'h0 - input_r);
				local_bb0_sub_valid_out_0_NO_SHIFT_REG <= local_bb0_sub_inputs_ready;
				local_bb0_sub_valid_out_1_NO_SHIFT_REG <= local_bb0_sub_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub_stall_in_0))
				begin
					local_bb0_sub_valid_out_0_NO_SHIFT_REG <= local_bb0_sub_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_sub_stall_in_1))
				begin
					local_bb0_sub_valid_out_1_NO_SHIFT_REG <= local_bb0_sub_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub_inputs_ready)
			begin
				local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u1_inputs_ready;
 reg local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u1_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u1_stall_in;
wire local_bb0_var__u1_output_regs_ready;
 reg [31:0] local_bb0_var__u1_NO_SHIFT_REG;
wire local_bb0_var__u1_causedstall;

assign local_bb0_var__u1_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign local_bb0_var__u1_output_regs_ready = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u1_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u1_stall_in))));
assign merge_node_stall_in_2 = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u1_output_regs_ready) | ~(local_bb0_var__u1_inputs_ready)));
assign local_bb0_var__u1_causedstall = (local_bb0_var__u1_inputs_ready && (~(local_bb0_var__u1_output_regs_ready) && !(~(local_bb0_var__u1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_NO_SHIFT_REG <= 'x;
		local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_NO_SHIFT_REG <= 'x;
			local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_output_regs_ready)
			begin
				local_bb0_var__u1_NO_SHIFT_REG <= input_e_d;
				local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u1_stall_in))
				begin
					local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_inputs_ready)
			begin
				local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u0_inputs_ready;
 reg local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u0_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u0_stall_in;
wire local_bb0_var__u0_output_regs_ready;
 reg [63:0] local_bb0_var__u0_NO_SHIFT_REG;
wire local_bb0_var__u0_causedstall;

assign local_bb0_var__u0_inputs_ready = merge_node_valid_out_4_NO_SHIFT_REG;
assign local_bb0_var__u0_output_regs_ready = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u0_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u0_stall_in))));
assign merge_node_stall_in_4 = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u0_output_regs_ready) | ~(local_bb0_var__u0_inputs_ready)));
assign local_bb0_var__u0_causedstall = (local_bb0_var__u0_inputs_ready && (~(local_bb0_var__u0_output_regs_ready) && !(~(local_bb0_var__u0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_NO_SHIFT_REG <= 'x;
		local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_NO_SHIFT_REG <= 'x;
			local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_output_regs_ready)
			begin
				local_bb0_var__u0_NO_SHIFT_REG <= $signed(input_r);
				local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u0_stall_in))
				begin
					local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_inputs_ready)
			begin
				local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp1017_inputs_ready;
 reg local_bb0_cmp1017_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp1017_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp1017_stall_in;
wire local_bb0_cmp1017_output_regs_ready;
 reg local_bb0_cmp1017_NO_SHIFT_REG;
wire local_bb0_cmp1017_causedstall;

assign local_bb0_cmp1017_inputs_ready = (local_bb0_sub_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign local_bb0_cmp1017_output_regs_ready = (~(local_bb0_cmp1017_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp1017_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp1017_stall_in))));
assign local_bb0_sub_stall_in_0 = (~(local_bb0_cmp1017_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp1017_output_regs_ready) | ~(local_bb0_cmp1017_inputs_ready)));
assign merge_node_stall_in_1 = (~(local_bb0_cmp1017_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp1017_output_regs_ready) | ~(local_bb0_cmp1017_inputs_ready)));
assign local_bb0_cmp1017_causedstall = (local_bb0_cmp1017_inputs_ready && (~(local_bb0_cmp1017_output_regs_ready) && !(~(local_bb0_cmp1017_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp1017_NO_SHIFT_REG <= 'x;
		local_bb0_cmp1017_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp1017_NO_SHIFT_REG <= 'x;
			local_bb0_cmp1017_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp1017_output_regs_ready)
			begin
				local_bb0_cmp1017_NO_SHIFT_REG <= ($signed(local_bb0_sub_NO_SHIFT_REG) > $signed(input_r));
				local_bb0_cmp1017_valid_out_NO_SHIFT_REG <= local_bb0_cmp1017_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp1017_stall_in))
				begin
					local_bb0_cmp1017_valid_out_NO_SHIFT_REG <= local_bb0_cmp1017_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp1017_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp1017_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp1017_inputs_ready)
			begin
				local_bb0_cmp1017_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__inputs_ready;
 reg local_bb0_var__wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__valid_out_NO_SHIFT_REG;
wire local_bb0_var__stall_in;
wire local_bb0_var__output_regs_ready;
 reg [63:0] local_bb0_var__NO_SHIFT_REG;
wire local_bb0_var__causedstall;

assign local_bb0_var__inputs_ready = local_bb0_sub_valid_out_1_NO_SHIFT_REG;
assign local_bb0_var__output_regs_ready = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__valid_out_NO_SHIFT_REG) | ~(local_bb0_var__stall_in))));
assign local_bb0_sub_stall_in_1 = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__output_regs_ready) | ~(local_bb0_var__inputs_ready)));
assign local_bb0_var__causedstall = (local_bb0_var__inputs_ready && (~(local_bb0_var__output_regs_ready) && !(~(local_bb0_var__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__NO_SHIFT_REG <= 'x;
		local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__NO_SHIFT_REG <= 'x;
			local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__output_regs_ready)
			begin
				local_bb0_var__NO_SHIFT_REG <= $signed(local_bb0_sub_NO_SHIFT_REG);
				local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__stall_in))
				begin
					local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__inputs_ready)
			begin
				local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_2to2_bb0_var__u1_valid_out_0;
wire rstag_2to2_bb0_var__u1_stall_in_0;
wire rstag_2to2_bb0_var__u1_valid_out_1;
wire rstag_2to2_bb0_var__u1_stall_in_1;
wire rstag_2to2_bb0_var__u1_valid_out_2;
wire rstag_2to2_bb0_var__u1_stall_in_2;
wire rstag_2to2_bb0_var__u1_inputs_ready;
wire rstag_2to2_bb0_var__u1_stall_local;
 reg rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG;
wire rstag_2to2_bb0_var__u1_combined_valid;
 reg [31:0] rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_2to2_bb0_var__u1;
 reg rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG;
 reg rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG;
 reg rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG;

assign rstag_2to2_bb0_var__u1_inputs_ready = local_bb0_var__u1_valid_out_NO_SHIFT_REG;
assign rstag_2to2_bb0_var__u1 = (rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG ? rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG : local_bb0_var__u1_NO_SHIFT_REG);
assign rstag_2to2_bb0_var__u1_combined_valid = (rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG | rstag_2to2_bb0_var__u1_inputs_ready);
assign rstag_2to2_bb0_var__u1_stall_local = ((rstag_2to2_bb0_var__u1_stall_in_0 & ~(rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG)) | (rstag_2to2_bb0_var__u1_stall_in_1 & ~(rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG)) | (rstag_2to2_bb0_var__u1_stall_in_2 & ~(rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG)));
assign rstag_2to2_bb0_var__u1_valid_out_0 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG));
assign rstag_2to2_bb0_var__u1_valid_out_1 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG));
assign rstag_2to2_bb0_var__u1_valid_out_2 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG));
assign local_bb0_var__u1_stall_in = (|rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_2to2_bb0_var__u1_stall_local)
			begin
				if (~(rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG))
				begin
					rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= rstag_2to2_bb0_var__u1_inputs_ready;
				end
			end
			else
			begin
				rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG))
		begin
			rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG <= local_bb0_var__u1_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_0)) & rstag_2to2_bb0_var__u1_stall_local);
			rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_1)) & rstag_2to2_bb0_var__u1_stall_local);
			rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_2)) & rstag_2to2_bb0_var__u1_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and33_i_inputs_ready;
 reg local_bb0_and33_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and33_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and33_i_stall_in;
wire local_bb0_and33_i_output_regs_ready;
 reg [31:0] local_bb0_and33_i_NO_SHIFT_REG;
wire local_bb0_and33_i_causedstall;

assign local_bb0_and33_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_0;
assign local_bb0_and33_i_output_regs_ready = (~(local_bb0_and33_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and33_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and33_i_stall_in))));
assign rstag_2to2_bb0_var__u1_stall_in_0 = (~(local_bb0_and33_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and33_i_output_regs_ready) | ~(local_bb0_and33_i_inputs_ready)));
assign local_bb0_and33_i_causedstall = (local_bb0_and33_i_inputs_ready && (~(local_bb0_and33_i_output_regs_ready) && !(~(local_bb0_and33_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and33_i_NO_SHIFT_REG <= 'x;
		local_bb0_and33_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and33_i_NO_SHIFT_REG <= 'x;
			local_bb0_and33_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and33_i_output_regs_ready)
			begin
				local_bb0_and33_i_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1 & 32'h807FFFFF);
				local_bb0_and33_i_valid_out_NO_SHIFT_REG <= local_bb0_and33_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and33_i_stall_in))
				begin
					local_bb0_and33_i_valid_out_NO_SHIFT_REG <= local_bb0_and33_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and33_i_inputs_ready)
			begin
				local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_and2_i_valid_out;
wire local_bb0_and2_i_stall_in;
wire local_bb0_and2_i_inputs_ready;
wire local_bb0_and2_i_stall_local;
wire [31:0] local_bb0_and2_i;

assign local_bb0_and2_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_1;
assign local_bb0_and2_i = (rstag_2to2_bb0_var__u1 & 32'h7FFFFF);
assign local_bb0_and2_i_valid_out = local_bb0_and2_i_inputs_ready;
assign local_bb0_and2_i_stall_local = local_bb0_and2_i_stall_in;
assign rstag_2to2_bb0_var__u1_stall_in_1 = (|local_bb0_and2_i_stall_local);

// This section implements a registered operation.
// 
wire local_bb0_shr_i_inputs_ready;
 reg local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_shr_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_shr_i_stall_in_0;
 reg local_bb0_shr_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_shr_i_stall_in_1;
wire local_bb0_shr_i_output_regs_ready;
 reg [31:0] local_bb0_shr_i_NO_SHIFT_REG;
wire local_bb0_shr_i_causedstall;

assign local_bb0_shr_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_2;
assign local_bb0_shr_i_output_regs_ready = (~(local_bb0_shr_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_shr_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_shr_i_stall_in_0)) & (~(local_bb0_shr_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_shr_i_stall_in_1))));
assign rstag_2to2_bb0_var__u1_stall_in_2 = (~(local_bb0_shr_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_shr_i_output_regs_ready) | ~(local_bb0_shr_i_inputs_ready)));
assign local_bb0_shr_i_causedstall = (local_bb0_shr_i_inputs_ready && (~(local_bb0_shr_i_output_regs_ready) && !(~(local_bb0_shr_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_shr_i_NO_SHIFT_REG <= 'x;
		local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_shr_i_NO_SHIFT_REG <= 'x;
			local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_shr_i_output_regs_ready)
			begin
				local_bb0_shr_i_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1 >> 32'h17);
				local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= local_bb0_shr_i_inputs_ready;
				local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= local_bb0_shr_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_shr_i_stall_in_0))
				begin
					local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_shr_i_stall_in_1))
				begin
					local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_shr_i_inputs_ready)
			begin
				local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_lnot6_i_inputs_ready;
 reg local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_lnot6_i_valid_out_NO_SHIFT_REG;
wire local_bb0_lnot6_i_stall_in;
wire local_bb0_lnot6_i_output_regs_ready;
 reg local_bb0_lnot6_i_NO_SHIFT_REG;
wire local_bb0_lnot6_i_causedstall;

assign local_bb0_lnot6_i_inputs_ready = local_bb0_and2_i_valid_out;
assign local_bb0_lnot6_i_output_regs_ready = (~(local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_lnot6_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_lnot6_i_stall_in))));
assign local_bb0_and2_i_stall_in = (~(local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_lnot6_i_output_regs_ready) | ~(local_bb0_lnot6_i_inputs_ready)));
assign local_bb0_lnot6_i_causedstall = (local_bb0_lnot6_i_inputs_ready && (~(local_bb0_lnot6_i_output_regs_ready) && !(~(local_bb0_lnot6_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_lnot6_i_NO_SHIFT_REG <= 'x;
		local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_lnot6_i_NO_SHIFT_REG <= 'x;
			local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_lnot6_i_output_regs_ready)
			begin
				local_bb0_lnot6_i_NO_SHIFT_REG <= ((local_bb0_and2_i & 32'h7FFFFF) != 32'h0);
				local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= local_bb0_lnot6_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_lnot6_i_stall_in))
				begin
					local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_lnot6_i_inputs_ready)
			begin
				local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and1_i_inputs_ready;
 reg local_bb0_and1_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and1_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and1_i_stall_in;
wire local_bb0_and1_i_output_regs_ready;
 reg [31:0] local_bb0_and1_i_NO_SHIFT_REG;
wire local_bb0_and1_i_causedstall;

assign local_bb0_and1_i_inputs_ready = local_bb0_shr_i_valid_out_0_NO_SHIFT_REG;
assign local_bb0_and1_i_output_regs_ready = (~(local_bb0_and1_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and1_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and1_i_stall_in))));
assign local_bb0_shr_i_stall_in_0 = (~(local_bb0_and1_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and1_i_output_regs_ready) | ~(local_bb0_and1_i_inputs_ready)));
assign local_bb0_and1_i_causedstall = (local_bb0_and1_i_inputs_ready && (~(local_bb0_and1_i_output_regs_ready) && !(~(local_bb0_and1_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and1_i_NO_SHIFT_REG <= 'x;
		local_bb0_and1_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and1_i_NO_SHIFT_REG <= 'x;
			local_bb0_and1_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and1_i_output_regs_ready)
			begin
				local_bb0_and1_i_NO_SHIFT_REG <= ((local_bb0_shr_i_NO_SHIFT_REG & 32'h1FF) & 32'hFF);
				local_bb0_and1_i_valid_out_NO_SHIFT_REG <= local_bb0_and1_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and1_i_stall_in))
				begin
					local_bb0_and1_i_valid_out_NO_SHIFT_REG <= local_bb0_and1_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and1_i_inputs_ready)
			begin
				local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_4to4_bb0_and1_i_valid_out_0;
wire rstag_4to4_bb0_and1_i_stall_in_0;
wire rstag_4to4_bb0_and1_i_valid_out_1;
wire rstag_4to4_bb0_and1_i_stall_in_1;
wire rstag_4to4_bb0_and1_i_valid_out_2;
wire rstag_4to4_bb0_and1_i_stall_in_2;
wire rstag_4to4_bb0_and1_i_inputs_ready;
wire rstag_4to4_bb0_and1_i_stall_local;
 reg rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG;
wire rstag_4to4_bb0_and1_i_combined_valid;
 reg [31:0] rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_4to4_bb0_and1_i;
 reg rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG;
 reg rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG;
 reg rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG;

assign rstag_4to4_bb0_and1_i_inputs_ready = local_bb0_and1_i_valid_out_NO_SHIFT_REG;
assign rstag_4to4_bb0_and1_i = (rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG ? rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG : (local_bb0_and1_i_NO_SHIFT_REG & 32'hFF));
assign rstag_4to4_bb0_and1_i_combined_valid = (rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG | rstag_4to4_bb0_and1_i_inputs_ready);
assign rstag_4to4_bb0_and1_i_stall_local = ((rstag_4to4_bb0_and1_i_stall_in_0 & ~(rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG)) | (rstag_4to4_bb0_and1_i_stall_in_1 & ~(rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG)) | (rstag_4to4_bb0_and1_i_stall_in_2 & ~(rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG)));
assign rstag_4to4_bb0_and1_i_valid_out_0 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG));
assign rstag_4to4_bb0_and1_i_valid_out_1 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG));
assign rstag_4to4_bb0_and1_i_valid_out_2 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG));
assign local_bb0_and1_i_stall_in = (|rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_4to4_bb0_and1_i_stall_local)
			begin
				if (~(rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= rstag_4to4_bb0_and1_i_inputs_ready;
				end
			end
			else
			begin
				rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG <= (local_bb0_and1_i_NO_SHIFT_REG & 32'hFF);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_0)) & rstag_4to4_bb0_and1_i_stall_local);
			rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_1)) & rstag_4to4_bb0_and1_i_stall_local);
			rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_2)) & rstag_4to4_bb0_and1_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp10_i_inputs_ready;
 reg local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_cmp10_i_stall_in_0;
 reg local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_cmp10_i_stall_in_1;
wire local_bb0_cmp10_i_output_regs_ready;
 reg local_bb0_cmp10_i_NO_SHIFT_REG;
wire local_bb0_cmp10_i_causedstall;

assign local_bb0_cmp10_i_inputs_ready = rstag_4to4_bb0_and1_i_valid_out_1;
assign local_bb0_cmp10_i_output_regs_ready = (~(local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_cmp10_i_stall_in_0)) & (~(local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_cmp10_i_stall_in_1))));
assign rstag_4to4_bb0_and1_i_stall_in_1 = (~(local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp10_i_output_regs_ready) | ~(local_bb0_cmp10_i_inputs_ready)));
assign local_bb0_cmp10_i_causedstall = (local_bb0_cmp10_i_inputs_ready && (~(local_bb0_cmp10_i_output_regs_ready) && !(~(local_bb0_cmp10_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp10_i_NO_SHIFT_REG <= 'x;
		local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp10_i_NO_SHIFT_REG <= 'x;
			local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp10_i_output_regs_ready)
			begin
				local_bb0_cmp10_i_NO_SHIFT_REG <= ((rstag_4to4_bb0_and1_i & 32'hFF) == 32'h0);
				local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp10_i_inputs_ready;
				local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp10_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp10_i_stall_in_0))
				begin
					local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_cmp10_i_stall_in_1))
				begin
					local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp10_i_inputs_ready)
			begin
				local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp_i_inputs_ready;
 reg local_bb0_cmp_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp_i_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp_i_stall_in;
wire local_bb0_cmp_i_output_regs_ready;
 reg local_bb0_cmp_i_NO_SHIFT_REG;
wire local_bb0_cmp_i_causedstall;

assign local_bb0_cmp_i_inputs_ready = rstag_4to4_bb0_and1_i_valid_out_2;
assign local_bb0_cmp_i_output_regs_ready = (~(local_bb0_cmp_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp_i_stall_in))));
assign rstag_4to4_bb0_and1_i_stall_in_2 = (~(local_bb0_cmp_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp_i_output_regs_ready) | ~(local_bb0_cmp_i_inputs_ready)));
assign local_bb0_cmp_i_causedstall = (local_bb0_cmp_i_inputs_ready && (~(local_bb0_cmp_i_output_regs_ready) && !(~(local_bb0_cmp_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp_i_NO_SHIFT_REG <= 'x;
		local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp_i_NO_SHIFT_REG <= 'x;
			local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp_i_output_regs_ready)
			begin
				local_bb0_cmp_i_NO_SHIFT_REG <= ((rstag_4to4_bb0_and1_i & 32'hFF) == 32'hFF);
				local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= local_bb0_cmp_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp_i_stall_in))
				begin
					local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= local_bb0_cmp_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp_i_inputs_ready)
			begin
				local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_not_cmp10_i_valid_out;
wire local_bb0_not_cmp10_i_stall_in;
wire local_bb0_not_cmp10_i_inputs_ready;
wire local_bb0_not_cmp10_i_stall_local;
wire local_bb0_not_cmp10_i;

assign local_bb0_not_cmp10_i_inputs_ready = local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG;
assign local_bb0_not_cmp10_i = (local_bb0_cmp10_i_NO_SHIFT_REG ^ 1'b1);
assign local_bb0_not_cmp10_i_valid_out = local_bb0_not_cmp10_i_inputs_ready;
assign local_bb0_not_cmp10_i_stall_local = local_bb0_not_cmp10_i_stall_in;
assign local_bb0_cmp10_i_stall_in_1 = (|local_bb0_not_cmp10_i_stall_local);

// This section implements a staging register.
// 
wire rstag_5to5_bb0_cmp_i_valid_out_0;
wire rstag_5to5_bb0_cmp_i_stall_in_0;
wire rstag_5to5_bb0_cmp_i_valid_out_1;
wire rstag_5to5_bb0_cmp_i_stall_in_1;
wire rstag_5to5_bb0_cmp_i_valid_out_2;
wire rstag_5to5_bb0_cmp_i_stall_in_2;
wire rstag_5to5_bb0_cmp_i_valid_out_3;
wire rstag_5to5_bb0_cmp_i_stall_in_3;
wire rstag_5to5_bb0_cmp_i_inputs_ready;
wire rstag_5to5_bb0_cmp_i_stall_local;
 reg rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb0_cmp_i_combined_valid;
 reg rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG;
wire rstag_5to5_bb0_cmp_i;
 reg rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG;

assign rstag_5to5_bb0_cmp_i_inputs_ready = local_bb0_cmp_i_valid_out_NO_SHIFT_REG;
assign rstag_5to5_bb0_cmp_i = (rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG : local_bb0_cmp_i_NO_SHIFT_REG);
assign rstag_5to5_bb0_cmp_i_combined_valid = (rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG | rstag_5to5_bb0_cmp_i_inputs_ready);
assign rstag_5to5_bb0_cmp_i_stall_local = ((rstag_5to5_bb0_cmp_i_stall_in_0 & ~(rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_1 & ~(rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_2 & ~(rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_3 & ~(rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG)));
assign rstag_5to5_bb0_cmp_i_valid_out_0 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_1 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_2 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_3 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG));
assign local_bb0_cmp_i_stall_in = (|rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_5to5_bb0_cmp_i_stall_local)
			begin
				if (~(rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb0_cmp_i_inputs_ready;
				end
			end
			else
			begin
				rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG <= local_bb0_cmp_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_0)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_1)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_2)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_3)) & rstag_5to5_bb0_cmp_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_conv22_i_inputs_ready;
 reg local_bb0_conv22_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_conv22_i_valid_out_NO_SHIFT_REG;
wire local_bb0_conv22_i_stall_in;
wire local_bb0_conv22_i_output_regs_ready;
 reg [31:0] local_bb0_conv22_i_NO_SHIFT_REG;
wire local_bb0_conv22_i_causedstall;

assign local_bb0_conv22_i_inputs_ready = rstag_5to5_bb0_cmp_i_valid_out_0;
assign local_bb0_conv22_i_output_regs_ready = (~(local_bb0_conv22_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_conv22_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_conv22_i_stall_in))));
assign rstag_5to5_bb0_cmp_i_stall_in_0 = (~(local_bb0_conv22_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_conv22_i_output_regs_ready) | ~(local_bb0_conv22_i_inputs_ready)));
assign local_bb0_conv22_i_causedstall = (local_bb0_conv22_i_inputs_ready && (~(local_bb0_conv22_i_output_regs_ready) && !(~(local_bb0_conv22_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_conv22_i_NO_SHIFT_REG <= 'x;
		local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_conv22_i_NO_SHIFT_REG <= 'x;
			local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_conv22_i_output_regs_ready)
			begin
				local_bb0_conv22_i_NO_SHIFT_REG <= rstag_5to5_bb0_cmp_i;
				local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= local_bb0_conv22_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_conv22_i_stall_in))
				begin
					local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= local_bb0_conv22_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_conv22_i_inputs_ready)
			begin
				local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__7_i_inputs_ready;
 reg local_bb0__7_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__7_i_valid_out_NO_SHIFT_REG;
wire local_bb0__7_i_stall_in;
wire local_bb0__7_i_output_regs_ready;
 reg local_bb0__7_i_NO_SHIFT_REG;
wire local_bb0__7_i_causedstall;

assign local_bb0__7_i_inputs_ready = (local_bb0_not_cmp10_i_valid_out & rstag_5to5_bb0_cmp_i_valid_out_1);
assign local_bb0__7_i_output_regs_ready = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__7_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__7_i_stall_in))));
assign local_bb0_not_cmp10_i_stall_in = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__7_i_output_regs_ready) | ~(local_bb0__7_i_inputs_ready)));
assign rstag_5to5_bb0_cmp_i_stall_in_1 = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__7_i_output_regs_ready) | ~(local_bb0__7_i_inputs_ready)));
assign local_bb0__7_i_causedstall = (local_bb0__7_i_inputs_ready && (~(local_bb0__7_i_output_regs_ready) && !(~(local_bb0__7_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__7_i_NO_SHIFT_REG <= 'x;
		local_bb0__7_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__7_i_NO_SHIFT_REG <= 'x;
			local_bb0__7_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__7_i_output_regs_ready)
			begin
				local_bb0__7_i_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i | local_bb0_not_cmp10_i);
				local_bb0__7_i_valid_out_NO_SHIFT_REG <= local_bb0__7_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__7_i_stall_in))
				begin
					local_bb0__7_i_valid_out_NO_SHIFT_REG <= local_bb0__7_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__7_i_inputs_ready)
			begin
				local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_not_cmp_i_valid_out;
wire local_bb0_not_cmp_i_stall_in;
wire local_bb0_not_cmp_i_inputs_ready;
wire local_bb0_not_cmp_i_stall_local;
wire local_bb0_not_cmp_i;

assign local_bb0_not_cmp_i_inputs_ready = rstag_5to5_bb0_cmp_i_valid_out_2;
assign local_bb0_not_cmp_i = (rstag_5to5_bb0_cmp_i ^ 1'b1);
assign local_bb0_not_cmp_i_valid_out = local_bb0_not_cmp_i_inputs_ready;
assign local_bb0_not_cmp_i_stall_local = local_bb0_not_cmp_i_stall_in;
assign rstag_5to5_bb0_cmp_i_stall_in_2 = (|local_bb0_not_cmp_i_stall_local);

// This section implements a registered operation.
// 
wire local_bb0___i_inputs_ready;
 reg local_bb0___i_wii_reg_NO_SHIFT_REG;
 reg local_bb0___i_valid_out_0_NO_SHIFT_REG;
wire local_bb0___i_stall_in_0;
 reg local_bb0___i_valid_out_1_NO_SHIFT_REG;
wire local_bb0___i_stall_in_1;
wire local_bb0___i_output_regs_ready;
 reg local_bb0___i_NO_SHIFT_REG;
wire local_bb0___i_causedstall;

assign local_bb0___i_inputs_ready = (local_bb0_lnot6_i_valid_out_NO_SHIFT_REG & rstag_5to5_bb0_cmp_i_valid_out_3);
assign local_bb0___i_output_regs_ready = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0___i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0___i_stall_in_0)) & (~(local_bb0___i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0___i_stall_in_1))));
assign local_bb0_lnot6_i_stall_in = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & (~(local_bb0___i_output_regs_ready) | ~(local_bb0___i_inputs_ready)));
assign rstag_5to5_bb0_cmp_i_stall_in_3 = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & (~(local_bb0___i_output_regs_ready) | ~(local_bb0___i_inputs_ready)));
assign local_bb0___i_causedstall = (local_bb0___i_inputs_ready && (~(local_bb0___i_output_regs_ready) && !(~(local_bb0___i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0___i_NO_SHIFT_REG <= 'x;
		local_bb0___i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0___i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0___i_NO_SHIFT_REG <= 'x;
			local_bb0___i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0___i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0___i_output_regs_ready)
			begin
				local_bb0___i_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i & local_bb0_lnot6_i_NO_SHIFT_REG);
				local_bb0___i_valid_out_0_NO_SHIFT_REG <= local_bb0___i_inputs_ready;
				local_bb0___i_valid_out_1_NO_SHIFT_REG <= local_bb0___i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0___i_stall_in_0))
				begin
					local_bb0___i_valid_out_0_NO_SHIFT_REG <= local_bb0___i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0___i_stall_in_1))
				begin
					local_bb0___i_valid_out_1_NO_SHIFT_REG <= local_bb0___i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0___i_inputs_ready)
			begin
				local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_6to6_bb0__7_i_valid_out_0;
wire rstag_6to6_bb0__7_i_stall_in_0;
wire rstag_6to6_bb0__7_i_valid_out_1;
wire rstag_6to6_bb0__7_i_stall_in_1;
wire rstag_6to6_bb0__7_i_inputs_ready;
wire rstag_6to6_bb0__7_i_stall_local;
 reg rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG;
wire rstag_6to6_bb0__7_i_combined_valid;
 reg rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG;
wire rstag_6to6_bb0__7_i;
 reg rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG;
 reg rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG;

assign rstag_6to6_bb0__7_i_inputs_ready = local_bb0__7_i_valid_out_NO_SHIFT_REG;
assign rstag_6to6_bb0__7_i = (rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG ? rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG : local_bb0__7_i_NO_SHIFT_REG);
assign rstag_6to6_bb0__7_i_combined_valid = (rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG | rstag_6to6_bb0__7_i_inputs_ready);
assign rstag_6to6_bb0__7_i_stall_local = ((rstag_6to6_bb0__7_i_stall_in_0 & ~(rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG)) | (rstag_6to6_bb0__7_i_stall_in_1 & ~(rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG)));
assign rstag_6to6_bb0__7_i_valid_out_0 = (rstag_6to6_bb0__7_i_combined_valid & ~(rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG));
assign rstag_6to6_bb0__7_i_valid_out_1 = (rstag_6to6_bb0__7_i_combined_valid & ~(rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__7_i_stall_in = (|rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_6to6_bb0__7_i_stall_local)
			begin
				if (~(rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= rstag_6to6_bb0__7_i_inputs_ready;
				end
			end
			else
			begin
				rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG <= local_bb0__7_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= (rstag_6to6_bb0__7_i_combined_valid & (rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG | ~(rstag_6to6_bb0__7_i_stall_in_0)) & rstag_6to6_bb0__7_i_stall_local);
			rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= (rstag_6to6_bb0__7_i_combined_valid & (rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG | ~(rstag_6to6_bb0__7_i_stall_in_1)) & rstag_6to6_bb0__7_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__4_i_inputs_ready;
 reg local_bb0__4_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__4_i_valid_out_NO_SHIFT_REG;
wire local_bb0__4_i_stall_in;
wire local_bb0__4_i_output_regs_ready;
 reg local_bb0__4_i_NO_SHIFT_REG;
wire local_bb0__4_i_causedstall;

assign local_bb0__4_i_inputs_ready = (local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG & local_bb0_not_cmp_i_valid_out);
assign local_bb0__4_i_output_regs_ready = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__4_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__4_i_stall_in))));
assign local_bb0_cmp10_i_stall_in_0 = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__4_i_output_regs_ready) | ~(local_bb0__4_i_inputs_ready)));
assign local_bb0_not_cmp_i_stall_in = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__4_i_output_regs_ready) | ~(local_bb0__4_i_inputs_ready)));
assign local_bb0__4_i_causedstall = (local_bb0__4_i_inputs_ready && (~(local_bb0__4_i_output_regs_ready) && !(~(local_bb0__4_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__4_i_NO_SHIFT_REG <= 'x;
		local_bb0__4_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__4_i_NO_SHIFT_REG <= 'x;
			local_bb0__4_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__4_i_output_regs_ready)
			begin
				local_bb0__4_i_NO_SHIFT_REG <= (local_bb0_cmp10_i_NO_SHIFT_REG & local_bb0_not_cmp_i);
				local_bb0__4_i_valid_out_NO_SHIFT_REG <= local_bb0__4_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__4_i_stall_in))
				begin
					local_bb0__4_i_valid_out_NO_SHIFT_REG <= local_bb0__4_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__4_i_inputs_ready)
			begin
				local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_conv44_i_stall_local;
wire [31:0] local_bb0_conv44_i;

assign local_bb0_conv44_i[31:1] = 31'h0;
assign local_bb0_conv44_i[0] = local_bb0___i_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb0_cond50_i_stall_local;
wire [31:0] local_bb0_cond50_i;

assign local_bb0_cond50_i = (local_bb0___i_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements a registered operation.
// 
wire local_bb0__12_i_inputs_ready;
 reg local_bb0__12_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__12_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0__12_i_stall_in_0;
 reg local_bb0__12_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0__12_i_stall_in_1;
wire local_bb0__12_i_output_regs_ready;
 reg local_bb0__12_i_NO_SHIFT_REG;
wire local_bb0__12_i_causedstall;

assign local_bb0__12_i_inputs_ready = rstag_6to6_bb0__7_i_valid_out_0;
assign local_bb0__12_i_output_regs_ready = (~(local_bb0__12_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0__12_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0__12_i_stall_in_0)) & (~(local_bb0__12_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0__12_i_stall_in_1))));
assign rstag_6to6_bb0__7_i_stall_in_0 = (~(local_bb0__12_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__12_i_output_regs_ready) | ~(local_bb0__12_i_inputs_ready)));
assign local_bb0__12_i_causedstall = (local_bb0__12_i_inputs_ready && (~(local_bb0__12_i_output_regs_ready) && !(~(local_bb0__12_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__12_i_NO_SHIFT_REG <= 'x;
		local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__12_i_NO_SHIFT_REG <= 'x;
			local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__12_i_output_regs_ready)
			begin
				local_bb0__12_i_NO_SHIFT_REG <= (1'b0 & rstag_6to6_bb0__7_i);
				local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= local_bb0__12_i_inputs_ready;
				local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= local_bb0__12_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__12_i_stall_in_0))
				begin
					local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= local_bb0__12_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0__12_i_stall_in_1))
				begin
					local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= local_bb0__12_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__12_i_inputs_ready)
			begin
				local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__8_i_inputs_ready;
 reg local_bb0__8_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__8_i_valid_out_NO_SHIFT_REG;
wire local_bb0__8_i_stall_in;
wire local_bb0__8_i_output_regs_ready;
 reg local_bb0__8_i_NO_SHIFT_REG;
wire local_bb0__8_i_causedstall;

assign local_bb0__8_i_inputs_ready = rstag_6to6_bb0__7_i_valid_out_1;
assign local_bb0__8_i_output_regs_ready = (~(local_bb0__8_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__8_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__8_i_stall_in))));
assign rstag_6to6_bb0__7_i_stall_in_1 = (~(local_bb0__8_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__8_i_output_regs_ready) | ~(local_bb0__8_i_inputs_ready)));
assign local_bb0__8_i_causedstall = (local_bb0__8_i_inputs_ready && (~(local_bb0__8_i_output_regs_ready) && !(~(local_bb0__8_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__8_i_NO_SHIFT_REG <= 'x;
		local_bb0__8_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__8_i_NO_SHIFT_REG <= 'x;
			local_bb0__8_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__8_i_output_regs_ready)
			begin
				local_bb0__8_i_NO_SHIFT_REG <= (1'b1 & rstag_6to6_bb0__7_i);
				local_bb0__8_i_valid_out_NO_SHIFT_REG <= local_bb0__8_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__8_i_stall_in))
				begin
					local_bb0__8_i_valid_out_NO_SHIFT_REG <= local_bb0__8_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__8_i_inputs_ready)
			begin
				local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_7to7_bb0__4_i_valid_out_0;
wire rstag_7to7_bb0__4_i_stall_in_0;
wire rstag_7to7_bb0__4_i_valid_out_1;
wire rstag_7to7_bb0__4_i_stall_in_1;
wire rstag_7to7_bb0__4_i_inputs_ready;
wire rstag_7to7_bb0__4_i_stall_local;
 reg rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG;
wire rstag_7to7_bb0__4_i_combined_valid;
 reg rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG;
wire rstag_7to7_bb0__4_i;
 reg rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG;
 reg rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG;

assign rstag_7to7_bb0__4_i_inputs_ready = local_bb0__4_i_valid_out_NO_SHIFT_REG;
assign rstag_7to7_bb0__4_i = (rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG ? rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG : local_bb0__4_i_NO_SHIFT_REG);
assign rstag_7to7_bb0__4_i_combined_valid = (rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG | rstag_7to7_bb0__4_i_inputs_ready);
assign rstag_7to7_bb0__4_i_stall_local = ((rstag_7to7_bb0__4_i_stall_in_0 & ~(rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG)) | (rstag_7to7_bb0__4_i_stall_in_1 & ~(rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG)));
assign rstag_7to7_bb0__4_i_valid_out_0 = (rstag_7to7_bb0__4_i_combined_valid & ~(rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG));
assign rstag_7to7_bb0__4_i_valid_out_1 = (rstag_7to7_bb0__4_i_combined_valid & ~(rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__4_i_stall_in = (|rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_7to7_bb0__4_i_stall_local)
			begin
				if (~(rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= rstag_7to7_bb0__4_i_inputs_ready;
				end
			end
			else
			begin
				rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG <= local_bb0__4_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= (rstag_7to7_bb0__4_i_combined_valid & (rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG | ~(rstag_7to7_bb0__4_i_stall_in_0)) & rstag_7to7_bb0__4_i_stall_local);
			rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= (rstag_7to7_bb0__4_i_combined_valid & (rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG | ~(rstag_7to7_bb0__4_i_stall_in_1)) & rstag_7to7_bb0__4_i_stall_local);
		end
	end
end


// This section implements a staging register.
// 
wire rstag_7to7_bb0__8_i_valid_out_0;
wire rstag_7to7_bb0__8_i_stall_in_0;
wire rstag_7to7_bb0__8_i_valid_out_1;
wire rstag_7to7_bb0__8_i_stall_in_1;
wire rstag_7to7_bb0__8_i_inputs_ready;
wire rstag_7to7_bb0__8_i_stall_local;
 reg rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG;
wire rstag_7to7_bb0__8_i_combined_valid;
 reg rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG;
wire rstag_7to7_bb0__8_i;
 reg rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG;
 reg rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG;

assign rstag_7to7_bb0__8_i_inputs_ready = local_bb0__8_i_valid_out_NO_SHIFT_REG;
assign rstag_7to7_bb0__8_i = (rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG ? rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG : local_bb0__8_i_NO_SHIFT_REG);
assign rstag_7to7_bb0__8_i_combined_valid = (rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG | rstag_7to7_bb0__8_i_inputs_ready);
assign rstag_7to7_bb0__8_i_stall_local = ((rstag_7to7_bb0__8_i_stall_in_0 & ~(rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG)) | (rstag_7to7_bb0__8_i_stall_in_1 & ~(rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG)));
assign rstag_7to7_bb0__8_i_valid_out_0 = (rstag_7to7_bb0__8_i_combined_valid & ~(rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG));
assign rstag_7to7_bb0__8_i_valid_out_1 = (rstag_7to7_bb0__8_i_combined_valid & ~(rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__8_i_stall_in = (|rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_7to7_bb0__8_i_stall_local)
			begin
				if (~(rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= rstag_7to7_bb0__8_i_inputs_ready;
				end
			end
			else
			begin
				rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG <= local_bb0__8_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i_combined_valid & (rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG | ~(rstag_7to7_bb0__8_i_stall_in_0)) & rstag_7to7_bb0__8_i_stall_local);
			rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i_combined_valid & (rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG | ~(rstag_7to7_bb0__8_i_stall_in_1)) & rstag_7to7_bb0__8_i_stall_local);
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0__17_i_stall_local;
wire [31:0] local_bb0__17_i;

assign local_bb0__17_i = (rstag_7to7_bb0__4_i ? 32'h0 : 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb0__5_i_valid_out;
wire local_bb0__5_i_stall_in;
wire local_bb0__5_i_inputs_ready;
wire local_bb0__5_i_stall_local;
wire [31:0] local_bb0__5_i;

assign local_bb0__5_i_inputs_ready = rstag_7to7_bb0__4_i_valid_out_1;
assign local_bb0__5_i[31:1] = 31'h0;
assign local_bb0__5_i[0] = rstag_7to7_bb0__4_i;
assign local_bb0__5_i_valid_out = local_bb0__5_i_inputs_ready;
assign local_bb0__5_i_stall_local = local_bb0__5_i_stall_in;
assign rstag_7to7_bb0__4_i_stall_in_1 = (|local_bb0__5_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0__18_i_valid_out;
wire local_bb0__18_i_stall_in;
wire local_bb0__18_i_inputs_ready;
wire local_bb0__18_i_stall_local;
wire [31:0] local_bb0__18_i;

assign local_bb0__18_i_inputs_ready = (rstag_7to7_bb0__4_i_valid_out_0 & rstag_7to7_bb0__8_i_valid_out_0);
assign local_bb0__18_i = (rstag_7to7_bb0__8_i ? 32'h1 : (local_bb0__17_i & 32'h100));
assign local_bb0__18_i_valid_out = local_bb0__18_i_inputs_ready;
assign local_bb0__18_i_stall_local = local_bb0__18_i_stall_in;
assign rstag_7to7_bb0__4_i_stall_in_0 = (local_bb0__18_i_stall_local | ~(local_bb0__18_i_inputs_ready));
assign rstag_7to7_bb0__8_i_stall_in_0 = (local_bb0__18_i_stall_local | ~(local_bb0__18_i_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb0__9_i_inputs_ready;
 reg local_bb0__9_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__9_i_valid_out_NO_SHIFT_REG;
wire local_bb0__9_i_stall_in;
wire local_bb0__9_i_output_regs_ready;
 reg [31:0] local_bb0__9_i_NO_SHIFT_REG;
wire local_bb0__9_i_causedstall;

assign local_bb0__9_i_inputs_ready = (local_bb0__5_i_valid_out & rstag_7to7_bb0__8_i_valid_out_1);
assign local_bb0__9_i_output_regs_ready = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__9_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__9_i_stall_in))));
assign local_bb0__5_i_stall_in = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__9_i_output_regs_ready) | ~(local_bb0__9_i_inputs_ready)));
assign rstag_7to7_bb0__8_i_stall_in_1 = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__9_i_output_regs_ready) | ~(local_bb0__9_i_inputs_ready)));
assign local_bb0__9_i_causedstall = (local_bb0__9_i_inputs_ready && (~(local_bb0__9_i_output_regs_ready) && !(~(local_bb0__9_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__9_i_NO_SHIFT_REG <= 'x;
		local_bb0__9_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__9_i_NO_SHIFT_REG <= 'x;
			local_bb0__9_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__9_i_output_regs_ready)
			begin
				local_bb0__9_i_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i ? 32'h0 : (local_bb0__5_i & 32'h1));
				local_bb0__9_i_valid_out_NO_SHIFT_REG <= local_bb0__9_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__9_i_stall_in))
				begin
					local_bb0__9_i_valid_out_NO_SHIFT_REG <= local_bb0__9_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__9_i_inputs_ready)
			begin
				local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__19_i_inputs_ready;
 reg local_bb0__19_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__19_i_valid_out_NO_SHIFT_REG;
wire local_bb0__19_i_stall_in;
wire local_bb0__19_i_output_regs_ready;
 reg [31:0] local_bb0__19_i_NO_SHIFT_REG;
wire local_bb0__19_i_causedstall;

assign local_bb0__19_i_inputs_ready = (local_bb0__12_i_valid_out_1_NO_SHIFT_REG & local_bb0__18_i_valid_out);
assign local_bb0__19_i_output_regs_ready = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__19_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__19_i_stall_in))));
assign local_bb0__12_i_stall_in_1 = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__19_i_output_regs_ready) | ~(local_bb0__19_i_inputs_ready)));
assign local_bb0__18_i_stall_in = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__19_i_output_regs_ready) | ~(local_bb0__19_i_inputs_ready)));
assign local_bb0__19_i_causedstall = (local_bb0__19_i_inputs_ready && (~(local_bb0__19_i_output_regs_ready) && !(~(local_bb0__19_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__19_i_NO_SHIFT_REG <= 'x;
		local_bb0__19_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__19_i_NO_SHIFT_REG <= 'x;
			local_bb0__19_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__19_i_output_regs_ready)
			begin
				local_bb0__19_i_NO_SHIFT_REG <= ((local_bb0__12_i_NO_SHIFT_REG & 1'b0) ? 32'hFFFFFF00 : (local_bb0__18_i & 32'h101));
				local_bb0__19_i_valid_out_NO_SHIFT_REG <= local_bb0__19_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__19_i_stall_in))
				begin
					local_bb0__19_i_valid_out_NO_SHIFT_REG <= local_bb0__19_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__19_i_inputs_ready)
			begin
				local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0__13_i_valid_out;
wire local_bb0__13_i_stall_in;
wire local_bb0__13_i_inputs_ready;
wire local_bb0__13_i_stall_local;
wire [31:0] local_bb0__13_i;

assign local_bb0__13_i_inputs_ready = (local_bb0__12_i_valid_out_0_NO_SHIFT_REG & local_bb0__9_i_valid_out_NO_SHIFT_REG);
assign local_bb0__13_i = ((local_bb0__12_i_NO_SHIFT_REG & 1'b0) ? 32'h0 : (local_bb0__9_i_NO_SHIFT_REG & 32'h1));
assign local_bb0__13_i_valid_out = local_bb0__13_i_inputs_ready;
assign local_bb0__13_i_stall_local = local_bb0__13_i_stall_in;
assign local_bb0__12_i_stall_in_0 = (local_bb0__13_i_stall_local | ~(local_bb0__13_i_inputs_ready));
assign local_bb0__9_i_stall_in = (local_bb0__13_i_stall_local | ~(local_bb0__13_i_inputs_ready));

// This section implements a staging register.
// 
wire rstag_8to8_bb0__19_i_valid_out_0;
wire rstag_8to8_bb0__19_i_stall_in_0;
wire rstag_8to8_bb0__19_i_valid_out_1;
wire rstag_8to8_bb0__19_i_stall_in_1;
wire rstag_8to8_bb0__19_i_inputs_ready;
wire rstag_8to8_bb0__19_i_stall_local;
 reg rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG;
wire rstag_8to8_bb0__19_i_combined_valid;
 reg [31:0] rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_8to8_bb0__19_i;
 reg rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG;
 reg rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG;

assign rstag_8to8_bb0__19_i_inputs_ready = local_bb0__19_i_valid_out_NO_SHIFT_REG;
assign rstag_8to8_bb0__19_i = (rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG ? rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG : (local_bb0__19_i_NO_SHIFT_REG & 32'hFFFFFF01));
assign rstag_8to8_bb0__19_i_combined_valid = (rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG | rstag_8to8_bb0__19_i_inputs_ready);
assign rstag_8to8_bb0__19_i_stall_local = ((rstag_8to8_bb0__19_i_stall_in_0 & ~(rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG)) | (rstag_8to8_bb0__19_i_stall_in_1 & ~(rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG)));
assign rstag_8to8_bb0__19_i_valid_out_0 = (rstag_8to8_bb0__19_i_combined_valid & ~(rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG));
assign rstag_8to8_bb0__19_i_valid_out_1 = (rstag_8to8_bb0__19_i_combined_valid & ~(rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__19_i_stall_in = (|rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_8to8_bb0__19_i_stall_local)
			begin
				if (~(rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= rstag_8to8_bb0__19_i_inputs_ready;
				end
			end
			else
			begin
				rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG <= (local_bb0__19_i_NO_SHIFT_REG & 32'hFFFFFF01);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= (rstag_8to8_bb0__19_i_combined_valid & (rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG | ~(rstag_8to8_bb0__19_i_stall_in_0)) & rstag_8to8_bb0__19_i_stall_local);
			rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= (rstag_8to8_bb0__19_i_combined_valid & (rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG | ~(rstag_8to8_bb0__19_i_stall_in_1)) & rstag_8to8_bb0__19_i_stall_local);
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_fold_i_valid_out;
wire local_bb0_fold_i_stall_in;
wire local_bb0_fold_i_inputs_ready;
wire local_bb0_fold_i_stall_local;
wire [31:0] local_bb0_fold_i;

assign local_bb0_fold_i_inputs_ready = (local_bb0_shr_i_valid_out_1_NO_SHIFT_REG & rstag_8to8_bb0__19_i_valid_out_0);
assign local_bb0_fold_i = ((rstag_8to8_bb0__19_i & 32'hFFFFFF01) + (local_bb0_shr_i_NO_SHIFT_REG & 32'h1FF));
assign local_bb0_fold_i_valid_out = local_bb0_fold_i_inputs_ready;
assign local_bb0_fold_i_stall_local = local_bb0_fold_i_stall_in;
assign local_bb0_shr_i_stall_in_1 = (local_bb0_fold_i_stall_local | ~(local_bb0_fold_i_inputs_ready));
assign rstag_8to8_bb0__19_i_stall_in_0 = (local_bb0_fold_i_stall_local | ~(local_bb0_fold_i_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb0_add_i_inputs_ready;
 reg local_bb0_add_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_add_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_add_i_stall_in_0;
 reg local_bb0_add_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_add_i_stall_in_1;
wire local_bb0_add_i_output_regs_ready;
 reg [31:0] local_bb0_add_i_NO_SHIFT_REG;
wire local_bb0_add_i_causedstall;

assign local_bb0_add_i_inputs_ready = (rstag_8to8_bb0__19_i_valid_out_1 & rstag_4to4_bb0_and1_i_valid_out_0);
assign local_bb0_add_i_output_regs_ready = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_add_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_add_i_stall_in_0)) & (~(local_bb0_add_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_add_i_stall_in_1))));
assign rstag_8to8_bb0__19_i_stall_in_1 = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_add_i_output_regs_ready) | ~(local_bb0_add_i_inputs_ready)));
assign rstag_4to4_bb0_and1_i_stall_in_0 = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_add_i_output_regs_ready) | ~(local_bb0_add_i_inputs_ready)));
assign local_bb0_add_i_causedstall = (local_bb0_add_i_inputs_ready && (~(local_bb0_add_i_output_regs_ready) && !(~(local_bb0_add_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add_i_NO_SHIFT_REG <= 'x;
		local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add_i_NO_SHIFT_REG <= 'x;
			local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add_i_output_regs_ready)
			begin
				local_bb0_add_i_NO_SHIFT_REG <= ((rstag_8to8_bb0__19_i & 32'hFFFFFF01) + (rstag_4to4_bb0_and1_i & 32'hFF));
				local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= local_bb0_add_i_inputs_ready;
				local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= local_bb0_add_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_add_i_stall_in_0))
				begin
					local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= local_bb0_add_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_add_i_stall_in_1))
				begin
					local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= local_bb0_add_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add_i_inputs_ready)
			begin
				local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and32_i_inputs_ready;
 reg local_bb0_and32_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and32_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and32_i_stall_in;
wire local_bb0_and32_i_output_regs_ready;
 reg [31:0] local_bb0_and32_i_NO_SHIFT_REG;
wire local_bb0_and32_i_causedstall;

assign local_bb0_and32_i_inputs_ready = local_bb0_fold_i_valid_out;
assign local_bb0_and32_i_output_regs_ready = (~(local_bb0_and32_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and32_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and32_i_stall_in))));
assign local_bb0_fold_i_stall_in = (~(local_bb0_and32_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and32_i_output_regs_ready) | ~(local_bb0_and32_i_inputs_ready)));
assign local_bb0_and32_i_causedstall = (local_bb0_and32_i_inputs_ready && (~(local_bb0_and32_i_output_regs_ready) && !(~(local_bb0_and32_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and32_i_NO_SHIFT_REG <= 'x;
		local_bb0_and32_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and32_i_NO_SHIFT_REG <= 'x;
			local_bb0_and32_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and32_i_output_regs_ready)
			begin
				local_bb0_and32_i_NO_SHIFT_REG <= (local_bb0_fold_i << 32'h17);
				local_bb0_and32_i_valid_out_NO_SHIFT_REG <= local_bb0_and32_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and32_i_stall_in))
				begin
					local_bb0_and32_i_valid_out_NO_SHIFT_REG <= local_bb0_and32_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and32_i_inputs_ready)
			begin
				local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_cmp20_i_stall_local;
wire local_bb0_cmp20_i;

assign local_bb0_cmp20_i = ($signed(local_bb0_add_i_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb0_cmp25_i_stall_local;
wire local_bb0_cmp25_i;

assign local_bb0_cmp25_i = ($signed(local_bb0_add_i_NO_SHIFT_REG) < $signed(32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_shl_i_stall_local;
wire [31:0] local_bb0_shl_i;

assign local_bb0_shl_i = ((local_bb0_and32_i_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb0_conv_i_valid_out;
wire local_bb0_conv_i_stall_in;
wire local_bb0_conv_i_inputs_ready;
wire local_bb0_conv_i_stall_local;
wire [31:0] local_bb0_conv_i;

assign local_bb0_conv_i_inputs_ready = local_bb0_add_i_valid_out_0_NO_SHIFT_REG;
assign local_bb0_conv_i[31:1] = 31'h0;
assign local_bb0_conv_i[0] = local_bb0_cmp20_i;
assign local_bb0_conv_i_valid_out = local_bb0_conv_i_inputs_ready;
assign local_bb0_conv_i_stall_local = local_bb0_conv_i_stall_in;
assign local_bb0_add_i_stall_in_0 = (|local_bb0_conv_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0_conv26_i_valid_out;
wire local_bb0_conv26_i_stall_in;
wire local_bb0_conv26_i_inputs_ready;
wire local_bb0_conv26_i_stall_local;
wire [31:0] local_bb0_conv26_i;

assign local_bb0_conv26_i_inputs_ready = local_bb0_add_i_valid_out_1_NO_SHIFT_REG;
assign local_bb0_conv26_i[31:1] = 31'h0;
assign local_bb0_conv26_i[0] = local_bb0_cmp25_i;
assign local_bb0_conv26_i_valid_out = local_bb0_conv26_i_inputs_ready;
assign local_bb0_conv26_i_stall_local = local_bb0_conv26_i_stall_in;
assign local_bb0_add_i_stall_in_1 = (|local_bb0_conv26_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0_or34_i_stall_local;
wire [31:0] local_bb0_or34_i;

assign local_bb0_or34_i = ((local_bb0_shl_i & 32'h7F800000) | (local_bb0_and33_i_NO_SHIFT_REG & 32'h807FFFFF));

// This section implements a registered operation.
// 
wire local_bb0_or_i_inputs_ready;
 reg local_bb0_or_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_or_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_or_i_stall_in_0;
 reg local_bb0_or_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_or_i_stall_in_1;
wire local_bb0_or_i_output_regs_ready;
 reg [31:0] local_bb0_or_i_NO_SHIFT_REG;
wire local_bb0_or_i_causedstall;

assign local_bb0_or_i_inputs_ready = (local_bb0_conv_i_valid_out & local_bb0_conv22_i_valid_out_NO_SHIFT_REG);
assign local_bb0_or_i_output_regs_ready = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_or_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_or_i_stall_in_0)) & (~(local_bb0_or_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_or_i_stall_in_1))));
assign local_bb0_conv_i_stall_in = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or_i_output_regs_ready) | ~(local_bb0_or_i_inputs_ready)));
assign local_bb0_conv22_i_stall_in = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or_i_output_regs_ready) | ~(local_bb0_or_i_inputs_ready)));
assign local_bb0_or_i_causedstall = (local_bb0_or_i_inputs_ready && (~(local_bb0_or_i_output_regs_ready) && !(~(local_bb0_or_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or_i_NO_SHIFT_REG <= 'x;
		local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or_i_NO_SHIFT_REG <= 'x;
			local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or_i_output_regs_ready)
			begin
				local_bb0_or_i_NO_SHIFT_REG <= ((local_bb0_conv_i & 32'h1) | (local_bb0_conv22_i_NO_SHIFT_REG & 32'h1));
				local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= local_bb0_or_i_inputs_ready;
				local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= local_bb0_or_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_or_i_stall_in_0))
				begin
					local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= local_bb0_or_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_or_i_stall_in_1))
				begin
					local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= local_bb0_or_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or_i_inputs_ready)
			begin
				local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_or29_i_inputs_ready;
 reg local_bb0_or29_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_or29_i_valid_out_NO_SHIFT_REG;
wire local_bb0_or29_i_stall_in;
wire local_bb0_or29_i_output_regs_ready;
 reg [31:0] local_bb0_or29_i_NO_SHIFT_REG;
wire local_bb0_or29_i_causedstall;

assign local_bb0_or29_i_inputs_ready = (local_bb0_conv26_i_valid_out & local_bb0__13_i_valid_out);
assign local_bb0_or29_i_output_regs_ready = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_or29_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_or29_i_stall_in))));
assign local_bb0_conv26_i_stall_in = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or29_i_output_regs_ready) | ~(local_bb0_or29_i_inputs_ready)));
assign local_bb0__13_i_stall_in = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or29_i_output_regs_ready) | ~(local_bb0_or29_i_inputs_ready)));
assign local_bb0_or29_i_causedstall = (local_bb0_or29_i_inputs_ready && (~(local_bb0_or29_i_output_regs_ready) && !(~(local_bb0_or29_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or29_i_NO_SHIFT_REG <= 'x;
		local_bb0_or29_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or29_i_NO_SHIFT_REG <= 'x;
			local_bb0_or29_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or29_i_output_regs_ready)
			begin
				local_bb0_or29_i_NO_SHIFT_REG <= ((local_bb0_conv26_i & 32'h1) | (local_bb0__13_i & 32'h1));
				local_bb0_or29_i_valid_out_NO_SHIFT_REG <= local_bb0_or29_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_or29_i_stall_in))
				begin
					local_bb0_or29_i_valid_out_NO_SHIFT_REG <= local_bb0_or29_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or29_i_inputs_ready)
			begin
				local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_or45_i_stall_local;
wire [31:0] local_bb0_or45_i;

assign local_bb0_or45_i = ((local_bb0_or_i_NO_SHIFT_REG & 32'h1) | (local_bb0_conv44_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_or39_i_stall_local;
wire [31:0] local_bb0_or39_i;

assign local_bb0_or39_i = ((local_bb0_or29_i_NO_SHIFT_REG & 32'h1) | (local_bb0_or_i_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_tobool46_i_stall_local;
wire local_bb0_tobool46_i;

assign local_bb0_tobool46_i = ((local_bb0_or45_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_tobool40_i_stall_local;
wire local_bb0_tobool40_i;

assign local_bb0_tobool40_i = ((local_bb0_or39_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_cond47_i_stall_local;
wire [31:0] local_bb0_cond47_i;

assign local_bb0_cond47_i = (local_bb0_tobool46_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_cond_i_stall_local;
wire [31:0] local_bb0_cond_i;

assign local_bb0_cond_i = (local_bb0_tobool40_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb0_or52_i_stall_local;
wire [31:0] local_bb0_or52_i;

assign local_bb0_or52_i = ((local_bb0_cond47_i & 32'h7F800000) | (local_bb0_cond50_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb0_and51_i_stall_local;
wire [31:0] local_bb0_and51_i;

assign local_bb0_and51_i = ((local_bb0_cond_i | 32'h80000000) & local_bb0_or34_i);

// This section implements an unregistered operation.
// 
wire local_bb0_or53_i_stall_local;
wire [31:0] local_bb0_or53_i;

assign local_bb0_or53_i = ((local_bb0_or52_i & 32'h7FC00000) | local_bb0_and51_i);

// This section implements an unregistered operation.
// 
wire local_bb0_var__u2_valid_out;
wire local_bb0_var__u2_stall_in;
wire local_bb0_var__u2_inputs_ready;
wire local_bb0_var__u2_stall_local;
wire [31:0] local_bb0_var__u2;

assign local_bb0_var__u2_inputs_ready = (local_bb0_and33_i_valid_out_NO_SHIFT_REG & local_bb0_and32_i_valid_out_NO_SHIFT_REG & local_bb0___i_valid_out_1_NO_SHIFT_REG & local_bb0___i_valid_out_0_NO_SHIFT_REG & local_bb0_or_i_valid_out_1_NO_SHIFT_REG & local_bb0_or29_i_valid_out_NO_SHIFT_REG & local_bb0_or_i_valid_out_0_NO_SHIFT_REG);
assign local_bb0_var__u2 = local_bb0_or53_i;
assign local_bb0_var__u2_valid_out = local_bb0_var__u2_inputs_ready;
assign local_bb0_var__u2_stall_local = local_bb0_var__u2_stall_in;
assign local_bb0_and33_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_and32_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0___i_stall_in_1 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0___i_stall_in_0 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or_i_stall_in_1 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or29_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or_i_stall_in_0 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));

// This section implements a staging register.
// 
wire rstag_10to10_bb0_var__u2_valid_out;
wire rstag_10to10_bb0_var__u2_stall_in;
wire rstag_10to10_bb0_var__u2_inputs_ready;
wire rstag_10to10_bb0_var__u2_stall_local;
 reg rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG;
wire rstag_10to10_bb0_var__u2_combined_valid;
 reg [31:0] rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_10to10_bb0_var__u2;

assign rstag_10to10_bb0_var__u2_inputs_ready = local_bb0_var__u2_valid_out;
assign rstag_10to10_bb0_var__u2 = (rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG ? rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG : local_bb0_var__u2);
assign rstag_10to10_bb0_var__u2_combined_valid = (rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG | rstag_10to10_bb0_var__u2_inputs_ready);
assign rstag_10to10_bb0_var__u2_valid_out = rstag_10to10_bb0_var__u2_combined_valid;
assign rstag_10to10_bb0_var__u2_stall_local = rstag_10to10_bb0_var__u2_stall_in;
assign local_bb0_var__u2_stall_in = (|rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_10to10_bb0_var__u2_stall_local)
			begin
				if (~(rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG))
				begin
					rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= rstag_10to10_bb0_var__u2_inputs_ready;
				end
			end
			else
			begin
				rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG))
		begin
			rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG <= local_bb0_var__u2;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_mul39_inputs_ready;
 reg local_bb0_mul39_wii_reg_NO_SHIFT_REG;
 reg local_bb0_mul39_valid_out_NO_SHIFT_REG;
wire local_bb0_mul39_stall_in;
wire local_bb0_mul39_output_regs_ready;
wire [31:0] local_bb0_mul39;
 reg local_bb0_mul39_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb0_mul39_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb0_mul39_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb0_mul39_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb0_mul39_valid_pipe_4_NO_SHIFT_REG;
wire local_bb0_mul39_causedstall;

acl_fp_mul_ll_s5 fp_module_local_bb0_mul39 (
	.clock(clock),
	.dataa(rstag_10to10_bb0_var__u2),
	.datab(input_e_d),
	.enable(local_bb0_mul39_output_regs_ready),
	.result(local_bb0_mul39)
);


assign local_bb0_mul39_inputs_ready = (merge_node_valid_out_3_NO_SHIFT_REG & rstag_10to10_bb0_var__u2_valid_out);
assign local_bb0_mul39_output_regs_ready = (~(local_bb0_mul39_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_mul39_valid_out_NO_SHIFT_REG) | ~(local_bb0_mul39_stall_in))));
assign merge_node_stall_in_3 = (~(local_bb0_mul39_wii_reg_NO_SHIFT_REG) & (~(local_bb0_mul39_output_regs_ready) | ~(local_bb0_mul39_inputs_ready)));
assign rstag_10to10_bb0_var__u2_stall_in = (~(local_bb0_mul39_wii_reg_NO_SHIFT_REG) & (~(local_bb0_mul39_output_regs_ready) | ~(local_bb0_mul39_inputs_ready)));
assign local_bb0_mul39_causedstall = (local_bb0_mul39_inputs_ready && (~(local_bb0_mul39_output_regs_ready) && !(~(local_bb0_mul39_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul39_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul39_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul39_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul39_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul39_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul39_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul39_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul39_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul39_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul39_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul39_output_regs_ready)
			begin
				local_bb0_mul39_valid_pipe_0_NO_SHIFT_REG <= local_bb0_mul39_inputs_ready;
				local_bb0_mul39_valid_pipe_1_NO_SHIFT_REG <= local_bb0_mul39_valid_pipe_0_NO_SHIFT_REG;
				local_bb0_mul39_valid_pipe_2_NO_SHIFT_REG <= local_bb0_mul39_valid_pipe_1_NO_SHIFT_REG;
				local_bb0_mul39_valid_pipe_3_NO_SHIFT_REG <= local_bb0_mul39_valid_pipe_2_NO_SHIFT_REG;
				local_bb0_mul39_valid_pipe_4_NO_SHIFT_REG <= local_bb0_mul39_valid_pipe_3_NO_SHIFT_REG;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul39_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul39_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul39_output_regs_ready)
			begin
				local_bb0_mul39_valid_out_NO_SHIFT_REG <= local_bb0_mul39_valid_pipe_4_NO_SHIFT_REG;
			end
			else
			begin
				if (~(local_bb0_mul39_stall_in))
				begin
					local_bb0_mul39_valid_out_NO_SHIFT_REG <= local_bb0_mul39_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul39_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul39_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul39_valid_pipe_4_NO_SHIFT_REG)
			begin
				local_bb0_mul39_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg lvb_bb0_cmp1017_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_mul39_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb0_var__reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb0_var__u0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb0_var__u0_valid_out_NO_SHIFT_REG & local_bb0_var__valid_out_NO_SHIFT_REG & local_bb0_mul39_valid_out_NO_SHIFT_REG & local_bb0_cmp1017_valid_out_NO_SHIFT_REG & merge_node_valid_out_5_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb0_var__u0_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_var__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_mul39_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_cmp1017_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign merge_node_stall_in_5 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb0_cmp1017 = lvb_bb0_cmp1017_reg_NO_SHIFT_REG;
assign lvb_bb0_mul39 = lvb_bb0_mul39_reg_NO_SHIFT_REG;
assign lvb_bb0_var_ = lvb_bb0_var__reg_NO_SHIFT_REG;
assign lvb_bb0_var__u0 = lvb_bb0_var__u0_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb0_cmp1017_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_mul39_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__u0_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb0_cmp1017_reg_NO_SHIFT_REG <= local_bb0_cmp1017_NO_SHIFT_REG;
			lvb_bb0_mul39_reg_NO_SHIFT_REG <= local_bb0_mul39;
			lvb_bb0_var__reg_NO_SHIFT_REG <= local_bb0_var__NO_SHIFT_REG;
			lvb_bb0_var__u0_reg_NO_SHIFT_REG <= local_bb0_var__u0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_1
	(
		input 		clock,
		input 		resetn,
		input 		input_wii_cmp1017,
		input [31:0] 		input_wii_mul39,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u3,
		input 		valid_in_0,
		output 		stall_out_0,
		input [63:0] 		input_indvars_iv33_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [63:0] 		input_indvars_iv33_1,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start,
		output [63:0] 		ffwd_0_0,
		output [31:0] 		ffwd_1_0,
		output 		ffwd_2_0,
		output [63:0] 		ffwd_3_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv33_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv33_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv33_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_indvars_iv33_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_indvars_iv33_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_indvars_iv33_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv33_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_indvars_iv33_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv33_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_indvars_iv33_NO_SHIFT_REG <= input_indvars_iv33_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_indvars_iv33_NO_SHIFT_REG <= input_indvars_iv33_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_indvars_iv33_NO_SHIFT_REG <= input_indvars_iv33_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_indvars_iv33_NO_SHIFT_REG <= input_indvars_iv33_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1_var__stall_local;
wire [31:0] local_bb1_var_;

assign local_bb1_var_ = local_lvm_indvars_iv33_NO_SHIFT_REG[31:0];

// This section implements an unregistered operation.
// 
wire local_bb1_var__u4_stall_local;
wire [63:0] local_bb1_var__u4;

assign local_bb1_var__u4 = (local_lvm_indvars_iv33_NO_SHIFT_REG << 64'h6);

// This section implements an unregistered operation.
// 
wire local_bb1_var__u5_stall_local;
wire [63:0] local_bb1_var__u5;

assign local_bb1_var__u5 = (local_lvm_indvars_iv33_NO_SHIFT_REG << 64'h8);

// This section implements an unregistered operation.
// 
wire local_bb1__indvars_iv33_valid_out;
wire local_bb1__indvars_iv33_stall_in;
wire local_bb1__indvars_iv33_inputs_ready;
wire local_bb1__indvars_iv33_stall_local;
 reg [63:0] ffwd_0_0_reg_NO_SHIFT_REG;

assign local_bb1__indvars_iv33_inputs_ready = merge_node_valid_out_3_NO_SHIFT_REG;
assign ffwd_0_0 = ffwd_0_0_reg_NO_SHIFT_REG;
assign local_bb1__indvars_iv33_valid_out = local_bb1__indvars_iv33_inputs_ready;
assign local_bb1__indvars_iv33_stall_local = local_bb1__indvars_iv33_stall_in;
assign merge_node_stall_in_3 = (|local_bb1__indvars_iv33_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb1__indvars_iv33_inputs_ready))
	begin
		ffwd_0_0_reg_NO_SHIFT_REG <= local_lvm_indvars_iv33_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1_cmp_stall_local;
wire local_bb1_cmp;

assign local_bb1_cmp = (local_bb1_var_ < 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb1___stall_local;
 reg [31:0] ffwd_1_0_reg_NO_SHIFT_REG;
wire local_bb1___inputs_ready;

assign ffwd_1_0 = ffwd_1_0_reg_NO_SHIFT_REG;

always @(posedge clock)
begin
	if ((1'b1 & local_bb1___inputs_ready))
	begin
		ffwd_1_0_reg_NO_SHIFT_REG <= local_bb1_var_;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1__add126_stall_local;
wire [63:0] local_bb1__add126;

assign local_bb1__add126 = ((local_bb1_var__u4 & 64'hFFFFFFFFFFFFFFC0) + (local_bb1_var__u5 & 64'hFFFFFFFFFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb1___valid_out;
wire local_bb1___stall_in;
wire local_bb1__cmp_valid_out;
wire local_bb1__cmp_stall_in;
wire local_bb1__cmp_inputs_ready;
wire local_bb1__cmp_stall_local;
 reg ffwd_2_0_reg_NO_SHIFT_REG;
 reg local_bb1___consumed_0_NO_SHIFT_REG;
 reg local_bb1__cmp_consumed_0_NO_SHIFT_REG;

assign local_bb1__cmp_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb1___inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign ffwd_2_0 = ffwd_2_0_reg_NO_SHIFT_REG;
assign local_bb1__cmp_stall_local = ((local_bb1___stall_in & ~(local_bb1___consumed_0_NO_SHIFT_REG)) | (local_bb1__cmp_stall_in & ~(local_bb1__cmp_consumed_0_NO_SHIFT_REG)));
assign local_bb1___valid_out = (local_bb1__cmp_inputs_ready & ~(local_bb1___consumed_0_NO_SHIFT_REG));
assign local_bb1__cmp_valid_out = (local_bb1__cmp_inputs_ready & ~(local_bb1__cmp_consumed_0_NO_SHIFT_REG));
assign merge_node_stall_in_0 = (|local_bb1__cmp_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb1__cmp_inputs_ready))
	begin
		ffwd_2_0_reg_NO_SHIFT_REG <= local_bb1_cmp;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1___consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb1__cmp_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb1___consumed_0_NO_SHIFT_REG <= (local_bb1__cmp_inputs_ready & (local_bb1___consumed_0_NO_SHIFT_REG | ~(local_bb1___stall_in)) & local_bb1__cmp_stall_local);
		local_bb1__cmp_consumed_0_NO_SHIFT_REG <= (local_bb1__cmp_inputs_ready & (local_bb1__cmp_consumed_0_NO_SHIFT_REG | ~(local_bb1__cmp_stall_in)) & local_bb1__cmp_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1___add126_valid_out;
wire local_bb1___add126_stall_in;
wire local_bb1___add126_inputs_ready;
wire local_bb1___add126_stall_local;
 reg [63:0] ffwd_3_0_reg_NO_SHIFT_REG;

assign local_bb1___add126_inputs_ready = (merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG);
assign ffwd_3_0 = ffwd_3_0_reg_NO_SHIFT_REG;
assign local_bb1___add126_valid_out = local_bb1___add126_inputs_ready;
assign local_bb1___add126_stall_local = local_bb1___add126_stall_in;
assign merge_node_stall_in_1 = (local_bb1___add126_stall_local | ~(local_bb1___add126_inputs_ready));
assign merge_node_stall_in_2 = (local_bb1___add126_stall_local | ~(local_bb1___add126_inputs_ready));

always @(posedge clock)
begin
	if ((1'b1 & local_bb1___add126_inputs_ready))
	begin
		ffwd_3_0_reg_NO_SHIFT_REG <= (local_bb1__add126 & 64'hFFFFFFFFFFFFFFC0);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb1___0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb1___0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb1___0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb1___0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1___0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1___0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb1___0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb1___0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb1___0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb1___0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb1___0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to2_bb1___0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb1___0_reg_2_fifo.DATA_WIDTH = 0;
defparam rnode_1to2_bb1___0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb1___0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb1___0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb1___valid_out;
assign local_bb1___stall_in = rnode_1to2_bb1___0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb1___0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb1___0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb1___0_valid_out_NO_SHIFT_REG = rnode_1to2_bb1___0_valid_out_reg_2_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb1__cmp_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb1__cmp_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb1__cmp_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb1__cmp_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1__cmp_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1__cmp_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb1__cmp_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb1__cmp_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb1__cmp_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb1__cmp_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb1__cmp_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to2_bb1__cmp_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb1__cmp_0_reg_2_fifo.DATA_WIDTH = 0;
defparam rnode_1to2_bb1__cmp_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb1__cmp_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb1__cmp_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb1__cmp_valid_out;
assign local_bb1__cmp_stall_in = rnode_1to2_bb1__cmp_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb1__cmp_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb1__cmp_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb1__cmp_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb1__cmp_0_valid_out_reg_2_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_1to2_rc0_bb1___add126_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to2_rc0_bb1___add126_0_stall_in_NO_SHIFT_REG;
 logic rcnode_1to2_rc0_bb1___add126_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rcnode_1to2_rc0_bb1___add126_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rcnode_1to2_rc0_bb1___add126_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rcnode_1to2_rc0_bb1___add126_0_stall_out_0_reg_2_IP_NO_SHIFT_REG;
 logic rcnode_1to2_rc0_bb1___add126_0_stall_out_0_reg_2_NO_SHIFT_REG;

acl_data_fifo rcnode_1to2_rc0_bb1___add126_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to2_rc0_bb1___add126_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to2_rc0_bb1___add126_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rcnode_1to2_rc0_bb1___add126_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rcnode_1to2_rc0_bb1___add126_0_stall_out_0_reg_2_IP_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rcnode_1to2_rc0_bb1___add126_0_reg_2_fifo.DEPTH = 1;
defparam rcnode_1to2_rc0_bb1___add126_0_reg_2_fifo.DATA_WIDTH = 0;
defparam rcnode_1to2_rc0_bb1___add126_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_1to2_rc0_bb1___add126_0_reg_2_fifo.IMPL = "ll_reg";

assign rcnode_1to2_rc0_bb1___add126_0_reg_2_inputs_ready_NO_SHIFT_REG = (local_bb1___add126_valid_out & local_bb1__indvars_iv33_valid_out);
assign rcnode_1to2_rc0_bb1___add126_0_stall_out_0_reg_2_NO_SHIFT_REG = (~(rcnode_1to2_rc0_bb1___add126_0_reg_2_inputs_ready_NO_SHIFT_REG) | rcnode_1to2_rc0_bb1___add126_0_stall_out_0_reg_2_IP_NO_SHIFT_REG);
assign local_bb1___add126_stall_in = rcnode_1to2_rc0_bb1___add126_0_stall_out_0_reg_2_NO_SHIFT_REG;
assign local_bb1__indvars_iv33_stall_in = rcnode_1to2_rc0_bb1___add126_0_stall_out_0_reg_2_NO_SHIFT_REG;
assign rcnode_1to2_rc0_bb1___add126_0_stall_in_reg_2_NO_SHIFT_REG = rcnode_1to2_rc0_bb1___add126_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to2_rc0_bb1___add126_0_valid_out_NO_SHIFT_REG = rcnode_1to2_rc0_bb1___add126_0_valid_out_reg_2_NO_SHIFT_REG;

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;

assign branch_var__inputs_ready = (rnode_1to2_bb1__cmp_0_valid_out_NO_SHIFT_REG & rnode_1to2_bb1___0_valid_out_NO_SHIFT_REG & rcnode_1to2_rc0_bb1___add126_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign rnode_1to2_bb1__cmp_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to2_bb1___0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_1to2_rc0_bb1___add126_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_2
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_in,
		input 		input_wii_cmp1017,
		input [31:0] 		input_wii_mul39,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u6,
		input 		valid_in_0,
		output 		stall_out_0,
		input [63:0] 		input_indvars_iv30_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [63:0] 		input_indvars_iv30_1,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start,
		input [63:0] 		ffwd_3_0,
		output [63:0] 		ffwd_4_0,
		output [31:0] 		ffwd_5_0,
		input 		ffwd_2_0,
		output [63:0] 		ffwd_7_0,
		output 		ffwd_6_0,
		input [511:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [32:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [511:0] 		avm_local_bb2_ld__writedata,
		output [63:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		output 		local_bb2_ld__active,
		input 		clock2x,
		output [31:0] 		ffwd_8_0,
		output 		ffwd_9_0,
		output 		ffwd_10_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv30_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv30_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv30_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_indvars_iv30_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_indvars_iv30_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_indvars_iv30_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv30_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_indvars_iv30_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv30_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_indvars_iv30_NO_SHIFT_REG <= input_indvars_iv30_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_indvars_iv30_NO_SHIFT_REG <= input_indvars_iv30_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_indvars_iv30_NO_SHIFT_REG <= input_indvars_iv30_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_indvars_iv30_NO_SHIFT_REG <= input_indvars_iv30_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__stall_local;
wire [31:0] local_bb2_var_;

assign local_bb2_var_ = local_lvm_indvars_iv30_NO_SHIFT_REG[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2__add126192_acl_ffwd_dest_i64_3_stall_local;
wire [63:0] local_bb2__add126192_acl_ffwd_dest_i64_3;

assign local_bb2__add126192_acl_ffwd_dest_i64_3 = ffwd_3_0;

// This section implements an unregistered operation.
// 
wire local_bb2__indvars_iv30_valid_out;
wire local_bb2__indvars_iv30_stall_in;
wire local_bb2__indvars_iv30_inputs_ready;
wire local_bb2__indvars_iv30_stall_local;
 reg [63:0] ffwd_4_0_reg_NO_SHIFT_REG;

assign local_bb2__indvars_iv30_inputs_ready = merge_node_valid_out_3_NO_SHIFT_REG;
assign ffwd_4_0 = ffwd_4_0_reg_NO_SHIFT_REG;
assign local_bb2__indvars_iv30_valid_out = local_bb2__indvars_iv30_inputs_ready;
assign local_bb2__indvars_iv30_stall_local = local_bb2__indvars_iv30_stall_in;
assign merge_node_stall_in_3 = (|local_bb2__indvars_iv30_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2__indvars_iv30_inputs_ready))
	begin
		ffwd_4_0_reg_NO_SHIFT_REG <= local_lvm_indvars_iv30_NO_SHIFT_REG;
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_fifo.DEPTH = 3;
defparam rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_reg_3_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_4_NO_SHIFT_REG;
assign merge_node_stall_in_4 = rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_in_reg_3_NO_SHIFT_REG = rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_in_NO_SHIFT_REG;
assign rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_valid_out_NO_SHIFT_REG = rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_valid_out_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp2_stall_local;
wire local_bb2_cmp2;

assign local_bb2_cmp2 = (local_bb2_var_ < 32'h140);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp2_valid_out;
wire local_bb2_cmp2_stall_in;
wire local_bb2___valid_out;
wire local_bb2___stall_in;
wire local_bb2___inputs_ready;
wire local_bb2___stall_local;
 reg [31:0] ffwd_5_0_reg_NO_SHIFT_REG;
 reg local_bb2_cmp2_consumed_0_NO_SHIFT_REG;
 reg local_bb2___consumed_0_NO_SHIFT_REG;

assign local_bb2___inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign ffwd_5_0 = ffwd_5_0_reg_NO_SHIFT_REG;
assign local_bb2___stall_local = ((local_bb2_cmp2_stall_in & ~(local_bb2_cmp2_consumed_0_NO_SHIFT_REG)) | (local_bb2___stall_in & ~(local_bb2___consumed_0_NO_SHIFT_REG)));
assign local_bb2_cmp2_valid_out = (local_bb2___inputs_ready & ~(local_bb2_cmp2_consumed_0_NO_SHIFT_REG));
assign local_bb2___valid_out = (local_bb2___inputs_ready & ~(local_bb2___consumed_0_NO_SHIFT_REG));
assign merge_node_stall_in_0 = (|local_bb2___stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___inputs_ready))
	begin
		ffwd_5_0_reg_NO_SHIFT_REG <= local_bb2_var_;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp2_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2___consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp2_consumed_0_NO_SHIFT_REG <= (local_bb2___inputs_ready & (local_bb2_cmp2_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp2_stall_in)) & local_bb2___stall_local);
		local_bb2___consumed_0_NO_SHIFT_REG <= (local_bb2___inputs_ready & (local_bb2___consumed_0_NO_SHIFT_REG | ~(local_bb2___stall_in)) & local_bb2___stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__u7_valid_out;
wire local_bb2_var__u7_stall_in;
wire local_bb2_var__u7_inputs_ready;
wire local_bb2_var__u7_stall_local;
wire [63:0] local_bb2_var__u7;

assign local_bb2_var__u7_inputs_ready = (merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG);
assign local_bb2_var__u7 = (local_lvm_indvars_iv30_NO_SHIFT_REG + local_bb2__add126192_acl_ffwd_dest_i64_3);
assign local_bb2_var__u7_valid_out = local_bb2_var__u7_inputs_ready;
assign local_bb2_var__u7_stall_local = local_bb2_var__u7_stall_in;
assign merge_node_stall_in_1 = (local_bb2_var__u7_stall_local | ~(local_bb2_var__u7_inputs_ready));
assign merge_node_stall_in_2 = (local_bb2_var__u7_stall_local | ~(local_bb2_var__u7_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb2_cmp191_acl_ffwd_dest_i1_2_stall_local;
wire local_bb2_cmp191_acl_ffwd_dest_i1_2;

assign local_bb2_cmp191_acl_ffwd_dest_i1_2 = ffwd_2_0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb2_cmp2_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp2_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp2_0_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp2_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp2_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp2_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp2_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp2_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb2_cmp2_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb2_cmp2_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb2_cmp2_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb2_cmp2_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb2_cmp2_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb2_cmp2),
	.data_out(rnode_1to3_bb2_cmp2_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb2_cmp2_0_reg_3_fifo.DEPTH = 3;
defparam rnode_1to3_bb2_cmp2_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb2_cmp2_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to3_bb2_cmp2_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_1to3_bb2_cmp2_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb2_cmp2_valid_out;
assign local_bb2_cmp2_stall_in = rnode_1to3_bb2_cmp2_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb2_cmp2_0_NO_SHIFT_REG = rnode_1to3_bb2_cmp2_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb2_cmp2_0_stall_in_reg_3_NO_SHIFT_REG = rnode_1to3_bb2_cmp2_0_stall_in_NO_SHIFT_REG;
assign rnode_1to3_bb2_cmp2_0_valid_out_NO_SHIFT_REG = rnode_1to3_bb2_cmp2_0_valid_out_reg_3_NO_SHIFT_REG;

// Register node:
//  * latency = 164
//  * capacity = 164
 logic rcnode_1to165_rc0_bb2__indvars_iv30_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_in_NO_SHIFT_REG;
 logic rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rcnode_1to165_rc0_bb2__indvars_iv30_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_out_0_reg_165_IP_NO_SHIFT_REG;
 logic rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_out_0_reg_165_NO_SHIFT_REG;

acl_data_fifo rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rcnode_1to165_rc0_bb2__indvars_iv30_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_out_0_reg_165_IP_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_fifo.DEPTH = 165;
defparam rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_fifo.DATA_WIDTH = 0;
defparam rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_fifo.IMPL = "ram";

assign rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_inputs_ready_NO_SHIFT_REG = (local_bb2__indvars_iv30_valid_out & local_bb2___valid_out);
assign rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_out_0_reg_165_NO_SHIFT_REG = (~(rcnode_1to165_rc0_bb2__indvars_iv30_0_reg_165_inputs_ready_NO_SHIFT_REG) | rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_out_0_reg_165_IP_NO_SHIFT_REG);
assign local_bb2__indvars_iv30_stall_in = rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_out_0_reg_165_NO_SHIFT_REG;
assign local_bb2___stall_in = rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_out_0_reg_165_NO_SHIFT_REG;
assign rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_in_reg_165_NO_SHIFT_REG = rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to165_rc0_bb2__indvars_iv30_0_valid_out_NO_SHIFT_REG = rcnode_1to165_rc0_bb2__indvars_iv30_0_valid_out_reg_165_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb2_var__u7_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u7_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb2_var__u7_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u7_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u7_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb2_var__u7_1_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u7_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb2_var__u7_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u7_0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u7_0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u7_0_stall_out_reg_2_NO_SHIFT_REG;
 reg rnode_1to2_bb2_var__u7_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to2_bb2_var__u7_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb2_var__u7_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb2_var__u7_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb2_var__u7_0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb2_var__u7_0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb2_var__u7_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb2_var__u7),
	.data_out(rnode_1to2_bb2_var__u7_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb2_var__u7_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb2_var__u7_0_reg_2_fifo.DATA_WIDTH = 64;
defparam rnode_1to2_bb2_var__u7_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb2_var__u7_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb2_var__u7_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb2_var__u7_valid_out;
assign local_bb2_var__u7_stall_in = rnode_1to2_bb2_var__u7_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u7_0_stall_in_0_reg_2_NO_SHIFT_REG = ((rnode_1to2_bb2_var__u7_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__u7_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to2_bb2_var__u7_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__u7_0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to2_bb2_var__u7_0_valid_out_0_NO_SHIFT_REG = (rnode_1to2_bb2_var__u7_0_valid_out_0_reg_2_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__u7_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to2_bb2_var__u7_0_valid_out_1_NO_SHIFT_REG = (rnode_1to2_bb2_var__u7_0_valid_out_0_reg_2_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__u7_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to2_bb2_var__u7_0_NO_SHIFT_REG = rnode_1to2_bb2_var__u7_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u7_1_NO_SHIFT_REG = rnode_1to2_bb2_var__u7_0_reg_2_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to2_bb2_var__u7_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to2_bb2_var__u7_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to2_bb2_var__u7_0_consumed_0_NO_SHIFT_REG <= (rnode_1to2_bb2_var__u7_0_valid_out_0_reg_2_NO_SHIFT_REG & (rnode_1to2_bb2_var__u7_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to2_bb2_var__u7_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to2_bb2_var__u7_0_stall_in_0_reg_2_NO_SHIFT_REG);
		rnode_1to2_bb2_var__u7_0_consumed_1_NO_SHIFT_REG <= (rnode_1to2_bb2_var__u7_0_valid_out_0_reg_2_NO_SHIFT_REG & (rnode_1to2_bb2_var__u7_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to2_bb2_var__u7_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to2_bb2_var__u7_0_stall_in_0_reg_2_NO_SHIFT_REG);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__u8_stall_local;
wire local_bb2_var__u8;

assign local_bb2_var__u8 = (local_bb2_cmp191_acl_ffwd_dest_i1_2 & rnode_1to3_bb2_cmp2_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx_valid_out;
wire local_bb2_arrayidx_stall_in;
wire local_bb2_arrayidx_inputs_ready;
wire local_bb2_arrayidx_stall_local;
wire [63:0] local_bb2_arrayidx;

assign local_bb2_arrayidx_inputs_ready = rnode_1to2_bb2_var__u7_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_arrayidx = ((input_in & 64'hFFFFFFFFFFFFFC00) + (rnode_1to2_bb2_var__u7_0_NO_SHIFT_REG << 6'h2));
assign local_bb2_arrayidx_valid_out = local_bb2_arrayidx_inputs_ready;
assign local_bb2_arrayidx_stall_local = local_bb2_arrayidx_stall_in;
assign rnode_1to2_bb2_var__u7_0_stall_in_0_NO_SHIFT_REG = (|local_bb2_arrayidx_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb2___u9_valid_out;
wire local_bb2___u9_stall_in;
wire local_bb2___u9_inputs_ready;
wire local_bb2___u9_stall_local;
 reg [63:0] ffwd_7_0_reg_NO_SHIFT_REG;

assign local_bb2___u9_inputs_ready = rnode_1to2_bb2_var__u7_0_valid_out_1_NO_SHIFT_REG;
assign ffwd_7_0 = ffwd_7_0_reg_NO_SHIFT_REG;
assign local_bb2___u9_valid_out = local_bb2___u9_inputs_ready;
assign local_bb2___u9_stall_local = local_bb2___u9_stall_in;
assign rnode_1to2_bb2_var__u7_0_stall_in_1_NO_SHIFT_REG = (|local_bb2___u9_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___u9_inputs_ready))
	begin
		ffwd_7_0_reg_NO_SHIFT_REG <= rnode_1to2_bb2_var__u7_1_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2__phi_decision_xor_stall_local;
wire local_bb2__phi_decision_xor;

assign local_bb2__phi_decision_xor = (local_bb2_var__u8 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__phi_decision_xor_valid_out;
wire local_bb2__phi_decision_xor_stall_in;
wire local_bb2___u10_valid_out;
wire local_bb2___u10_stall_in;
wire local_bb2___u10_inputs_ready;
wire local_bb2___u10_stall_local;
 reg ffwd_6_0_reg_NO_SHIFT_REG;
 reg local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG;
 reg local_bb2___u10_consumed_0_NO_SHIFT_REG;

assign local_bb2___u10_inputs_ready = (rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_valid_out_NO_SHIFT_REG & rnode_1to3_bb2_cmp2_0_valid_out_NO_SHIFT_REG);
assign ffwd_6_0 = ffwd_6_0_reg_NO_SHIFT_REG;
assign local_bb2___u10_stall_local = ((local_bb2__phi_decision_xor_stall_in & ~(local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG)) | (local_bb2___u10_stall_in & ~(local_bb2___u10_consumed_0_NO_SHIFT_REG)));
assign local_bb2__phi_decision_xor_valid_out = (local_bb2___u10_inputs_ready & ~(local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG));
assign local_bb2___u10_valid_out = (local_bb2___u10_inputs_ready & ~(local_bb2___u10_consumed_0_NO_SHIFT_REG));
assign rnode_1to3_bb2_cmp191_acl_ffwd_dest_i1_2_0_stall_in_NO_SHIFT_REG = (local_bb2___u10_stall_local | ~(local_bb2___u10_inputs_ready));
assign rnode_1to3_bb2_cmp2_0_stall_in_NO_SHIFT_REG = (local_bb2___u10_stall_local | ~(local_bb2___u10_inputs_ready));

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___u10_inputs_ready))
	begin
		ffwd_6_0_reg_NO_SHIFT_REG <= local_bb2_var__u8;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2___u10_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= (local_bb2___u10_inputs_ready & (local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG | ~(local_bb2__phi_decision_xor_stall_in)) & local_bb2___u10_stall_local);
		local_bb2___u10_consumed_0_NO_SHIFT_REG <= (local_bb2___u10_inputs_ready & (local_bb2___u10_consumed_0_NO_SHIFT_REG | ~(local_bb2___u10_stall_in)) & local_bb2___u10_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb2_arrayidx_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb2_arrayidx_0_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb2_arrayidx_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb2_arrayidx_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb2_arrayidx_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb2_arrayidx_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb2_arrayidx_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb2_arrayidx_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in((local_bb2_arrayidx & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_2to3_bb2_arrayidx_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.DEPTH = 2;
defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.DATA_WIDTH = 64;
defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_2to3_bb2_arrayidx_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb2_arrayidx_valid_out;
assign local_bb2_arrayidx_stall_in = rnode_2to3_bb2_arrayidx_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx_0_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx_0_stall_in_reg_3_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx_0_stall_in_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx_0_valid_out_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx_0_valid_out_reg_3_NO_SHIFT_REG;

// Register node:
//  * latency = 163
//  * capacity = 163
 logic rnode_2to165_bb2___u9_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to165_bb2___u9_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to165_bb2___u9_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to165_bb2___u9_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_2to165_bb2___u9_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_2to165_bb2___u9_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_2to165_bb2___u9_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to165_bb2___u9_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to165_bb2___u9_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_2to165_bb2___u9_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_2to165_bb2___u9_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to165_bb2___u9_0_reg_165_fifo.DEPTH = 164;
defparam rnode_2to165_bb2___u9_0_reg_165_fifo.DATA_WIDTH = 0;
defparam rnode_2to165_bb2___u9_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_2to165_bb2___u9_0_reg_165_fifo.IMPL = "ram";

assign rnode_2to165_bb2___u9_0_reg_165_inputs_ready_NO_SHIFT_REG = local_bb2___u9_valid_out;
assign local_bb2___u9_stall_in = rnode_2to165_bb2___u9_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_2to165_bb2___u9_0_stall_in_reg_165_NO_SHIFT_REG = rnode_2to165_bb2___u9_0_stall_in_NO_SHIFT_REG;
assign rnode_2to165_bb2___u9_0_valid_out_NO_SHIFT_REG = rnode_2to165_bb2___u9_0_valid_out_reg_165_NO_SHIFT_REG;

// This section implements a staging register.
// 
wire rstag_3to3_bb2__phi_decision_xor_valid_out_0;
wire rstag_3to3_bb2__phi_decision_xor_stall_in_0;
wire rstag_3to3_bb2__phi_decision_xor_valid_out_1;
wire rstag_3to3_bb2__phi_decision_xor_stall_in_1;
wire rstag_3to3_bb2__phi_decision_xor_inputs_ready;
wire rstag_3to3_bb2__phi_decision_xor_stall_local;
 reg rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG;
wire rstag_3to3_bb2__phi_decision_xor_combined_valid;
 reg rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG;
wire rstag_3to3_bb2__phi_decision_xor;
 reg rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG;
 reg rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG;

assign rstag_3to3_bb2__phi_decision_xor_inputs_ready = local_bb2__phi_decision_xor_valid_out;
assign rstag_3to3_bb2__phi_decision_xor = (rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG ? rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG : local_bb2__phi_decision_xor);
assign rstag_3to3_bb2__phi_decision_xor_combined_valid = (rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG | rstag_3to3_bb2__phi_decision_xor_inputs_ready);
assign rstag_3to3_bb2__phi_decision_xor_stall_local = ((rstag_3to3_bb2__phi_decision_xor_stall_in_0 & ~(rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG)) | (rstag_3to3_bb2__phi_decision_xor_stall_in_1 & ~(rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG)));
assign rstag_3to3_bb2__phi_decision_xor_valid_out_0 = (rstag_3to3_bb2__phi_decision_xor_combined_valid & ~(rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG));
assign rstag_3to3_bb2__phi_decision_xor_valid_out_1 = (rstag_3to3_bb2__phi_decision_xor_combined_valid & ~(rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG));
assign local_bb2__phi_decision_xor_stall_in = (|rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_3to3_bb2__phi_decision_xor_stall_local)
		begin
			if (~(rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG))
			begin
				rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG <= rstag_3to3_bb2__phi_decision_xor_inputs_ready;
			end
		end
		else
		begin
			rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG))
		begin
			rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG <= local_bb2__phi_decision_xor;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= (rstag_3to3_bb2__phi_decision_xor_combined_valid & (rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG | ~(rstag_3to3_bb2__phi_decision_xor_stall_in_0)) & rstag_3to3_bb2__phi_decision_xor_stall_local);
		rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG <= (rstag_3to3_bb2__phi_decision_xor_combined_valid & (rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG | ~(rstag_3to3_bb2__phi_decision_xor_stall_in_1)) & rstag_3to3_bb2__phi_decision_xor_stall_local);
	end
end


// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_3to165_bb2___u10_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u10_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u10_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u10_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u10_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u10_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_3to165_bb2___u10_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to165_bb2___u10_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to165_bb2___u10_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_3to165_bb2___u10_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_3to165_bb2___u10_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to165_bb2___u10_0_reg_165_fifo.DEPTH = 163;
defparam rnode_3to165_bb2___u10_0_reg_165_fifo.DATA_WIDTH = 0;
defparam rnode_3to165_bb2___u10_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_3to165_bb2___u10_0_reg_165_fifo.IMPL = "ram";

assign rnode_3to165_bb2___u10_0_reg_165_inputs_ready_NO_SHIFT_REG = local_bb2___u10_valid_out;
assign local_bb2___u10_stall_in = rnode_3to165_bb2___u10_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_3to165_bb2___u10_0_stall_in_reg_165_NO_SHIFT_REG = rnode_3to165_bb2___u10_0_stall_in_NO_SHIFT_REG;
assign rnode_3to165_bb2___u10_0_valid_out_NO_SHIFT_REG = rnode_3to165_bb2___u10_0_valid_out_reg_165_NO_SHIFT_REG;

// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_3to165_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to165_bb2__phi_decision_xor_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to165_bb2__phi_decision_xor_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_3to165_bb2__phi_decision_xor_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_3to165_bb2__phi_decision_xor_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(rstag_3to3_bb2__phi_decision_xor),
	.data_out(rnode_3to165_bb2__phi_decision_xor_0_reg_165_NO_SHIFT_REG)
);

defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.DEPTH = 163;
defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.DATA_WIDTH = 1;
defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.IMPL = "ram";

assign rnode_3to165_bb2__phi_decision_xor_0_reg_165_inputs_ready_NO_SHIFT_REG = rstag_3to3_bb2__phi_decision_xor_valid_out_0;
assign rstag_3to3_bb2__phi_decision_xor_stall_in_0 = rnode_3to165_bb2__phi_decision_xor_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_reg_165_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_stall_in_reg_165_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_valid_out_reg_165_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb2_ld__inputs_ready;
 reg local_bb2_ld__valid_out_NO_SHIFT_REG;
wire local_bb2_ld__stall_in;
wire local_bb2_ld__output_regs_ready;
wire local_bb2_ld__fu_stall_out;
wire local_bb2_ld__fu_valid_out;
wire [31:0] local_bb2_ld__lsu_dataout;
 reg [31:0] local_bb2_ld__NO_SHIFT_REG;
wire local_bb2_ld__causedstall;

lsu_top lsu_local_bb2_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld__fu_stall_out),
	.i_valid(local_bb2_ld__inputs_ready),
	.i_address((rnode_2to3_bb2_arrayidx_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_3to3_bb2__phi_decision_xor),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld__output_regs_ready)),
	.o_valid(local_bb2_ld__fu_valid_out),
	.o_readdata(local_bb2_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld__active),
	.avm_address(avm_local_bb2_ld__address),
	.avm_read(avm_local_bb2_ld__read),
	.avm_readdata(avm_local_bb2_ld__readdata),
	.avm_write(avm_local_bb2_ld__write),
	.avm_writeack(avm_local_bb2_ld__writeack),
	.avm_burstcount(avm_local_bb2_ld__burstcount),
	.avm_writedata(avm_local_bb2_ld__writedata),
	.avm_byteenable(avm_local_bb2_ld__byteenable),
	.avm_waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld_.AWIDTH = 33;
defparam lsu_local_bb2_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb2_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb2_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb2_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld_.READ = 1;
defparam lsu_local_bb2_ld_.ATOMIC = 0;
defparam lsu_local_bb2_ld_.WIDTH = 32;
defparam lsu_local_bb2_ld_.MWIDTH = 512;
defparam lsu_local_bb2_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld_.MEMORY_SIDE_MEM_LATENCY = 148;
defparam lsu_local_bb2_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb2_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld_.USECACHING = 0;
defparam lsu_local_bb2_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld_.ADDRSPACE = 1;
defparam lsu_local_bb2_ld_.STYLE = "BURST-COALESCED";

assign local_bb2_ld__inputs_ready = (rnode_2to3_bb2_arrayidx_0_valid_out_NO_SHIFT_REG & rstag_3to3_bb2__phi_decision_xor_valid_out_1);
assign local_bb2_ld__output_regs_ready = (&(~(local_bb2_ld__valid_out_NO_SHIFT_REG) | ~(local_bb2_ld__stall_in)));
assign rnode_2to3_bb2_arrayidx_0_stall_in_NO_SHIFT_REG = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign rstag_3to3_bb2__phi_decision_xor_stall_in_1 = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign local_bb2_ld__causedstall = (local_bb2_ld__inputs_ready && (local_bb2_ld__fu_stall_out && !(~(local_bb2_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld__NO_SHIFT_REG <= 'x;
		local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld__output_regs_ready)
		begin
			local_bb2_ld__NO_SHIFT_REG <= local_bb2_ld__lsu_dataout;
			local_bb2_ld__valid_out_NO_SHIFT_REG <= local_bb2_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld__stall_in))
			begin
				local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_165to166_rc0_bb2__indvars_iv30_0_valid_out_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_in_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv30_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_165to166_rc0_bb2__indvars_iv30_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_fifo.DEPTH = 1;
defparam rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_fifo.DATA_WIDTH = 0;
defparam rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_fifo.IMPL = "ll_reg";

assign rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_inputs_ready_NO_SHIFT_REG = (rnode_2to165_bb2___u9_0_valid_out_NO_SHIFT_REG & rnode_3to165_bb2___u10_0_valid_out_NO_SHIFT_REG & rcnode_1to165_rc0_bb2__indvars_iv30_0_valid_out_NO_SHIFT_REG);
assign rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_165to166_rc0_bb2__indvars_iv30_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign rnode_2to165_bb2___u9_0_stall_in_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rnode_3to165_bb2___u10_0_stall_in_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_1to165_rc0_bb2__indvars_iv30_0_stall_in_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_in_NO_SHIFT_REG;
assign rcnode_165to166_rc0_bb2__indvars_iv30_0_valid_out_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv30_0_valid_out_reg_166_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_reg_166_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_165to166_bb2__phi_decision_xor_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_165to166_bb2__phi_decision_xor_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_165to166_bb2__phi_decision_xor_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_165to166_bb2__phi_decision_xor_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(rnode_3to165_bb2__phi_decision_xor_0_NO_SHIFT_REG),
	.data_out(rnode_165to166_bb2__phi_decision_xor_0_reg_166_NO_SHIFT_REG)
);

defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.DEPTH = 1;
defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.DATA_WIDTH = 1;
defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.IMPL = "ll_reg";

assign rnode_165to166_bb2__phi_decision_xor_0_reg_166_inputs_ready_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_165to166_bb2__phi_decision_xor_0_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_reg_166_NO_SHIFT_REG;
assign rnode_165to166_bb2__phi_decision_xor_0_stall_in_reg_166_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
assign rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements a staging register.
// 
wire rstag_163to163_bb2_ld__valid_out_0;
wire rstag_163to163_bb2_ld__stall_in_0;
wire rstag_163to163_bb2_ld__valid_out_1;
wire rstag_163to163_bb2_ld__stall_in_1;
wire rstag_163to163_bb2_ld__inputs_ready;
wire rstag_163to163_bb2_ld__stall_local;
 reg rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG;
wire rstag_163to163_bb2_ld__combined_valid;
 reg [31:0] rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_163to163_bb2_ld_;
 reg rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG;
 reg rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG;

assign rstag_163to163_bb2_ld__inputs_ready = local_bb2_ld__valid_out_NO_SHIFT_REG;
assign rstag_163to163_bb2_ld_ = (rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG ? rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG : local_bb2_ld__NO_SHIFT_REG);
assign rstag_163to163_bb2_ld__combined_valid = (rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG | rstag_163to163_bb2_ld__inputs_ready);
assign rstag_163to163_bb2_ld__stall_local = ((rstag_163to163_bb2_ld__stall_in_0 & ~(rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG)) | (rstag_163to163_bb2_ld__stall_in_1 & ~(rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG)));
assign rstag_163to163_bb2_ld__valid_out_0 = (rstag_163to163_bb2_ld__combined_valid & ~(rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG));
assign rstag_163to163_bb2_ld__valid_out_1 = (rstag_163to163_bb2_ld__combined_valid & ~(rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG));
assign local_bb2_ld__stall_in = (|rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_163to163_bb2_ld__stall_local)
		begin
			if (~(rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG <= rstag_163to163_bb2_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG <= local_bb2_ld__NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG <= (rstag_163to163_bb2_ld__combined_valid & (rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG | ~(rstag_163to163_bb2_ld__stall_in_0)) & rstag_163to163_bb2_ld__stall_local);
		rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG <= (rstag_163to163_bb2_ld__combined_valid & (rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG | ~(rstag_163to163_bb2_ld__stall_in_1)) & rstag_163to163_bb2_ld__stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2___u11_valid_out;
wire local_bb2___u11_stall_in;
wire local_bb2___u11_inputs_ready;
wire local_bb2___u11_stall_local;
 reg [31:0] ffwd_8_0_reg_NO_SHIFT_REG;

assign local_bb2___u11_inputs_ready = rstag_163to163_bb2_ld__valid_out_0;
assign ffwd_8_0 = ffwd_8_0_reg_NO_SHIFT_REG;
assign local_bb2___u11_valid_out = local_bb2___u11_inputs_ready;
assign local_bb2___u11_stall_local = local_bb2___u11_stall_in;
assign rstag_163to163_bb2_ld__stall_in_0 = (|local_bb2___u11_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___u11_inputs_ready))
	begin
		ffwd_8_0_reg_NO_SHIFT_REG <= rstag_163to163_bb2_ld_;
	end
end


// This section implements a registered operation.
// 
wire local_bb2_cmp4_inputs_ready;
 reg local_bb2_cmp4_valid_out_NO_SHIFT_REG;
wire local_bb2_cmp4_stall_in;
wire local_bb2_cmp4_output_regs_ready;
wire local_bb2_cmp4;
 reg local_bb2_cmp4_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_cmp4_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_cmp4_causedstall;

acl_fp_cmp fp_module_local_bb2_cmp4 (
	.clock(clock),
	.dataa(rstag_163to163_bb2_ld_),
	.datab(32'h0),
	.enable(local_bb2_cmp4_output_regs_ready),
	.result(local_bb2_cmp4)
);

defparam fp_module_local_bb2_cmp4.COMPARISON_MODE = 0;

assign local_bb2_cmp4_inputs_ready = rstag_163to163_bb2_ld__valid_out_1;
assign local_bb2_cmp4_output_regs_ready = (&(~(local_bb2_cmp4_valid_out_NO_SHIFT_REG) | ~(local_bb2_cmp4_stall_in)));
assign rstag_163to163_bb2_ld__stall_in_1 = (~(local_bb2_cmp4_output_regs_ready) | ~(local_bb2_cmp4_inputs_ready));
assign local_bb2_cmp4_causedstall = (local_bb2_cmp4_inputs_ready && (~(local_bb2_cmp4_output_regs_ready) && !(~(local_bb2_cmp4_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp4_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp4_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_cmp4_output_regs_ready)
		begin
			local_bb2_cmp4_valid_pipe_0_NO_SHIFT_REG <= local_bb2_cmp4_inputs_ready;
			local_bb2_cmp4_valid_pipe_1_NO_SHIFT_REG <= local_bb2_cmp4_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp4_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_cmp4_output_regs_ready)
		begin
			local_bb2_cmp4_valid_out_NO_SHIFT_REG <= local_bb2_cmp4_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb2_cmp4_stall_in))
			begin
				local_bb2_cmp4_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_163to166_bb2___u11_0_valid_out_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u11_0_stall_in_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u11_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u11_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u11_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u11_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_163to166_bb2___u11_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_163to166_bb2___u11_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_163to166_bb2___u11_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_163to166_bb2___u11_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_163to166_bb2___u11_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_163to166_bb2___u11_0_reg_166_fifo.DEPTH = 4;
defparam rnode_163to166_bb2___u11_0_reg_166_fifo.DATA_WIDTH = 0;
defparam rnode_163to166_bb2___u11_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_163to166_bb2___u11_0_reg_166_fifo.IMPL = "ll_reg";

assign rnode_163to166_bb2___u11_0_reg_166_inputs_ready_NO_SHIFT_REG = local_bb2___u11_valid_out;
assign local_bb2___u11_stall_in = rnode_163to166_bb2___u11_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_163to166_bb2___u11_0_stall_in_reg_166_NO_SHIFT_REG = rnode_163to166_bb2___u11_0_stall_in_NO_SHIFT_REG;
assign rnode_163to166_bb2___u11_0_valid_out_NO_SHIFT_REG = rnode_163to166_bb2___u11_0_valid_out_reg_166_NO_SHIFT_REG;

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_166to166_bb2_cmp4_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_1_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_reg_166_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_valid_out_0_reg_166_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_stall_in_0_reg_166_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp4_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_166to166_bb2_cmp4_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to166_bb2_cmp4_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to166_bb2_cmp4_0_stall_in_0_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_166to166_bb2_cmp4_0_valid_out_0_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_166to166_bb2_cmp4_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(local_bb2_cmp4),
	.data_out(rnode_166to166_bb2_cmp4_0_reg_166_NO_SHIFT_REG)
);

defparam rnode_166to166_bb2_cmp4_0_reg_166_fifo.DEPTH = 3;
defparam rnode_166to166_bb2_cmp4_0_reg_166_fifo.DATA_WIDTH = 1;
defparam rnode_166to166_bb2_cmp4_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_166to166_bb2_cmp4_0_reg_166_fifo.IMPL = "zl_reg";

assign rnode_166to166_bb2_cmp4_0_reg_166_inputs_ready_NO_SHIFT_REG = local_bb2_cmp4_valid_out_NO_SHIFT_REG;
assign local_bb2_cmp4_stall_in = rnode_166to166_bb2_cmp4_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp4_0_stall_in_0_reg_166_NO_SHIFT_REG = (rnode_166to166_bb2_cmp4_0_stall_in_0_NO_SHIFT_REG | rnode_166to166_bb2_cmp4_0_stall_in_1_NO_SHIFT_REG);
assign rnode_166to166_bb2_cmp4_0_valid_out_0_NO_SHIFT_REG = rnode_166to166_bb2_cmp4_0_valid_out_0_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp4_0_valid_out_1_NO_SHIFT_REG = rnode_166to166_bb2_cmp4_0_valid_out_0_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp4_0_NO_SHIFT_REG = rnode_166to166_bb2_cmp4_0_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp4_1_NO_SHIFT_REG = rnode_166to166_bb2_cmp4_0_reg_166_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__cmp4_stall_local;
 reg ffwd_9_0_reg_NO_SHIFT_REG;
wire local_bb2__cmp4_inputs_ready;

assign ffwd_9_0 = ffwd_9_0_reg_NO_SHIFT_REG;

always @(posedge clock)
begin
	if ((1'b1 & local_bb2__cmp4_inputs_ready))
	begin
		ffwd_9_0_reg_NO_SHIFT_REG <= rnode_166to166_bb2_cmp4_0_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__u12_stall_local;
wire local_bb2_var__u12;

assign local_bb2_var__u12 = (rnode_166to166_bb2_cmp4_1_NO_SHIFT_REG | rnode_165to166_bb2__phi_decision_xor_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u13_stall_local;
wire local_bb2_var__u13;

assign local_bb2_var__u13 = (local_bb2_var__u12 | input_wii_cmp1017);

// This section implements an unregistered operation.
// 
wire local_bb2___u14_valid_out;
wire local_bb2___u14_stall_in;
wire local_bb2__cmp4_valid_out;
wire local_bb2__cmp4_stall_in;
wire local_bb2___u14_inputs_ready;
wire local_bb2___u14_stall_local;
 reg ffwd_10_0_reg_NO_SHIFT_REG;

assign local_bb2___u14_inputs_ready = (rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG & rnode_166to166_bb2_cmp4_0_valid_out_1_NO_SHIFT_REG & rnode_166to166_bb2_cmp4_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__cmp4_inputs_ready = (rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG & rnode_166to166_bb2_cmp4_0_valid_out_1_NO_SHIFT_REG & rnode_166to166_bb2_cmp4_0_valid_out_0_NO_SHIFT_REG);
assign ffwd_10_0 = ffwd_10_0_reg_NO_SHIFT_REG;
assign local_bb2___u14_stall_local = (local_bb2___u14_stall_in | local_bb2__cmp4_stall_in);
assign local_bb2___u14_valid_out = local_bb2___u14_inputs_ready;
assign local_bb2__cmp4_valid_out = local_bb2___u14_inputs_ready;
assign rnode_165to166_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG = (local_bb2___u14_stall_local | ~(local_bb2___u14_inputs_ready));
assign rnode_166to166_bb2_cmp4_0_stall_in_1_NO_SHIFT_REG = (local_bb2___u14_stall_local | ~(local_bb2___u14_inputs_ready));
assign rnode_166to166_bb2_cmp4_0_stall_in_0_NO_SHIFT_REG = (local_bb2___u14_stall_local | ~(local_bb2___u14_inputs_ready));

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___u14_inputs_ready))
	begin
		ffwd_10_0_reg_NO_SHIFT_REG <= local_bb2_var__u13;
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;

assign branch_var__inputs_ready = (local_bb2___u14_valid_out & local_bb2__cmp4_valid_out & rnode_163to166_bb2___u11_0_valid_out_NO_SHIFT_REG & rcnode_165to166_rc0_bb2__indvars_iv30_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb2___u14_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb2__cmp4_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_163to166_bb2___u11_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_165to166_rc0_bb2__indvars_iv30_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_3
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_gaussian,
		input [31:0] 		input_r,
		input 		input_wii_cmp1017,
		input [31:0] 		input_wii_mul39,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u15,
		input 		valid_in_0,
		output 		stall_out_0,
		input 		input_forked_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input 		input_forked_1,
		output 		valid_out,
		input 		stall_in,
		output [31:0] 		lvb_bb3_c0_exe1,
		output [63:0] 		lvb_bb3_c0_exe2,
		output 		lvb_bb3_c0_exe3,
		output 		lvb_bb3_c0_exe4,
		output [31:0] 		lvb_bb3_t_219_pop5_,
		output [31:0] 		lvb_bb3_sum_218_pop6_,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		feedback_valid_in_5,
		output 		feedback_stall_out_5,
		input [31:0] 		feedback_data_in_5,
		input 		feedback_valid_in_6,
		output 		feedback_stall_out_6,
		input [31:0] 		feedback_data_in_6,
		input 		feedback_valid_in_4,
		output 		feedback_stall_out_4,
		input [63:0] 		feedback_data_in_4,
		input 		ffwd_10_0,
		output 		feedback_stall_out_2,
		input 		feedback_valid_in_3,
		output 		feedback_stall_out_3,
		input 		feedback_data_in_3,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		input [31:0] 		ffwd_5_0,
		output 		feedback_valid_out_3,
		input 		feedback_stall_in_3,
		output 		feedback_data_out_3,
		output 		feedback_valid_out_4,
		input 		feedback_stall_in_4,
		output [63:0] 		feedback_data_out_4
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg input_forked_0_staging_reg_NO_SHIFT_REG;
 reg local_lvm_forked_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg input_forked_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_forked_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_forked_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_forked_0_staging_reg_NO_SHIFT_REG <= input_forked_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_forked_1_staging_reg_NO_SHIFT_REG <= input_forked_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni1_stall_local;
wire [15:0] local_bb3_c0_eni1;

assign local_bb3_c0_eni1[7:0] = 8'bx;
assign local_bb3_c0_eni1[8] = local_lvm_forked_NO_SHIFT_REG;
assign local_bb3_c0_eni1[15:9] = 7'bx;

// Register node:
//  * latency = 8
//  * capacity = 8
 logic rnode_1to9_forked_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to9_forked_1_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_reg_9_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_out_reg_9_NO_SHIFT_REG;
 reg rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_1to9_forked_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to9_forked_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_1to9_forked_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(local_lvm_forked_NO_SHIFT_REG),
	.data_out(rnode_1to9_forked_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_1to9_forked_0_reg_9_fifo.DEPTH = 9;
defparam rnode_1to9_forked_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_1to9_forked_0_reg_9_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to9_forked_0_reg_9_fifo.IMPL = "ram_plus_reg";

assign rnode_1to9_forked_0_reg_9_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign merge_node_stall_in_1 = rnode_1to9_forked_0_stall_out_reg_9_NO_SHIFT_REG;
assign rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG = ((rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to9_forked_0_valid_out_0_NO_SHIFT_REG = (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to9_forked_0_valid_out_1_NO_SHIFT_REG = (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to9_forked_0_NO_SHIFT_REG = rnode_1to9_forked_0_reg_9_NO_SHIFT_REG;
assign rnode_1to9_forked_1_NO_SHIFT_REG = rnode_1to9_forked_0_reg_9_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG <= (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & (rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG);
		rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG <= (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & (rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_valid_out_1;
wire local_bb3_c0_ene1_stall_in_1;
wire SFC_1_VALID_1_1_0_valid_out_0;
wire SFC_1_VALID_1_1_0_stall_in_0;
wire local_bb3_indvars_iv26_pop4__valid_out;
wire local_bb3_indvars_iv26_pop4__stall_in;
wire local_bb3_c0_enter_c0_eni1_inputs_ready;
wire local_bb3_c0_enter_c0_eni1_stall_local;
wire local_bb3_c0_enter_c0_eni1_input_accepted;
wire [15:0] local_bb3_c0_enter_c0_eni1;
wire local_bb3_c0_exit_c0_exi4_entry_stall;
wire local_bb3_c0_enter_c0_eni1_valid_bit;
wire local_bb3_c0_exit_c0_exi4_output_regs_ready;
wire local_bb3_c0_exit_c0_exi4_valid_in;
wire local_bb3_c0_exit_c0_exi4_phases;
wire local_bb3_c0_enter_c0_eni1_inc_pipelined_thread;
wire local_bb3_c0_enter_c0_eni1_dec_pipelined_thread;
wire local_bb3_c0_enter_c0_eni1_fu_stall_out;

assign local_bb3_c0_enter_c0_eni1_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb3_c0_enter_c0_eni1 = local_bb3_c0_eni1;
assign local_bb3_c0_enter_c0_eni1_input_accepted = (local_bb3_c0_enter_c0_eni1_inputs_ready && !(local_bb3_c0_exit_c0_exi4_entry_stall));
assign local_bb3_c0_enter_c0_eni1_valid_bit = local_bb3_c0_enter_c0_eni1_input_accepted;
assign local_bb3_c0_enter_c0_eni1_inc_pipelined_thread = 1'b1;
assign local_bb3_c0_enter_c0_eni1_dec_pipelined_thread = ~(1'b0);
assign local_bb3_c0_enter_c0_eni1_fu_stall_out = (~(local_bb3_c0_enter_c0_eni1_inputs_ready) | local_bb3_c0_exit_c0_exi4_entry_stall);
assign local_bb3_c0_enter_c0_eni1_stall_local = (local_bb3_c0_ene1_stall_in_1 | SFC_1_VALID_1_1_0_stall_in_0 | local_bb3_indvars_iv26_pop4__stall_in);
assign local_bb3_c0_ene1_valid_out_1 = local_bb3_c0_enter_c0_eni1_inputs_ready;
assign SFC_1_VALID_1_1_0_valid_out_0 = local_bb3_c0_enter_c0_eni1_inputs_ready;
assign local_bb3_indvars_iv26_pop4__valid_out = local_bb3_c0_enter_c0_eni1_inputs_ready;
assign merge_node_stall_in_0 = (|local_bb3_c0_enter_c0_eni1_fu_stall_out);

// This section implements a registered operation.
// 
wire local_bb3_t_219_pop5__inputs_ready;
 reg local_bb3_t_219_pop5__valid_out_NO_SHIFT_REG;
wire local_bb3_t_219_pop5__stall_in;
wire local_bb3_t_219_pop5__output_regs_ready;
wire [31:0] local_bb3_t_219_pop5__result;
wire local_bb3_t_219_pop5__fu_valid_out;
wire local_bb3_t_219_pop5__fu_stall_out;
 reg [31:0] local_bb3_t_219_pop5__NO_SHIFT_REG;
wire local_bb3_t_219_pop5__causedstall;

acl_pop local_bb3_t_219_pop5__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to9_forked_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(32'h0),
	.stall_out(local_bb3_t_219_pop5__fu_stall_out),
	.valid_in(local_bb3_t_219_pop5__inputs_ready),
	.valid_out(local_bb3_t_219_pop5__fu_valid_out),
	.stall_in(~(local_bb3_t_219_pop5__output_regs_ready)),
	.data_out(local_bb3_t_219_pop5__result),
	.feedback_in(feedback_data_in_5),
	.feedback_valid_in(feedback_valid_in_5),
	.feedback_stall_out(feedback_stall_out_5)
);

defparam local_bb3_t_219_pop5__feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_t_219_pop5__feedback.DATA_WIDTH = 32;
defparam local_bb3_t_219_pop5__feedback.STYLE = "REGULAR";

assign local_bb3_t_219_pop5__inputs_ready = rnode_1to9_forked_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_t_219_pop5__output_regs_ready = (&(~(local_bb3_t_219_pop5__valid_out_NO_SHIFT_REG) | ~(local_bb3_t_219_pop5__stall_in)));
assign rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG = (local_bb3_t_219_pop5__fu_stall_out | ~(local_bb3_t_219_pop5__inputs_ready));
assign local_bb3_t_219_pop5__causedstall = (local_bb3_t_219_pop5__inputs_ready && (local_bb3_t_219_pop5__fu_stall_out && !(~(local_bb3_t_219_pop5__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_t_219_pop5__NO_SHIFT_REG <= 'x;
		local_bb3_t_219_pop5__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_t_219_pop5__output_regs_ready)
		begin
			local_bb3_t_219_pop5__NO_SHIFT_REG <= local_bb3_t_219_pop5__result;
			local_bb3_t_219_pop5__valid_out_NO_SHIFT_REG <= local_bb3_t_219_pop5__fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_t_219_pop5__stall_in))
			begin
				local_bb3_t_219_pop5__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_sum_218_pop6__inputs_ready;
 reg local_bb3_sum_218_pop6__valid_out_NO_SHIFT_REG;
wire local_bb3_sum_218_pop6__stall_in;
wire local_bb3_sum_218_pop6__output_regs_ready;
wire [31:0] local_bb3_sum_218_pop6__result;
wire local_bb3_sum_218_pop6__fu_valid_out;
wire local_bb3_sum_218_pop6__fu_stall_out;
 reg [31:0] local_bb3_sum_218_pop6__NO_SHIFT_REG;
wire local_bb3_sum_218_pop6__causedstall;

acl_pop local_bb3_sum_218_pop6__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to9_forked_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(32'h0),
	.stall_out(local_bb3_sum_218_pop6__fu_stall_out),
	.valid_in(local_bb3_sum_218_pop6__inputs_ready),
	.valid_out(local_bb3_sum_218_pop6__fu_valid_out),
	.stall_in(~(local_bb3_sum_218_pop6__output_regs_ready)),
	.data_out(local_bb3_sum_218_pop6__result),
	.feedback_in(feedback_data_in_6),
	.feedback_valid_in(feedback_valid_in_6),
	.feedback_stall_out(feedback_stall_out_6)
);

defparam local_bb3_sum_218_pop6__feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_sum_218_pop6__feedback.DATA_WIDTH = 32;
defparam local_bb3_sum_218_pop6__feedback.STYLE = "REGULAR";

assign local_bb3_sum_218_pop6__inputs_ready = rnode_1to9_forked_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_sum_218_pop6__output_regs_ready = (&(~(local_bb3_sum_218_pop6__valid_out_NO_SHIFT_REG) | ~(local_bb3_sum_218_pop6__stall_in)));
assign rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG = (local_bb3_sum_218_pop6__fu_stall_out | ~(local_bb3_sum_218_pop6__inputs_ready));
assign local_bb3_sum_218_pop6__causedstall = (local_bb3_sum_218_pop6__inputs_ready && (local_bb3_sum_218_pop6__fu_stall_out && !(~(local_bb3_sum_218_pop6__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_sum_218_pop6__NO_SHIFT_REG <= 'x;
		local_bb3_sum_218_pop6__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_sum_218_pop6__output_regs_ready)
		begin
			local_bb3_sum_218_pop6__NO_SHIFT_REG <= local_bb3_sum_218_pop6__result;
			local_bb3_sum_218_pop6__valid_out_NO_SHIFT_REG <= local_bb3_sum_218_pop6__fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_sum_218_pop6__stall_in))
			begin
				local_bb3_sum_218_pop6__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_stall_local;
wire local_bb3_c0_ene1;

assign local_bb3_c0_ene1 = local_bb3_c0_enter_c0_eni1[8];

// This section implements an unregistered operation.
// 
wire SFC_1_VALID_1_1_0_stall_local;
wire SFC_1_VALID_1_1_0;

assign SFC_1_VALID_1_1_0 = local_bb3_c0_enter_c0_eni1_valid_bit;

// This section implements an unregistered operation.
// 
wire local_bb3_indvars_iv26_pop4__stall_local;
wire [63:0] local_bb3_indvars_iv26_pop4_;
wire local_bb3_indvars_iv26_pop4__fu_valid_out;
wire local_bb3_indvars_iv26_pop4__fu_stall_out;

acl_pop local_bb3_indvars_iv26_pop4__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_c0_ene1),
	.predicate(1'b0),
	.data_in(input_wii_var_),
	.stall_out(local_bb3_indvars_iv26_pop4__fu_stall_out),
	.valid_in(SFC_1_VALID_1_1_0),
	.valid_out(local_bb3_indvars_iv26_pop4__fu_valid_out),
	.stall_in(local_bb3_indvars_iv26_pop4__stall_local),
	.data_out(local_bb3_indvars_iv26_pop4_),
	.feedback_in(feedback_data_in_4),
	.feedback_valid_in(feedback_valid_in_4),
	.feedback_stall_out(feedback_stall_out_4)
);

defparam local_bb3_indvars_iv26_pop4__feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_indvars_iv26_pop4__feedback.DATA_WIDTH = 64;
defparam local_bb3_indvars_iv26_pop4__feedback.STYLE = "REGULAR";

assign local_bb3_indvars_iv26_pop4__stall_local = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_c0_ene1_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_c0_ene1_0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_c0_ene1_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene1),
	.data_out(rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene1_stall_in_1 = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_1_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_2_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_1_VALID_1_2_0_inputs_ready;
 reg SFC_1_VALID_1_2_0_valid_out_0_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_0;
 reg SFC_1_VALID_1_2_0_valid_out_1_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_1;
 reg SFC_1_VALID_1_2_0_valid_out_2_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_2;
 reg SFC_1_VALID_1_2_0_valid_out_3_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_3;
wire SFC_1_VALID_1_2_0_output_regs_ready;
 reg SFC_1_VALID_1_2_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_1_2_0_causedstall;

assign SFC_1_VALID_1_2_0_inputs_ready = 1'b1;
assign SFC_1_VALID_1_2_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_1_1_0_stall_in_0 = 1'b0;
assign SFC_1_VALID_1_2_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_1_2_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_1_2_0_output_regs_ready)
		begin
			SFC_1_VALID_1_2_0_NO_SHIFT_REG <= SFC_1_VALID_1_1_0;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb3_indvars_iv26_pop4__0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb3_indvars_iv26_pop4__1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv26_pop4__0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_indvars_iv26_pop4__0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_indvars_iv26_pop4__0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_indvars_iv26_pop4__0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_indvars_iv26_pop4_),
	.data_out(rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_fifo.DATA_WIDTH = 64;
defparam rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_indvars_iv26_pop4__stall_in = 1'b0;
assign rnode_1to2_bb3_indvars_iv26_pop4__0_stall_in_0_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_indvars_iv26_pop4__0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_indvars_iv26_pop4__0_NO_SHIFT_REG = rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_indvars_iv26_pop4__0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_indvars_iv26_pop4__1_NO_SHIFT_REG = rnode_1to2_bb3_indvars_iv26_pop4__0_reg_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__acl_ffwd_dest_i1_10_stall_local;
wire local_bb3__acl_ffwd_dest_i1_10;

assign local_bb3__acl_ffwd_dest_i1_10 = ffwd_10_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_c0_ene1_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_c0_ene1_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_c0_ene1_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_c0_ene1_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb3_c0_ene1_2_NO_SHIFT_REG),
	.data_out(rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_2_3_0_inputs_ready;
 reg SFC_1_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in;
wire SFC_1_VALID_2_3_0_output_regs_ready;
 reg SFC_1_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_2_3_0_causedstall;

assign SFC_1_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_1_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_1_2_0_stall_in_0 = 1'b0;
assign SFC_1_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_2_3_0_output_regs_ready)
		begin
			SFC_1_VALID_2_3_0_NO_SHIFT_REG <= SFC_1_VALID_1_2_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_keep_going200_acl_pipeline_1_inputs_ready;
 reg local_bb3_keep_going200_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb3_keep_going200_acl_pipeline_1_stall_in;
wire local_bb3_keep_going200_acl_pipeline_1_output_regs_ready;
wire local_bb3_keep_going200_acl_pipeline_1_keep_going;
wire local_bb3_keep_going200_acl_pipeline_1_fu_valid_out;
wire local_bb3_keep_going200_acl_pipeline_1_fu_stall_out;
 reg local_bb3_keep_going200_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb3_keep_going200_acl_pipeline_1_feedback_pipelined;
wire local_bb3_keep_going200_acl_pipeline_1_causedstall;

acl_pipeline local_bb3_keep_going200_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb3_keep_going200_acl_pipeline_1_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_keep_going200_acl_pipeline_1_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_keep_going200_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_2),
	.not_exitcond_in(feedback_data_in_3),
	.not_exitcond_valid_in(feedback_valid_in_3),
	.not_exitcond_stall_out(feedback_stall_out_3),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb3_keep_going200_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb3_keep_going200_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb3_keep_going200_acl_pipeline_1_inputs_ready = 1'b1;
assign local_bb3_keep_going200_acl_pipeline_1_output_regs_ready = 1'b1;
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign SFC_1_VALID_1_2_0_stall_in_1 = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb3_keep_going200_acl_pipeline_1_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_keep_going200_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb3_keep_going200_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_keep_going200_acl_pipeline_1_output_regs_ready)
		begin
			local_bb3_keep_going200_acl_pipeline_1_NO_SHIFT_REG <= local_bb3_keep_going200_acl_pipeline_1_keep_going;
			local_bb3_keep_going200_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_keep_going200_acl_pipeline_1_stall_in))
			begin
				local_bb3_keep_going200_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_indvars_iv_next27_stall_local;
wire [63:0] local_bb3_indvars_iv_next27;

assign local_bb3_indvars_iv_next27 = (rnode_1to2_bb3_indvars_iv26_pop4__0_NO_SHIFT_REG + 64'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb3_indvars_iv26_pop4__0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb3_indvars_iv26_pop4__1_NO_SHIFT_REG;
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_stall_in_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_indvars_iv26_pop4__0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_indvars_iv26_pop4__0_stall_in_0_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_0_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_indvars_iv26_pop4__0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb3_indvars_iv26_pop4__1_NO_SHIFT_REG),
	.data_out(rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_fifo.DATA_WIDTH = 64;
defparam rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_indvars_iv26_pop4__0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_indvars_iv26_pop4__0_stall_in_0_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_indvars_iv26_pop4__0_NO_SHIFT_REG = rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_indvars_iv26_pop4__1_NO_SHIFT_REG = rnode_2to3_bb3_indvars_iv26_pop4__0_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__acl_ffwd_dest_i32_5_stall_local;
wire [31:0] local_bb3__acl_ffwd_dest_i32_5;

assign local_bb3__acl_ffwd_dest_i32_5 = ffwd_5_0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_3_4_0_inputs_ready;
 reg SFC_1_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_3_4_0_stall_in;
wire SFC_1_VALID_3_4_0_output_regs_ready;
 reg SFC_1_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_3_4_0_causedstall;

assign SFC_1_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_1_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in = 1'b0;
assign SFC_1_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_3_4_0_output_regs_ready)
		begin
			SFC_1_VALID_3_4_0_NO_SHIFT_REG <= SFC_1_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_keep_going200_acl_pipeline_1_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_keep_going200_acl_pipeline_1_stall_in = 1'b0;
assign rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_NO_SHIFT_REG = rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__stall_local;
wire [31:0] local_bb3_var_;

assign local_bb3_var_ = local_bb3_indvars_iv_next27[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_var__u16_stall_local;
wire [31:0] local_bb3_var__u16;

assign local_bb3_var__u16 = rnode_2to3_bb3_indvars_iv26_pop4__0_NO_SHIFT_REG[31:0];

// This section implements an unregistered operation.
// 
wire local_bb3_var__u17_valid_out;
wire local_bb3_var__u17_stall_in;
wire local_bb3_var__u17_inputs_ready;
wire local_bb3_var__u17_stall_local;
wire [63:0] local_bb3_var__u17;

assign local_bb3_var__u17_inputs_ready = rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_var__u17 = (rnode_2to3_bb3_indvars_iv26_pop4__1_NO_SHIFT_REG + input_wii_var__u15);
assign local_bb3_var__u17_valid_out = 1'b1;
assign rnode_2to3_bb3_indvars_iv26_pop4__0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_4_5_0_inputs_ready;
 reg SFC_1_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_4_5_0_stall_in;
wire SFC_1_VALID_4_5_0_output_regs_ready;
 reg SFC_1_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_4_5_0_causedstall;

assign SFC_1_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_1_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_3_4_0_stall_in = 1'b0;
assign SFC_1_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_4_5_0_output_regs_ready)
		begin
			SFC_1_VALID_4_5_0_NO_SHIFT_REG <= SFC_1_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_cmp10_stall_local;
wire local_bb3_cmp10;

assign local_bb3_cmp10 = ($signed(local_bb3_var_) > $signed(input_r));

// This section implements an unregistered operation.
// 
wire local_bb3_add16_valid_out;
wire local_bb3_add16_stall_in;
wire local_bb3_add16_inputs_ready;
wire local_bb3_add16_stall_local;
wire [31:0] local_bb3_add16;

assign local_bb3_add16_inputs_ready = (rnode_2to3_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_indvars_iv26_pop4__0_valid_out_0_NO_SHIFT_REG);
assign local_bb3_add16 = (local_bb3_var__u16 + local_bb3__acl_ffwd_dest_i32_5);
assign local_bb3_add16_valid_out = 1'b1;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_indvars_iv26_pop4__0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_var__u17_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u17_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_3to4_bb3_var__u17_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u17_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_3to4_bb3_var__u17_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u17_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u17_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u17_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_var__u17_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_var__u17_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_var__u17_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_var__u17_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_var__u17_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_var__u17),
	.data_out(rnode_3to4_bb3_var__u17_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_var__u17_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_var__u17_0_reg_4_fifo.DATA_WIDTH = 64;
defparam rnode_3to4_bb3_var__u17_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_var__u17_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_var__u17_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u17_stall_in = 1'b0;
assign rnode_3to4_bb3_var__u17_0_NO_SHIFT_REG = rnode_3to4_bb3_var__u17_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_var__u17_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_var__u17_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u18_stall_local;
wire local_bb3_var__u18;

assign local_bb3_var__u18 = (local_bb3__acl_ffwd_dest_i1_10 | local_bb3_cmp10);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_add16_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add16_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_add16_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add16_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add16_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_add16_1_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add16_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_add16_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add16_0_valid_out_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add16_0_stall_in_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add16_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_add16_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_add16_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_add16_0_stall_in_0_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_add16_0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_add16_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_add16),
	.data_out(rnode_3to4_bb3_add16_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_add16_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_add16_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3_add16_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_add16_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_add16_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add16_stall_in = 1'b0;
assign rnode_3to4_bb3_add16_0_stall_in_0_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_add16_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_add16_0_NO_SHIFT_REG = rnode_3to4_bb3_add16_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_add16_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_add16_1_NO_SHIFT_REG = rnode_3to4_bb3_add16_0_reg_4_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_arrayidx32_valid_out;
wire local_bb3_arrayidx32_stall_in;
wire local_bb3_arrayidx32_inputs_ready;
wire local_bb3_arrayidx32_stall_local;
wire [63:0] local_bb3_arrayidx32;

assign local_bb3_arrayidx32_inputs_ready = rnode_3to4_bb3_var__u17_0_valid_out_NO_SHIFT_REG;
assign local_bb3_arrayidx32 = ((input_gaussian & 64'hFFFFFFFFFFFFFC00) + (rnode_3to4_bb3_var__u17_0_NO_SHIFT_REG << 6'h2));
assign local_bb3_arrayidx32_valid_out = 1'b1;
assign rnode_3to4_bb3_var__u17_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u18_valid_out_1;
wire local_bb3_var__u18_stall_in_1;
wire local_bb3_notexit202_valid_out_0;
wire local_bb3_notexit202_stall_in_0;
wire local_bb3_notexit202_valid_out_1;
wire local_bb3_notexit202_stall_in_1;
wire local_bb3_indvars_iv_next27_valid_out_1;
wire local_bb3_indvars_iv_next27_stall_in_1;
wire local_bb3_notexit202_inputs_ready;
wire local_bb3_notexit202_stall_local;
wire local_bb3_notexit202;

assign local_bb3_notexit202_inputs_ready = (rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG & rnode_1to2_bb3_indvars_iv26_pop4__0_valid_out_0_NO_SHIFT_REG);
assign local_bb3_notexit202 = (local_bb3_var__u18 ^ 1'b1);
assign local_bb3_var__u18_valid_out_1 = 1'b1;
assign local_bb3_notexit202_valid_out_0 = 1'b1;
assign local_bb3_notexit202_valid_out_1 = 1'b1;
assign local_bb3_indvars_iv_next27_valid_out_1 = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_indvars_iv26_pop4__0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp1_i_stall_local;
wire local_bb3_cmp1_i;

assign local_bb3_cmp1_i = (rnode_3to4_bb3_add16_0_NO_SHIFT_REG > 32'h13F);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_arrayidx32_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_arrayidx32_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb3_arrayidx32_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_arrayidx32_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb3_arrayidx32_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_arrayidx32_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_arrayidx32_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_arrayidx32_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_arrayidx32_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_arrayidx32_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_arrayidx32_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_arrayidx32_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_arrayidx32_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in((local_bb3_arrayidx32 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_4to5_bb3_arrayidx32_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_arrayidx32_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_arrayidx32_0_reg_5_fifo.DATA_WIDTH = 64;
defparam rnode_4to5_bb3_arrayidx32_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_arrayidx32_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_arrayidx32_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_arrayidx32_stall_in = 1'b0;
assign rnode_4to5_bb3_arrayidx32_0_NO_SHIFT_REG = rnode_4to5_bb3_arrayidx32_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_arrayidx32_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_arrayidx32_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_var__u18_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u18_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u18_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u18_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u18_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u18_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u18_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u18_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_var__u18_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_var__u18_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_var__u18_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_var__u18_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_var__u18_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_var__u18),
	.data_out(rnode_2to3_bb3_var__u18_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_var__u18_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_var__u18_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_var__u18_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_var__u18_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_var__u18_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u18_stall_in_1 = 1'b0;
assign rnode_2to3_bb3_var__u18_0_NO_SHIFT_REG = rnode_2to3_bb3_var__u18_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_var__u18_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_var__u18_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb3_notexitcond201_notexit202_inputs_ready;
 reg local_bb3_notexitcond201_notexit202_valid_out_NO_SHIFT_REG;
wire local_bb3_notexitcond201_notexit202_stall_in;
wire local_bb3_notexitcond201_notexit202_output_regs_ready;
wire local_bb3_notexitcond201_notexit202_result;
wire local_bb3_notexitcond201_notexit202_fu_valid_out;
wire local_bb3_notexitcond201_notexit202_fu_stall_out;
 reg local_bb3_notexitcond201_notexit202_NO_SHIFT_REG;
wire local_bb3_notexitcond201_notexit202_causedstall;

acl_push local_bb3_notexitcond201_notexit202_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(local_bb3_notexit202),
	.stall_out(local_bb3_notexitcond201_notexit202_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notexitcond201_notexit202_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_notexitcond201_notexit202_result),
	.feedback_out(feedback_data_out_3),
	.feedback_valid_out(feedback_valid_out_3),
	.feedback_stall_in(feedback_stall_in_3)
);

defparam local_bb3_notexitcond201_notexit202_feedback.STALLFREE = 1;
defparam local_bb3_notexitcond201_notexit202_feedback.DATA_WIDTH = 1;
defparam local_bb3_notexitcond201_notexit202_feedback.FIFO_DEPTH = 1;
defparam local_bb3_notexitcond201_notexit202_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb3_notexitcond201_notexit202_feedback.STYLE = "REGULAR";

assign local_bb3_notexitcond201_notexit202_inputs_ready = 1'b1;
assign local_bb3_notexitcond201_notexit202_output_regs_ready = 1'b1;
assign local_bb3_notexit202_stall_in_0 = 1'b0;
assign SFC_1_VALID_1_2_0_stall_in_2 = 1'b0;
assign local_bb3_notexitcond201_notexit202_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_notexitcond201_notexit202_NO_SHIFT_REG <= 'x;
		local_bb3_notexitcond201_notexit202_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_notexitcond201_notexit202_output_regs_ready)
		begin
			local_bb3_notexitcond201_notexit202_NO_SHIFT_REG <= local_bb3_notexitcond201_notexit202_result;
			local_bb3_notexitcond201_notexit202_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_notexitcond201_notexit202_stall_in))
			begin
				local_bb3_notexitcond201_notexit202_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_indvars_iv26_push4_indvars_iv_next27_inputs_ready;
 reg local_bb3_indvars_iv26_push4_indvars_iv_next27_valid_out_NO_SHIFT_REG;
wire local_bb3_indvars_iv26_push4_indvars_iv_next27_stall_in;
wire local_bb3_indvars_iv26_push4_indvars_iv_next27_output_regs_ready;
wire [63:0] local_bb3_indvars_iv26_push4_indvars_iv_next27_result;
wire local_bb3_indvars_iv26_push4_indvars_iv_next27_fu_valid_out;
wire local_bb3_indvars_iv26_push4_indvars_iv_next27_fu_stall_out;
 reg [63:0] local_bb3_indvars_iv26_push4_indvars_iv_next27_NO_SHIFT_REG;
wire local_bb3_indvars_iv26_push4_indvars_iv_next27_causedstall;

acl_push local_bb3_indvars_iv26_push4_indvars_iv_next27_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexit202),
	.predicate(1'b0),
	.data_in(local_bb3_indvars_iv_next27),
	.stall_out(local_bb3_indvars_iv26_push4_indvars_iv_next27_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_indvars_iv26_push4_indvars_iv_next27_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_indvars_iv26_push4_indvars_iv_next27_result),
	.feedback_out(feedback_data_out_4),
	.feedback_valid_out(feedback_valid_out_4),
	.feedback_stall_in(feedback_stall_in_4)
);

defparam local_bb3_indvars_iv26_push4_indvars_iv_next27_feedback.STALLFREE = 1;
defparam local_bb3_indvars_iv26_push4_indvars_iv_next27_feedback.DATA_WIDTH = 64;
defparam local_bb3_indvars_iv26_push4_indvars_iv_next27_feedback.FIFO_DEPTH = 2;
defparam local_bb3_indvars_iv26_push4_indvars_iv_next27_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb3_indvars_iv26_push4_indvars_iv_next27_feedback.STYLE = "REGULAR";

assign local_bb3_indvars_iv26_push4_indvars_iv_next27_inputs_ready = 1'b1;
assign local_bb3_indvars_iv26_push4_indvars_iv_next27_output_regs_ready = 1'b1;
assign local_bb3_indvars_iv_next27_stall_in_1 = 1'b0;
assign local_bb3_notexit202_stall_in_1 = 1'b0;
assign SFC_1_VALID_1_2_0_stall_in_3 = 1'b0;
assign local_bb3_indvars_iv26_push4_indvars_iv_next27_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_indvars_iv26_push4_indvars_iv_next27_NO_SHIFT_REG <= 'x;
		local_bb3_indvars_iv26_push4_indvars_iv_next27_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_indvars_iv26_push4_indvars_iv_next27_output_regs_ready)
		begin
			local_bb3_indvars_iv26_push4_indvars_iv_next27_NO_SHIFT_REG <= local_bb3_indvars_iv26_push4_indvars_iv_next27_result;
			local_bb3_indvars_iv26_push4_indvars_iv_next27_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_indvars_iv26_push4_indvars_iv_next27_stall_in))
			begin
				local_bb3_indvars_iv26_push4_indvars_iv_next27_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_sub17_add16_valid_out;
wire local_bb3_sub17_add16_stall_in;
wire local_bb3_sub17_add16_inputs_ready;
wire local_bb3_sub17_add16_stall_local;
wire [31:0] local_bb3_sub17_add16;

assign local_bb3_sub17_add16_inputs_ready = (rnode_3to4_bb3_add16_0_valid_out_0_NO_SHIFT_REG & rnode_3to4_bb3_add16_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_sub17_add16 = (local_bb3_cmp1_i ? 32'h13F : rnode_3to4_bb3_add16_1_NO_SHIFT_REG);
assign local_bb3_sub17_add16_valid_out = 1'b1;
assign rnode_3to4_bb3_add16_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_add16_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_var__u18_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u18_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u18_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u18_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u18_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u18_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u18_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u18_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_var__u18_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_var__u18_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_var__u18_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_var__u18_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_var__u18_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(rnode_2to3_bb3_var__u18_0_NO_SHIFT_REG),
	.data_out(rnode_3to4_bb3_var__u18_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_var__u18_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_var__u18_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_var__u18_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_var__u18_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_var__u18_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_var__u18_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_var__u18_0_NO_SHIFT_REG = rnode_3to4_bb3_var__u18_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_var__u18_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_var__u18_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond201_notexit202_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb3_notexitcond201_notexit202_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb3_notexitcond201_notexit202_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb3_notexitcond201_notexit202_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_notexitcond201_notexit202_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notexitcond201_notexit202_stall_in = 1'b0;
assign rnode_3to5_bb3_notexitcond201_notexit202_0_NO_SHIFT_REG = rnode_3to5_bb3_notexitcond201_notexit202_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb3_notexitcond201_notexit202_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_notexitcond201_notexit202_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_indvars_iv26_push4_indvars_iv_next27_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_fifo.DATA_WIDTH = 64;
defparam rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_indvars_iv26_push4_indvars_iv_next27_stall_in = 1'b0;
assign rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_NO_SHIFT_REG = rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_sub17_add16_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_sub17_add16_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_sub17_add16_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_sub17_add16_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_sub17_add16_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_sub17_add16_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_sub17_add16_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_sub17_add16_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_sub17_add16_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_sub17_add16_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_sub17_add16_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_sub17_add16_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_sub17_add16_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_sub17_add16),
	.data_out(rnode_4to5_bb3_sub17_add16_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_sub17_add16_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_sub17_add16_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3_sub17_add16_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_sub17_add16_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_sub17_add16_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_sub17_add16_stall_in = 1'b0;
assign rnode_4to5_bb3_sub17_add16_0_NO_SHIFT_REG = rnode_4to5_bb3_sub17_add16_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_sub17_add16_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_sub17_add16_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_var__u18_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u18_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u18_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u18_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u18_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u18_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u18_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u18_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_var__u18_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_var__u18_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_var__u18_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_var__u18_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_var__u18_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_var__u18_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_var__u18_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_var__u18_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_var__u18_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_var__u18_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_var__u18_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_var__u18_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_var__u18_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_var__u18_0_NO_SHIFT_REG = rnode_4to5_bb3_var__u18_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_var__u18_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_var__u18_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi1_stall_local;
wire [191:0] local_bb3_c0_exi1;

assign local_bb3_c0_exi1[31:0] = 32'bx;
assign local_bb3_c0_exi1[63:32] = rnode_4to5_bb3_sub17_add16_0_NO_SHIFT_REG;
assign local_bb3_c0_exi1[191:64] = 128'bx;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi2_stall_local;
wire [191:0] local_bb3_c0_exi2;

assign local_bb3_c0_exi2[63:0] = local_bb3_c0_exi1[63:0];
assign local_bb3_c0_exi2[127:64] = (rnode_4to5_bb3_arrayidx32_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign local_bb3_c0_exi2[191:128] = local_bb3_c0_exi1[191:128];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi3_stall_local;
wire [191:0] local_bb3_c0_exi3;

assign local_bb3_c0_exi3[127:0] = local_bb3_c0_exi2[127:0];
assign local_bb3_c0_exi3[128] = rnode_4to5_bb3_var__u18_0_NO_SHIFT_REG;
assign local_bb3_c0_exi3[191:129] = local_bb3_c0_exi2[191:129];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi4_valid_out;
wire local_bb3_c0_exi4_stall_in;
wire local_bb3_c0_exi4_inputs_ready;
wire local_bb3_c0_exi4_stall_local;
wire [191:0] local_bb3_c0_exi4;

assign local_bb3_c0_exi4_inputs_ready = (rnode_3to5_bb3_notexitcond201_notexit202_0_valid_out_NO_SHIFT_REG & rnode_4to5_bb3_var__u18_0_valid_out_NO_SHIFT_REG & rnode_4to5_bb3_arrayidx32_0_valid_out_NO_SHIFT_REG & rnode_4to5_bb3_sub17_add16_0_valid_out_NO_SHIFT_REG);
assign local_bb3_c0_exi4[135:0] = local_bb3_c0_exi3[135:0];
assign local_bb3_c0_exi4[136] = rnode_3to5_bb3_notexitcond201_notexit202_0_NO_SHIFT_REG;
assign local_bb3_c0_exi4[191:137] = local_bb3_c0_exi3[191:137];
assign local_bb3_c0_exi4_valid_out = 1'b1;
assign rnode_3to5_bb3_notexitcond201_notexit202_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_var__u18_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_arrayidx32_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_sub17_add16_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb3_c0_exit_c0_exi4_inputs_ready;
 reg local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_0;
 reg local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_1;
 reg local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_2;
 reg local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_3;
 reg [191:0] local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG;
wire [191:0] local_bb3_c0_exit_c0_exi4_in;
wire local_bb3_c0_exit_c0_exi4_valid;
wire local_bb3_c0_exit_c0_exi4_causedstall;

acl_stall_free_sink local_bb3_c0_exit_c0_exi4_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb3_c0_exi4),
	.data_out(local_bb3_c0_exit_c0_exi4_in),
	.input_accepted(local_bb3_c0_enter_c0_eni1_input_accepted),
	.valid_out(local_bb3_c0_exit_c0_exi4_valid),
	.stall_in(~(local_bb3_c0_exit_c0_exi4_output_regs_ready)),
	.stall_entry(local_bb3_c0_exit_c0_exi4_entry_stall),
	.valid_in(local_bb3_c0_exit_c0_exi4_valid_in),
	.IIphases(local_bb3_c0_exit_c0_exi4_phases),
	.inc_pipelined_thread(local_bb3_c0_enter_c0_eni1_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb3_c0_enter_c0_eni1_dec_pipelined_thread)
);

defparam local_bb3_c0_exit_c0_exi4_instance.DATA_WIDTH = 192;
defparam local_bb3_c0_exit_c0_exi4_instance.PIPELINE_DEPTH = 9;
defparam local_bb3_c0_exit_c0_exi4_instance.SHARINGII = 1;
defparam local_bb3_c0_exit_c0_exi4_instance.SCHEDULEII = 1;
defparam local_bb3_c0_exit_c0_exi4_instance.ALWAYS_THROTTLE = 0;

assign local_bb3_c0_exit_c0_exi4_inputs_ready = 1'b1;
assign local_bb3_c0_exit_c0_exi4_output_regs_ready = ((~(local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_0)) & (~(local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_1)) & (~(local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_2)) & (~(local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_3)));
assign local_bb3_c0_exit_c0_exi4_valid_in = SFC_1_VALID_4_5_0_NO_SHIFT_REG;
assign local_bb3_c0_exi4_stall_in = 1'b0;
assign SFC_1_VALID_4_5_0_stall_in = 1'b0;
assign rnode_3to5_bb3_keep_going200_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_indvars_iv26_push4_indvars_iv_next27_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb3_c0_exit_c0_exi4_causedstall = (1'b1 && (1'b0 && !(~(local_bb3_c0_exit_c0_exi4_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG <= 'x;
		local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_c0_exit_c0_exi4_output_regs_ready)
		begin
			local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_in;
			local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
			local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
			local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
			local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
		end
		else
		begin
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_0))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_1))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_2))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_3))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe1_stall_local;
wire [31:0] local_bb3_c0_exe1;

assign local_bb3_c0_exe1 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe2_stall_local;
wire [63:0] local_bb3_c0_exe2;

assign local_bb3_c0_exe2 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[127:64];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe3_stall_local;
wire local_bb3_c0_exe3;

assign local_bb3_c0_exe3 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[128];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe4_valid_out;
wire local_bb3_c0_exe4_stall_in;
wire local_bb3_c0_exe3_valid_out;
wire local_bb3_c0_exe3_stall_in;
wire local_bb3_c0_exe2_valid_out;
wire local_bb3_c0_exe2_stall_in;
wire local_bb3_c0_exe1_valid_out;
wire local_bb3_c0_exe1_stall_in;
wire local_bb3_c0_exe4_inputs_ready;
wire local_bb3_c0_exe4_stall_local;
wire local_bb3_c0_exe4;

assign local_bb3_c0_exe4_inputs_ready = (local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG);
assign local_bb3_c0_exe4 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[136];
assign local_bb3_c0_exe4_stall_local = (local_bb3_c0_exe4_stall_in | local_bb3_c0_exe3_stall_in | local_bb3_c0_exe2_stall_in | local_bb3_c0_exe1_stall_in);
assign local_bb3_c0_exe4_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exe3_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exe2_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exe1_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exit_c0_exi4_stall_in_3 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));
assign local_bb3_c0_exit_c0_exi4_stall_in_2 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));
assign local_bb3_c0_exit_c0_exi4_stall_in_1 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));
assign local_bb3_c0_exit_c0_exi4_stall_in_0 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [31:0] lvb_bb3_c0_exe1_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb3_c0_exe2_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe3_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe4_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_t_219_pop5__reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_sum_218_pop6__reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb3_sum_218_pop6__valid_out_NO_SHIFT_REG & local_bb3_t_219_pop5__valid_out_NO_SHIFT_REG & local_bb3_c0_exe4_valid_out & local_bb3_c0_exe3_valid_out & local_bb3_c0_exe2_valid_out & local_bb3_c0_exe1_valid_out);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb3_sum_218_pop6__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_t_219_pop5__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe4_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe3_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb3_c0_exe1 = lvb_bb3_c0_exe1_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe2 = lvb_bb3_c0_exe2_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe3 = lvb_bb3_c0_exe3_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe4 = lvb_bb3_c0_exe4_reg_NO_SHIFT_REG;
assign lvb_bb3_t_219_pop5_ = lvb_bb3_t_219_pop5__reg_NO_SHIFT_REG;
assign lvb_bb3_sum_218_pop6_ = lvb_bb3_sum_218_pop6__reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb3_c0_exe1_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe2_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe3_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe4_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_t_219_pop5__reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_sum_218_pop6__reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb3_c0_exe1_reg_NO_SHIFT_REG <= local_bb3_c0_exe1;
			lvb_bb3_c0_exe2_reg_NO_SHIFT_REG <= (local_bb3_c0_exe2 & 64'hFFFFFFFFFFFFFFFC);
			lvb_bb3_c0_exe3_reg_NO_SHIFT_REG <= local_bb3_c0_exe3;
			lvb_bb3_c0_exe4_reg_NO_SHIFT_REG <= local_bb3_c0_exe4;
			lvb_bb3_t_219_pop5__reg_NO_SHIFT_REG <= local_bb3_t_219_pop5__NO_SHIFT_REG;
			lvb_bb3_sum_218_pop6__reg_NO_SHIFT_REG <= local_bb3_sum_218_pop6__NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_4
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_in,
		input [63:0] 		input_gaussian,
		input [31:0] 		input_r,
		input 		input_wii_cmp1017,
		input [31:0] 		input_wii_mul39,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u19,
		input 		valid_in_0,
		output 		stall_out_0,
		input [31:0] 		input_t_313_0,
		input [31:0] 		input_sum_312_0,
		input 		input_forked203_0,
		input [31:0] 		input_sub17_add16204_0,
		input [63:0] 		input_arrayidx32205_0,
		input 		input_var__u20_0,
		input 		input_notexitcond201206_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [31:0] 		input_t_313_1,
		input [31:0] 		input_sum_312_1,
		input 		input_forked203_1,
		input [31:0] 		input_sub17_add16204_1,
		input [63:0] 		input_arrayidx32205_1,
		input 		input_var__u20_1,
		input 		input_notexitcond201206_1,
		output 		valid_out_0,
		input 		stall_in_0,
		output [319:0] 		lvb_bb4_c0_exit214_c0_exi7_0,
		output 		lvb_bb4_c0_exe7_0,
		output [95:0] 		lvb_bb4_c1_exit_c1_exi2_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [319:0] 		lvb_bb4_c0_exit214_c0_exi7_1,
		output 		lvb_bb4_c0_exe7_1,
		output [95:0] 		lvb_bb4_c1_exit_c1_exi2_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		ffwd_10_0,
		input [31:0] 		ffwd_1_0,
		input 		feedback_valid_in_7,
		output 		feedback_stall_out_7,
		input [63:0] 		feedback_data_in_7,
		output 		feedback_stall_out_0,
		input 		feedback_valid_in_1,
		output 		feedback_stall_out_1,
		input 		feedback_data_in_1,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		input 		feedback_valid_in_10,
		output 		feedback_stall_out_10,
		input [31:0] 		feedback_data_in_10,
		input 		feedback_valid_in_11,
		output 		feedback_stall_out_11,
		input [63:0] 		feedback_data_in_11,
		input 		feedback_valid_in_12,
		output 		feedback_stall_out_12,
		input 		feedback_data_in_12,
		input 		feedback_valid_in_13,
		output 		feedback_stall_out_13,
		input 		feedback_data_in_13,
		output 		feedback_valid_out_1,
		input 		feedback_stall_in_1,
		output 		feedback_data_out_1,
		output 		feedback_valid_out_7,
		input 		feedback_stall_in_7,
		output [63:0] 		feedback_data_out_7,
		output 		feedback_valid_out_11,
		input 		feedback_stall_in_11,
		output [63:0] 		feedback_data_out_11,
		output 		feedback_valid_out_12,
		input 		feedback_stall_in_12,
		output 		feedback_data_out_12,
		output 		feedback_valid_out_13,
		input 		feedback_stall_in_13,
		output 		feedback_data_out_13,
		output 		feedback_valid_out_10,
		input 		feedback_stall_in_10,
		output [31:0] 		feedback_data_out_10,
		input [511:0] 		avm_local_bb4_ld__readdata,
		input 		avm_local_bb4_ld__readdatavalid,
		input 		avm_local_bb4_ld__waitrequest,
		output [32:0] 		avm_local_bb4_ld__address,
		output 		avm_local_bb4_ld__read,
		output 		avm_local_bb4_ld__write,
		input 		avm_local_bb4_ld__writeack,
		output [511:0] 		avm_local_bb4_ld__writedata,
		output [63:0] 		avm_local_bb4_ld__byteenable,
		output [4:0] 		avm_local_bb4_ld__burstcount,
		output 		local_bb4_ld__active,
		input 		clock2x,
		input [511:0] 		avm_local_bb4_ld__u28_readdata,
		input 		avm_local_bb4_ld__u28_readdatavalid,
		input 		avm_local_bb4_ld__u28_waitrequest,
		output [32:0] 		avm_local_bb4_ld__u28_address,
		output 		avm_local_bb4_ld__u28_read,
		output 		avm_local_bb4_ld__u28_write,
		input 		avm_local_bb4_ld__u28_writeack,
		output [511:0] 		avm_local_bb4_ld__u28_writedata,
		output [63:0] 		avm_local_bb4_ld__u28_byteenable,
		output [4:0] 		avm_local_bb4_ld__u28_burstcount,
		output 		local_bb4_ld__u28_active,
		input [511:0] 		avm_local_bb4_ld__u29_readdata,
		input 		avm_local_bb4_ld__u29_readdatavalid,
		input 		avm_local_bb4_ld__u29_waitrequest,
		output [32:0] 		avm_local_bb4_ld__u29_address,
		output 		avm_local_bb4_ld__u29_read,
		output 		avm_local_bb4_ld__u29_write,
		input 		avm_local_bb4_ld__u29_writeack,
		output [511:0] 		avm_local_bb4_ld__u29_writedata,
		output [63:0] 		avm_local_bb4_ld__u29_byteenable,
		output [4:0] 		avm_local_bb4_ld__u29_burstcount,
		output 		local_bb4_ld__u29_active,
		input [31:0] 		ffwd_8_0,
		input 		feedback_valid_in_9,
		output 		feedback_stall_out_9,
		input [31:0] 		feedback_data_in_9,
		input 		feedback_valid_in_8,
		output 		feedback_stall_out_8,
		input [31:0] 		feedback_data_in_8,
		output 		feedback_valid_out_9,
		input 		feedback_stall_in_9,
		output [31:0] 		feedback_data_out_9,
		output [31:0] 		ffwd_11_0,
		output 		feedback_valid_out_8,
		input 		feedback_stall_in_8,
		output [31:0] 		feedback_data_out_8,
		output [31:0] 		ffwd_12_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_313_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_312_0_staging_reg_NO_SHIFT_REG;
 reg input_forked203_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sub17_add16204_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_arrayidx32205_0_staging_reg_NO_SHIFT_REG;
 reg input_var__u20_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond201206_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_t_313_NO_SHIFT_REG;
 reg [31:0] local_lvm_sum_312_NO_SHIFT_REG;
 reg local_lvm_forked203_NO_SHIFT_REG;
 reg [31:0] local_lvm_sub17_add16204_NO_SHIFT_REG;
 reg [63:0] local_lvm_arrayidx32205_NO_SHIFT_REG;
 reg local_lvm_var__u20_NO_SHIFT_REG;
 reg local_lvm_notexitcond201206_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_313_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_312_1_staging_reg_NO_SHIFT_REG;
 reg input_forked203_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sub17_add16204_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_arrayidx32205_1_staging_reg_NO_SHIFT_REG;
 reg input_var__u20_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond201206_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_t_313_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_312_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_forked203_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_sub17_add16204_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_arrayidx32205_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u20_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond201206_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_t_313_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_312_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_forked203_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_sub17_add16204_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_arrayidx32205_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u20_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond201206_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_t_313_0_staging_reg_NO_SHIFT_REG <= input_t_313_0;
				input_sum_312_0_staging_reg_NO_SHIFT_REG <= input_sum_312_0;
				input_forked203_0_staging_reg_NO_SHIFT_REG <= input_forked203_0;
				input_sub17_add16204_0_staging_reg_NO_SHIFT_REG <= input_sub17_add16204_0;
				input_arrayidx32205_0_staging_reg_NO_SHIFT_REG <= input_arrayidx32205_0;
				input_var__u20_0_staging_reg_NO_SHIFT_REG <= input_var__u20_0;
				input_notexitcond201206_0_staging_reg_NO_SHIFT_REG <= input_notexitcond201206_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_t_313_1_staging_reg_NO_SHIFT_REG <= input_t_313_1;
				input_sum_312_1_staging_reg_NO_SHIFT_REG <= input_sum_312_1;
				input_forked203_1_staging_reg_NO_SHIFT_REG <= input_forked203_1;
				input_sub17_add16204_1_staging_reg_NO_SHIFT_REG <= input_sub17_add16204_1;
				input_arrayidx32205_1_staging_reg_NO_SHIFT_REG <= input_arrayidx32205_1;
				input_var__u20_1_staging_reg_NO_SHIFT_REG <= input_var__u20_1;
				input_notexitcond201206_1_staging_reg_NO_SHIFT_REG <= input_notexitcond201206_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_t_313_NO_SHIFT_REG <= input_t_313_0_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_312_NO_SHIFT_REG <= input_sum_312_0_staging_reg_NO_SHIFT_REG;
					local_lvm_forked203_NO_SHIFT_REG <= input_forked203_0_staging_reg_NO_SHIFT_REG;
					local_lvm_sub17_add16204_NO_SHIFT_REG <= input_sub17_add16204_0_staging_reg_NO_SHIFT_REG;
					local_lvm_arrayidx32205_NO_SHIFT_REG <= input_arrayidx32205_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond201206_NO_SHIFT_REG <= input_notexitcond201206_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_t_313_NO_SHIFT_REG <= input_t_313_0;
					local_lvm_sum_312_NO_SHIFT_REG <= input_sum_312_0;
					local_lvm_forked203_NO_SHIFT_REG <= input_forked203_0;
					local_lvm_sub17_add16204_NO_SHIFT_REG <= input_sub17_add16204_0;
					local_lvm_arrayidx32205_NO_SHIFT_REG <= input_arrayidx32205_0;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_0;
					local_lvm_notexitcond201206_NO_SHIFT_REG <= input_notexitcond201206_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_t_313_NO_SHIFT_REG <= input_t_313_1_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_312_NO_SHIFT_REG <= input_sum_312_1_staging_reg_NO_SHIFT_REG;
					local_lvm_forked203_NO_SHIFT_REG <= input_forked203_1_staging_reg_NO_SHIFT_REG;
					local_lvm_sub17_add16204_NO_SHIFT_REG <= input_sub17_add16204_1_staging_reg_NO_SHIFT_REG;
					local_lvm_arrayidx32205_NO_SHIFT_REG <= input_arrayidx32205_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond201206_NO_SHIFT_REG <= input_notexitcond201206_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_t_313_NO_SHIFT_REG <= input_t_313_1;
					local_lvm_sum_312_NO_SHIFT_REG <= input_sum_312_1;
					local_lvm_forked203_NO_SHIFT_REG <= input_forked203_1;
					local_lvm_sub17_add16204_NO_SHIFT_REG <= input_sub17_add16204_1;
					local_lvm_arrayidx32205_NO_SHIFT_REG <= input_arrayidx32205_1;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_1;
					local_lvm_notexitcond201206_NO_SHIFT_REG <= input_notexitcond201206_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni1207_stall_local;
wire [191:0] local_bb4_c0_eni1207;

assign local_bb4_c0_eni1207[7:0] = 8'bx;
assign local_bb4_c0_eni1207[8] = local_lvm_forked203_NO_SHIFT_REG;
assign local_bb4_c0_eni1207[191:9] = 183'bx;

// Register node:
//  * latency = 14
//  * capacity = 14
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_fifo.DEPTH = 15;
defparam rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_fifo.IMPL = "ram";

assign rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_reg_15_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign merge_node_stall_in_5 = rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_out_reg_15_NO_SHIFT_REG;
assign rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_in_reg_15_NO_SHIFT_REG = rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_in_NO_SHIFT_REG;
assign rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_valid_out_NO_SHIFT_REG = rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_valid_out_reg_15_NO_SHIFT_REG;

// Register node:
//  * latency = 177
//  * capacity = 177
 logic rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_out_reg_178_NO_SHIFT_REG;
wire [64:0] rci_rcnode_1to338_rc7_t_313_0_reg_1;

acl_data_fifo rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_fifo.DEPTH = 178;
defparam rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_fifo.DATA_WIDTH = 0;
defparam rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_fifo.IMPL = "ram";

assign rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_reg_178_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_6_NO_SHIFT_REG;
assign merge_node_stall_in_6 = rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_out_reg_178_NO_SHIFT_REG;
assign rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_reg_178_NO_SHIFT_REG = rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_NO_SHIFT_REG;
assign rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_NO_SHIFT_REG = rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_reg_178_NO_SHIFT_REG;
assign rci_rcnode_1to338_rc7_t_313_0_reg_1[31:0] = local_lvm_t_313_NO_SHIFT_REG;
assign rci_rcnode_1to338_rc7_t_313_0_reg_1[32] = local_lvm_forked203_NO_SHIFT_REG;
assign rci_rcnode_1to338_rc7_t_313_0_reg_1[64:33] = local_lvm_sum_312_NO_SHIFT_REG;

// Register node:
//  * latency = 337
//  * capacity = 337
 logic rcnode_1to338_rc7_t_313_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to338_rc7_t_313_0_stall_in_NO_SHIFT_REG;
 logic [64:0] rcnode_1to338_rc7_t_313_0_NO_SHIFT_REG;
 logic rcnode_1to338_rc7_t_313_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [64:0] rcnode_1to338_rc7_t_313_0_reg_338_NO_SHIFT_REG;
 logic rcnode_1to338_rc7_t_313_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rcnode_1to338_rc7_t_313_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rcnode_1to338_rc7_t_313_0_stall_out_reg_338_IP_NO_SHIFT_REG;
 logic rcnode_1to338_rc7_t_313_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rcnode_1to338_rc7_t_313_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to338_rc7_t_313_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to338_rc7_t_313_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rcnode_1to338_rc7_t_313_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rcnode_1to338_rc7_t_313_0_stall_out_reg_338_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to338_rc7_t_313_0_reg_1),
	.data_out(rcnode_1to338_rc7_t_313_0_reg_338_NO_SHIFT_REG)
);

defparam rcnode_1to338_rc7_t_313_0_reg_338_fifo.DEPTH = 338;
defparam rcnode_1to338_rc7_t_313_0_reg_338_fifo.DATA_WIDTH = 65;
defparam rcnode_1to338_rc7_t_313_0_reg_338_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to338_rc7_t_313_0_reg_338_fifo.IMPL = "ram";

assign rcnode_1to338_rc7_t_313_0_reg_338_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_7_NO_SHIFT_REG;
assign rcnode_1to338_rc7_t_313_0_stall_out_reg_338_NO_SHIFT_REG = (~(rcnode_1to338_rc7_t_313_0_reg_338_inputs_ready_NO_SHIFT_REG) | rcnode_1to338_rc7_t_313_0_stall_out_reg_338_IP_NO_SHIFT_REG);
assign merge_node_stall_in_7 = rcnode_1to338_rc7_t_313_0_stall_out_reg_338_NO_SHIFT_REG;
assign rcnode_1to338_rc7_t_313_0_NO_SHIFT_REG = rcnode_1to338_rc7_t_313_0_reg_338_NO_SHIFT_REG;
assign rcnode_1to338_rc7_t_313_0_stall_in_reg_338_NO_SHIFT_REG = rcnode_1to338_rc7_t_313_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to338_rc7_t_313_0_valid_out_NO_SHIFT_REG = rcnode_1to338_rc7_t_313_0_valid_out_reg_338_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni2_stall_local;
wire [191:0] local_bb4_c0_eni2;

assign local_bb4_c0_eni2[31:0] = local_bb4_c0_eni1207[31:0];
assign local_bb4_c0_eni2[63:32] = local_lvm_sub17_add16204_NO_SHIFT_REG;
assign local_bb4_c0_eni2[191:64] = local_bb4_c0_eni1207[191:64];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_fifo.DEPTH = 2;
defparam rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_fifo.IMPL = "ll_reg";

assign rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_reg_16_inputs_ready_NO_SHIFT_REG = rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_valid_out_NO_SHIFT_REG;
assign rnode_1to15_bb4__acl_ffwd_dest_i1_10_0_stall_in_NO_SHIFT_REG = rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_out_reg_16_NO_SHIFT_REG;
assign rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_in_reg_16_NO_SHIFT_REG = rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_in_NO_SHIFT_REG;
assign rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_valid_out_NO_SHIFT_REG = rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_valid_out_reg_16_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_fifo.DATA_WIDTH = 0;
defparam rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_fifo.IMPL = "ll_reg";

assign rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_reg_179_inputs_ready_NO_SHIFT_REG = rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_NO_SHIFT_REG;
assign rnode_1to178_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_NO_SHIFT_REG = rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_out_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_reg_179_NO_SHIFT_REG = rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_NO_SHIFT_REG;
assign rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_NO_SHIFT_REG = rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_reg_179_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni3_stall_local;
wire [191:0] local_bb4_c0_eni3;

assign local_bb4_c0_eni3[63:0] = local_bb4_c0_eni2[63:0];
assign local_bb4_c0_eni3[127:64] = local_lvm_arrayidx32205_NO_SHIFT_REG;
assign local_bb4_c0_eni3[191:128] = local_bb4_c0_eni2[191:128];

// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_i1_10_valid_out;
wire local_bb4__acl_ffwd_dest_i1_10_stall_in;
wire local_bb4__acl_ffwd_dest_i1_10_inputs_ready;
wire local_bb4__acl_ffwd_dest_i1_10_stall_local;
wire local_bb4__acl_ffwd_dest_i1_10;

assign local_bb4__acl_ffwd_dest_i1_10_inputs_ready = rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_valid_out_NO_SHIFT_REG;
assign local_bb4__acl_ffwd_dest_i1_10 = ffwd_10_0;
assign local_bb4__acl_ffwd_dest_i1_10_valid_out = local_bb4__acl_ffwd_dest_i1_10_inputs_ready;
assign local_bb4__acl_ffwd_dest_i1_10_stall_local = local_bb4__acl_ffwd_dest_i1_10_stall_in;
assign rnode_15to16_bb4__acl_ffwd_dest_i1_10_0_stall_in_NO_SHIFT_REG = (|local_bb4__acl_ffwd_dest_i1_10_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_i1_10_u21_stall_local;
wire local_bb4__acl_ffwd_dest_i1_10_u21;

assign local_bb4__acl_ffwd_dest_i1_10_u21 = ffwd_10_0;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni4_stall_local;
wire [191:0] local_bb4_c0_eni4;

assign local_bb4_c0_eni4[127:0] = local_bb4_c0_eni3[127:0];
assign local_bb4_c0_eni4[128] = local_lvm_var__u20_NO_SHIFT_REG;
assign local_bb4_c0_eni4[191:129] = local_bb4_c0_eni3[191:129];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni5_stall_local;
wire [191:0] local_bb4_c0_eni5;

assign local_bb4_c0_eni5[135:0] = local_bb4_c0_eni4[135:0];
assign local_bb4_c0_eni5[136] = local_lvm_notexitcond201206_NO_SHIFT_REG;
assign local_bb4_c0_eni5[191:137] = local_bb4_c0_eni4[191:137];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene1209_valid_out;
wire local_bb4_c0_ene1209_stall_in;
wire local_bb4_c0_ene2_valid_out;
wire local_bb4_c0_ene2_stall_in;
wire local_bb4_c0_ene3_valid_out;
wire local_bb4_c0_ene3_stall_in;
wire local_bb4_c0_ene4_valid_out;
wire local_bb4_c0_ene4_stall_in;
wire local_bb4_c0_ene5_valid_out;
wire local_bb4_c0_ene5_stall_in;
wire SFC_2_VALID_1_1_0_valid_out;
wire SFC_2_VALID_1_1_0_stall_in;
wire local_bb4_c0_enter208_c0_eni5_inputs_ready;
wire local_bb4_c0_enter208_c0_eni5_stall_local;
wire local_bb4_c0_enter208_c0_eni5_input_accepted;
wire [191:0] local_bb4_c0_enter208_c0_eni5;
wire local_bb4_c0_exit214_c0_exi7_entry_stall;
wire local_bb4_c0_enter208_c0_eni5_valid_bit;
wire local_bb4_c0_exit214_c0_exi7_output_regs_ready;
wire local_bb4_c0_exit214_c0_exi7_valid_in;
wire local_bb4_c0_exit214_c0_exi7_phases;
wire local_bb4_c0_enter208_c0_eni5_inc_pipelined_thread;
wire local_bb4_c0_enter208_c0_eni5_dec_pipelined_thread;
wire local_bb4_c0_enter208_c0_eni5_fu_stall_out;

assign local_bb4_c0_enter208_c0_eni5_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_3_NO_SHIFT_REG & merge_node_valid_out_4_NO_SHIFT_REG);
assign local_bb4_c0_enter208_c0_eni5 = local_bb4_c0_eni5;
assign local_bb4_c0_enter208_c0_eni5_input_accepted = (local_bb4_c0_enter208_c0_eni5_inputs_ready && !(local_bb4_c0_exit214_c0_exi7_entry_stall));
assign local_bb4_c0_enter208_c0_eni5_valid_bit = local_bb4_c0_enter208_c0_eni5_input_accepted;
assign local_bb4_c0_enter208_c0_eni5_inc_pipelined_thread = 1'b1;
assign local_bb4_c0_enter208_c0_eni5_dec_pipelined_thread = ~(1'b0);
assign local_bb4_c0_enter208_c0_eni5_fu_stall_out = (~(local_bb4_c0_enter208_c0_eni5_inputs_ready) | local_bb4_c0_exit214_c0_exi7_entry_stall);
assign local_bb4_c0_enter208_c0_eni5_stall_local = (local_bb4_c0_ene1209_stall_in | local_bb4_c0_ene2_stall_in | local_bb4_c0_ene3_stall_in | local_bb4_c0_ene4_stall_in | local_bb4_c0_ene5_stall_in | SFC_2_VALID_1_1_0_stall_in);
assign local_bb4_c0_ene1209_valid_out = local_bb4_c0_enter208_c0_eni5_inputs_ready;
assign local_bb4_c0_ene2_valid_out = local_bb4_c0_enter208_c0_eni5_inputs_ready;
assign local_bb4_c0_ene3_valid_out = local_bb4_c0_enter208_c0_eni5_inputs_ready;
assign local_bb4_c0_ene4_valid_out = local_bb4_c0_enter208_c0_eni5_inputs_ready;
assign local_bb4_c0_ene5_valid_out = local_bb4_c0_enter208_c0_eni5_inputs_ready;
assign SFC_2_VALID_1_1_0_valid_out = local_bb4_c0_enter208_c0_eni5_inputs_ready;
assign merge_node_stall_in_0 = (local_bb4_c0_enter208_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter208_c0_eni5_inputs_ready));
assign merge_node_stall_in_1 = (local_bb4_c0_enter208_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter208_c0_eni5_inputs_ready));
assign merge_node_stall_in_2 = (local_bb4_c0_enter208_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter208_c0_eni5_inputs_ready));
assign merge_node_stall_in_3 = (local_bb4_c0_enter208_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter208_c0_eni5_inputs_ready));
assign merge_node_stall_in_4 = (local_bb4_c0_enter208_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter208_c0_eni5_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene1209_stall_local;
wire local_bb4_c0_ene1209;

assign local_bb4_c0_ene1209 = local_bb4_c0_enter208_c0_eni5[8];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene2_stall_local;
wire [31:0] local_bb4_c0_ene2;

assign local_bb4_c0_ene2 = local_bb4_c0_enter208_c0_eni5[63:32];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene3_stall_local;
wire [63:0] local_bb4_c0_ene3;

assign local_bb4_c0_ene3 = local_bb4_c0_enter208_c0_eni5[127:64];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene4_stall_local;
wire local_bb4_c0_ene4;

assign local_bb4_c0_ene4 = local_bb4_c0_enter208_c0_eni5[128];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene5_stall_local;
wire local_bb4_c0_ene5;

assign local_bb4_c0_ene5 = local_bb4_c0_enter208_c0_eni5[136];

// This section implements an unregistered operation.
// 
wire SFC_2_VALID_1_1_0_stall_local;
wire SFC_2_VALID_1_1_0;

assign SFC_2_VALID_1_1_0 = local_bb4_c0_enter208_c0_eni5_valid_bit;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene1209_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1209_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1209_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1209_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1209_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1209_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1209_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1209_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene1209_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene1209_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene1209_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene1209_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene1209_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene1209),
	.data_out(rnode_1to2_bb4_c0_ene1209_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene1209_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene1209_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene1209_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene1209_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene1209_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene1209_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene1209_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene1209_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene1209_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene1209_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene2_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene2_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene2_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene2_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene2_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene2_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene2),
	.data_out(rnode_1to2_bb4_c0_ene2_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene2_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene2_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene2_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene2_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene2_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb4_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb4_c0_ene3_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene3_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene3_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene3_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene3_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene3_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene3),
	.data_out(rnode_1to2_bb4_c0_ene3_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.DATA_WIDTH = 64;
defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene3_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene3_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene3_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene3_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene3_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene4_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene4_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene4_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene4_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene4_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene4),
	.data_out(rnode_1to2_bb4_c0_ene4_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene4_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene4_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene4_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene4_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene4_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene5_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene5_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene5_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene5_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene5_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene5),
	.data_out(rnode_1to2_bb4_c0_ene5_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene5_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene5_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene5_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene5_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene5_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_1_2_0_inputs_ready;
 reg SFC_2_VALID_1_2_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_1_2_0_stall_in;
wire SFC_2_VALID_1_2_0_output_regs_ready;
 reg SFC_2_VALID_1_2_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_1_2_0_causedstall;

assign SFC_2_VALID_1_2_0_inputs_ready = 1'b1;
assign SFC_2_VALID_1_2_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_1_1_0_stall_in = 1'b0;
assign SFC_2_VALID_1_2_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_1_2_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_1_2_0_output_regs_ready)
		begin
			SFC_2_VALID_1_2_0_NO_SHIFT_REG <= SFC_2_VALID_1_1_0;
		end
	end
end


// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_2to6_bb4_c0_ene1209_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene1209_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene1209_0_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene1209_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene1209_0_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene1209_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene1209_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene1209_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_2to6_bb4_c0_ene1209_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to6_bb4_c0_ene1209_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to6_bb4_c0_ene1209_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_2to6_bb4_c0_ene1209_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_2to6_bb4_c0_ene1209_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene1209_0_NO_SHIFT_REG),
	.data_out(rnode_2to6_bb4_c0_ene1209_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_2to6_bb4_c0_ene1209_0_reg_6_fifo.DEPTH = 4;
defparam rnode_2to6_bb4_c0_ene1209_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_2to6_bb4_c0_ene1209_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to6_bb4_c0_ene1209_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_2to6_bb4_c0_ene1209_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene1209_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to6_bb4_c0_ene1209_0_NO_SHIFT_REG = rnode_2to6_bb4_c0_ene1209_0_reg_6_NO_SHIFT_REG;
assign rnode_2to6_bb4_c0_ene1209_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_2to6_bb4_c0_ene1209_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_2to8_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to8_bb4_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to8_bb4_c0_ene2_0_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_2to8_bb4_c0_ene2_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to8_bb4_c0_ene2_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to8_bb4_c0_ene2_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_2to8_bb4_c0_ene2_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_2to8_bb4_c0_ene2_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_2to8_bb4_c0_ene2_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.DEPTH = 6;
defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_2to8_bb4_c0_ene2_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene2_0_NO_SHIFT_REG = rnode_2to8_bb4_c0_ene2_0_reg_8_NO_SHIFT_REG;
assign rnode_2to8_bb4_c0_ene2_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_2to9_bb4_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene3_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_2to9_bb4_c0_ene3_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene3_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene3_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene3_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene3_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene3_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene3_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene3_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene3_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene3_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene3_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene3_0_reg_9_fifo.DATA_WIDTH = 64;
defparam rnode_2to9_bb4_c0_ene3_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene3_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene3_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene3_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene3_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene3_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene4_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene4_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene4_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene4_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene4_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene4_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene4_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene4_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene4_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene4_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene5_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene5_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene5_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene5_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene5_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene5_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene5_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene5_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene5_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene5_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_2_3_0_inputs_ready;
 reg SFC_2_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_2_3_0_stall_in;
wire SFC_2_VALID_2_3_0_output_regs_ready;
 reg SFC_2_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_2_3_0_causedstall;

assign SFC_2_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_1_2_0_stall_in = 1'b0;
assign SFC_2_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_2_3_0_output_regs_ready)
		begin
			SFC_2_VALID_2_3_0_NO_SHIFT_REG <= SFC_2_VALID_1_2_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_1_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_2_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_valid_out_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_stall_in_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene1209_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_c0_ene1209_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_c0_ene1209_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_c0_ene1209_0_stall_in_0_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_c0_ene1209_0_valid_out_0_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_c0_ene1209_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(rnode_2to6_bb4_c0_ene1209_0_NO_SHIFT_REG),
	.data_out(rnode_6to7_bb4_c0_ene1209_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_c0_ene1209_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_c0_ene1209_0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_6to7_bb4_c0_ene1209_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_c0_ene1209_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_c0_ene1209_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to6_bb4_c0_ene1209_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene1209_0_stall_in_0_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene1209_0_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene1209_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene1209_1_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene1209_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene1209_2_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene1209_0_reg_7_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_c0_ene2_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_c0_ene2_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_c0_ene2_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_c0_ene2_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_c0_ene2_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_c0_ene2_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_2to8_bb4_c0_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_c0_ene2_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_c0_ene2_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to8_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene2_0_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene2_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_c0_ene2_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_9to10_bb4_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene3_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_9to10_bb4_c0_ene3_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene3_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene3_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene3_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene3_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene3_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene3_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene3_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene3_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene3_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene3_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene3_0_reg_10_fifo.DATA_WIDTH = 64;
defparam rnode_9to10_bb4_c0_ene3_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene3_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene3_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene3_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene3_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene3_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene4_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene4_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene4_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene4_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene4_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene4_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene4_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene4_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene4_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene4_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene5_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene5_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene5_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene5_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene5_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene5_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene5_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene5_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene5_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene5_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_3_4_0_inputs_ready;
 reg SFC_2_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_3_4_0_stall_in;
wire SFC_2_VALID_3_4_0_output_regs_ready;
 reg SFC_2_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_3_4_0_causedstall;

assign SFC_2_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_stall_in = 1'b0;
assign SFC_2_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_3_4_0_output_regs_ready)
		begin
			SFC_2_VALID_3_4_0_NO_SHIFT_REG <= SFC_2_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_i32_1_stall_local;
wire [31:0] local_bb4__acl_ffwd_dest_i32_1;

assign local_bb4__acl_ffwd_dest_i32_1 = ffwd_1_0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_7to9_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_1_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_2_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_3_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_valid_out_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_stall_in_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene1209_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_7to9_bb4_c0_ene1209_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to9_bb4_c0_ene1209_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to9_bb4_c0_ene1209_0_stall_in_0_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_7to9_bb4_c0_ene1209_0_valid_out_0_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_7to9_bb4_c0_ene1209_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_c0_ene1209_2_NO_SHIFT_REG),
	.data_out(rnode_7to9_bb4_c0_ene1209_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_7to9_bb4_c0_ene1209_0_reg_9_fifo.DEPTH = 2;
defparam rnode_7to9_bb4_c0_ene1209_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_7to9_bb4_c0_ene1209_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to9_bb4_c0_ene1209_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_7to9_bb4_c0_ene1209_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene1209_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_7to9_bb4_c0_ene1209_0_stall_in_0_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_7to9_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene1209_0_NO_SHIFT_REG = rnode_7to9_bb4_c0_ene1209_0_reg_9_NO_SHIFT_REG;
assign rnode_7to9_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene1209_1_NO_SHIFT_REG = rnode_7to9_bb4_c0_ene1209_0_reg_9_NO_SHIFT_REG;
assign rnode_7to9_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene1209_2_NO_SHIFT_REG = rnode_7to9_bb4_c0_ene1209_0_reg_9_NO_SHIFT_REG;
assign rnode_7to9_bb4_c0_ene1209_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene1209_3_NO_SHIFT_REG = rnode_7to9_bb4_c0_ene1209_0_reg_9_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_2_VALID_4_5_0_inputs_ready;
 reg SFC_2_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_4_5_0_stall_in;
wire SFC_2_VALID_4_5_0_output_regs_ready;
 reg SFC_2_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_4_5_0_causedstall;

assign SFC_2_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_stall_in = 1'b0;
assign SFC_2_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_4_5_0_output_regs_ready)
		begin
			SFC_2_VALID_4_5_0_NO_SHIFT_REG <= SFC_2_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_i1_10_u22_stall_local;
wire local_bb4__acl_ffwd_dest_i1_10_u22;

assign local_bb4__acl_ffwd_dest_i1_10_u22 = ffwd_10_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_2_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_valid_out_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_stall_in_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1209_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene1209_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene1209_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene1209_0_stall_in_0_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene1209_0_valid_out_0_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene1209_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_7to9_bb4_c0_ene1209_3_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene1209_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene1209_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene1209_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene1209_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene1209_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene1209_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene1209_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1209_0_stall_in_0_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene1209_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene1209_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene1209_1_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene1209_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene1209_2_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene1209_0_reg_10_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_2_VALID_5_6_0_inputs_ready;
 reg SFC_2_VALID_5_6_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_5_6_0_stall_in;
wire SFC_2_VALID_5_6_0_output_regs_ready;
 reg SFC_2_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_5_6_0_causedstall;

assign SFC_2_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_stall_in = 1'b0;
assign SFC_2_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_5_6_0_output_regs_ready)
		begin
			SFC_2_VALID_5_6_0_NO_SHIFT_REG <= SFC_2_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_6_7_0_inputs_ready;
 reg SFC_2_VALID_6_7_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_6_7_0_stall_in_0;
 reg SFC_2_VALID_6_7_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_6_7_0_stall_in_1;
wire SFC_2_VALID_6_7_0_output_regs_ready;
 reg SFC_2_VALID_6_7_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_6_7_0_causedstall;

assign SFC_2_VALID_6_7_0_inputs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_stall_in = 1'b0;
assign SFC_2_VALID_6_7_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_6_7_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_6_7_0_output_regs_ready)
		begin
			SFC_2_VALID_6_7_0_NO_SHIFT_REG <= SFC_2_VALID_5_6_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_7_8_0_inputs_ready;
 reg SFC_2_VALID_7_8_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_7_8_0_stall_in;
wire SFC_2_VALID_7_8_0_output_regs_ready;
 reg SFC_2_VALID_7_8_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_7_8_0_causedstall;

assign SFC_2_VALID_7_8_0_inputs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_7_8_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_7_8_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_7_8_0_output_regs_ready)
		begin
			SFC_2_VALID_7_8_0_NO_SHIFT_REG <= SFC_2_VALID_6_7_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_indvars_iv_pop7__stall_local;
wire [63:0] local_bb4_indvars_iv_pop7_;
wire local_bb4_indvars_iv_pop7__fu_valid_out;
wire local_bb4_indvars_iv_pop7__fu_stall_out;

acl_pop local_bb4_indvars_iv_pop7__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_6to7_bb4_c0_ene1209_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(input_wii_var_),
	.stall_out(local_bb4_indvars_iv_pop7__fu_stall_out),
	.valid_in(SFC_2_VALID_6_7_0_NO_SHIFT_REG),
	.valid_out(local_bb4_indvars_iv_pop7__fu_valid_out),
	.stall_in(local_bb4_indvars_iv_pop7__stall_local),
	.data_out(local_bb4_indvars_iv_pop7_),
	.feedback_in(feedback_data_in_7),
	.feedback_valid_in(feedback_valid_in_7),
	.feedback_stall_out(feedback_stall_out_7)
);

defparam local_bb4_indvars_iv_pop7__feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_indvars_iv_pop7__feedback.DATA_WIDTH = 64;
defparam local_bb4_indvars_iv_pop7__feedback.STYLE = "REGULAR";

assign local_bb4_indvars_iv_pop7__stall_local = 1'b0;

// This section implements a registered operation.
// 
wire SFC_2_VALID_8_9_0_inputs_ready;
 reg SFC_2_VALID_8_9_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_0;
 reg SFC_2_VALID_8_9_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_1;
 reg SFC_2_VALID_8_9_0_valid_out_2_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_2;
 reg SFC_2_VALID_8_9_0_valid_out_3_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_3;
 reg SFC_2_VALID_8_9_0_valid_out_4_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_4;
wire SFC_2_VALID_8_9_0_output_regs_ready;
 reg SFC_2_VALID_8_9_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_8_9_0_causedstall;

assign SFC_2_VALID_8_9_0_inputs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_stall_in = 1'b0;
assign SFC_2_VALID_8_9_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_8_9_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_8_9_0_output_regs_ready)
		begin
			SFC_2_VALID_8_9_0_NO_SHIFT_REG <= SFC_2_VALID_7_8_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__stall_local;
wire [31:0] local_bb4_var_;

assign local_bb4_var_ = local_bb4_indvars_iv_pop7_[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u23_stall_local;
wire [63:0] local_bb4_var__u23;

assign local_bb4_var__u23 = (local_bb4_indvars_iv_pop7_ + input_wii_var__u19);

// This section implements an unregistered operation.
// 
wire local_bb4_indvars_iv_next_stall_local;
wire [63:0] local_bb4_indvars_iv_next;

assign local_bb4_indvars_iv_next = (local_bb4_indvars_iv_pop7_ + 64'h1);

// This section implements a registered operation.
// 
wire SFC_2_VALID_9_10_0_inputs_ready;
 reg SFC_2_VALID_9_10_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_0;
 reg SFC_2_VALID_9_10_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_1;
 reg SFC_2_VALID_9_10_0_valid_out_2_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_2;
 reg SFC_2_VALID_9_10_0_valid_out_3_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_3;
 reg SFC_2_VALID_9_10_0_valid_out_4_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_4;
 reg SFC_2_VALID_9_10_0_valid_out_5_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_5;
 reg SFC_2_VALID_9_10_0_valid_out_6_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_6;
 reg SFC_2_VALID_9_10_0_valid_out_7_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_7;
wire SFC_2_VALID_9_10_0_output_regs_ready;
 reg SFC_2_VALID_9_10_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_9_10_0_causedstall;

assign SFC_2_VALID_9_10_0_inputs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_9_10_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_9_10_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_9_10_0_output_regs_ready)
		begin
			SFC_2_VALID_9_10_0_NO_SHIFT_REG <= SFC_2_VALID_8_9_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_keep_going_acl_pipeline_1_inputs_ready;
 reg local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb4_keep_going_acl_pipeline_1_stall_in;
wire local_bb4_keep_going_acl_pipeline_1_output_regs_ready;
wire local_bb4_keep_going_acl_pipeline_1_keep_going;
wire local_bb4_keep_going_acl_pipeline_1_fu_valid_out;
wire local_bb4_keep_going_acl_pipeline_1_fu_stall_out;
 reg local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb4_keep_going_acl_pipeline_1_feedback_pipelined;
wire local_bb4_keep_going_acl_pipeline_1_causedstall;

acl_pipeline local_bb4_keep_going_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb4_keep_going_acl_pipeline_1_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_keep_going_acl_pipeline_1_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_keep_going_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_0),
	.not_exitcond_in(feedback_data_in_1),
	.not_exitcond_valid_in(feedback_valid_in_1),
	.not_exitcond_stall_out(feedback_stall_out_1),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb4_keep_going_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb4_keep_going_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb4_keep_going_acl_pipeline_1_inputs_ready = 1'b1;
assign local_bb4_keep_going_acl_pipeline_1_output_regs_ready = 1'b1;
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign SFC_2_VALID_8_9_0_stall_in_1 = 1'b0;
assign rnode_7to9_bb4_c0_ene1209_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb4_keep_going_acl_pipeline_1_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_keep_going_acl_pipeline_1_output_regs_ready)
		begin
			local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG <= local_bb4_keep_going_acl_pipeline_1_keep_going;
			local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_keep_going_acl_pipeline_1_stall_in))
			begin
				local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_sub17_add16204_pop10_c0_ene2_stall_local;
wire [31:0] local_bb4_sub17_add16204_pop10_c0_ene2;
wire local_bb4_sub17_add16204_pop10_c0_ene2_fu_valid_out;
wire local_bb4_sub17_add16204_pop10_c0_ene2_fu_stall_out;

acl_pop local_bb4_sub17_add16204_pop10_c0_ene2_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_7to9_bb4_c0_ene1209_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_8to9_bb4_c0_ene2_0_NO_SHIFT_REG),
	.stall_out(local_bb4_sub17_add16204_pop10_c0_ene2_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sub17_add16204_pop10_c0_ene2_fu_valid_out),
	.stall_in(local_bb4_sub17_add16204_pop10_c0_ene2_stall_local),
	.data_out(local_bb4_sub17_add16204_pop10_c0_ene2),
	.feedback_in(feedback_data_in_10),
	.feedback_valid_in(feedback_valid_in_10),
	.feedback_stall_out(feedback_stall_out_10)
);

defparam local_bb4_sub17_add16204_pop10_c0_ene2_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_sub17_add16204_pop10_c0_ene2_feedback.DATA_WIDTH = 32;
defparam local_bb4_sub17_add16204_pop10_c0_ene2_feedback.STYLE = "REGULAR";

assign local_bb4_sub17_add16204_pop10_c0_ene2_stall_local = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_add18_stall_local;
wire [31:0] local_bb4_add18;

assign local_bb4_add18 = (local_bb4_var_ + local_bb4__acl_ffwd_dest_i32_1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u23_valid_out;
wire local_bb4_var__u23_stall_in;
wire local_bb4_indvars_iv_next_valid_out_1;
wire local_bb4_indvars_iv_next_stall_in_1;
wire local_bb4_add18_valid_out;
wire local_bb4_add18_stall_in;
wire local_bb4_var__u24_valid_out;
wire local_bb4_var__u24_stall_in;
wire local_bb4_var__u24_inputs_ready;
wire local_bb4_var__u24_stall_local;
wire [31:0] local_bb4_var__u24;

assign local_bb4_var__u24_inputs_ready = (SFC_2_VALID_6_7_0_valid_out_1_NO_SHIFT_REG & rnode_6to7_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG & rnode_6to7_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_var__u24 = local_bb4_indvars_iv_next[31:0];
assign local_bb4_var__u23_valid_out = 1'b1;
assign local_bb4_indvars_iv_next_valid_out_1 = 1'b1;
assign local_bb4_add18_valid_out = 1'b1;
assign local_bb4_var__u24_valid_out = 1'b1;
assign SFC_2_VALID_6_7_0_stall_in_1 = 1'b0;
assign rnode_6to7_bb4_c0_ene1209_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene1209_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_2_VALID_10_11_0_inputs_ready;
 reg SFC_2_VALID_10_11_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_10_11_0_stall_in;
wire SFC_2_VALID_10_11_0_output_regs_ready;
 reg SFC_2_VALID_10_11_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_10_11_0_causedstall;

assign SFC_2_VALID_10_11_0_inputs_ready = 1'b1;
assign SFC_2_VALID_10_11_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_10_11_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_10_11_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_10_11_0_output_regs_ready)
		begin
			SFC_2_VALID_10_11_0_NO_SHIFT_REG <= SFC_2_VALID_9_10_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_arrayidx32205_pop11_c0_ene3_valid_out_0;
wire local_bb4_arrayidx32205_pop11_c0_ene3_stall_in_0;
wire local_bb4_arrayidx32205_pop11_c0_ene3_valid_out_1;
wire local_bb4_arrayidx32205_pop11_c0_ene3_stall_in_1;
wire local_bb4_arrayidx32205_pop11_c0_ene3_inputs_ready;
wire local_bb4_arrayidx32205_pop11_c0_ene3_stall_local;
wire [63:0] local_bb4_arrayidx32205_pop11_c0_ene3;
wire local_bb4_arrayidx32205_pop11_c0_ene3_fu_valid_out;
wire local_bb4_arrayidx32205_pop11_c0_ene3_fu_stall_out;

acl_pop local_bb4_arrayidx32205_pop11_c0_ene3_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene1209_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene3_0_NO_SHIFT_REG),
	.stall_out(local_bb4_arrayidx32205_pop11_c0_ene3_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_arrayidx32205_pop11_c0_ene3_fu_valid_out),
	.stall_in(local_bb4_arrayidx32205_pop11_c0_ene3_stall_local),
	.data_out(local_bb4_arrayidx32205_pop11_c0_ene3),
	.feedback_in(feedback_data_in_11),
	.feedback_valid_in(feedback_valid_in_11),
	.feedback_stall_out(feedback_stall_out_11)
);

defparam local_bb4_arrayidx32205_pop11_c0_ene3_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_arrayidx32205_pop11_c0_ene3_feedback.DATA_WIDTH = 64;
defparam local_bb4_arrayidx32205_pop11_c0_ene3_feedback.STYLE = "REGULAR";

assign local_bb4_arrayidx32205_pop11_c0_ene3_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_1_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene1209_0_valid_out_0_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG);
assign local_bb4_arrayidx32205_pop11_c0_ene3_stall_local = 1'b0;
assign local_bb4_arrayidx32205_pop11_c0_ene3_valid_out_0 = 1'b1;
assign local_bb4_arrayidx32205_pop11_c0_ene3_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_1 = 1'b0;
assign rnode_9to10_bb4_c0_ene1209_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__pop12_c0_ene4_valid_out_0;
wire local_bb4__pop12_c0_ene4_stall_in_0;
wire local_bb4__pop12_c0_ene4_valid_out_1;
wire local_bb4__pop12_c0_ene4_stall_in_1;
wire local_bb4__pop12_c0_ene4_inputs_ready;
wire local_bb4__pop12_c0_ene4_stall_local;
wire local_bb4__pop12_c0_ene4;
wire local_bb4__pop12_c0_ene4_fu_valid_out;
wire local_bb4__pop12_c0_ene4_fu_stall_out;

acl_pop local_bb4__pop12_c0_ene4_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene1209_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene4_0_NO_SHIFT_REG),
	.stall_out(local_bb4__pop12_c0_ene4_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__pop12_c0_ene4_fu_valid_out),
	.stall_in(local_bb4__pop12_c0_ene4_stall_local),
	.data_out(local_bb4__pop12_c0_ene4),
	.feedback_in(feedback_data_in_12),
	.feedback_valid_in(feedback_valid_in_12),
	.feedback_stall_out(feedback_stall_out_12)
);

defparam local_bb4__pop12_c0_ene4_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4__pop12_c0_ene4_feedback.DATA_WIDTH = 1;
defparam local_bb4__pop12_c0_ene4_feedback.STYLE = "REGULAR";

assign local_bb4__pop12_c0_ene4_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_2_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG);
assign local_bb4__pop12_c0_ene4_stall_local = 1'b0;
assign local_bb4__pop12_c0_ene4_valid_out_0 = 1'b1;
assign local_bb4__pop12_c0_ene4_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_2 = 1'b0;
assign rnode_9to10_bb4_c0_ene1209_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notexitcond201206_pop13_c0_ene5_valid_out_0;
wire local_bb4_notexitcond201206_pop13_c0_ene5_stall_in_0;
wire local_bb4_notexitcond201206_pop13_c0_ene5_valid_out_1;
wire local_bb4_notexitcond201206_pop13_c0_ene5_stall_in_1;
wire local_bb4_notexitcond201206_pop13_c0_ene5_inputs_ready;
wire local_bb4_notexitcond201206_pop13_c0_ene5_stall_local;
wire local_bb4_notexitcond201206_pop13_c0_ene5;
wire local_bb4_notexitcond201206_pop13_c0_ene5_fu_valid_out;
wire local_bb4_notexitcond201206_pop13_c0_ene5_fu_stall_out;

acl_pop local_bb4_notexitcond201206_pop13_c0_ene5_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene1209_2_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene5_0_NO_SHIFT_REG),
	.stall_out(local_bb4_notexitcond201206_pop13_c0_ene5_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond201206_pop13_c0_ene5_fu_valid_out),
	.stall_in(local_bb4_notexitcond201206_pop13_c0_ene5_stall_local),
	.data_out(local_bb4_notexitcond201206_pop13_c0_ene5),
	.feedback_in(feedback_data_in_13),
	.feedback_valid_in(feedback_valid_in_13),
	.feedback_stall_out(feedback_stall_out_13)
);

defparam local_bb4_notexitcond201206_pop13_c0_ene5_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_notexitcond201206_pop13_c0_ene5_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond201206_pop13_c0_ene5_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond201206_pop13_c0_ene5_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_3_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notexitcond201206_pop13_c0_ene5_stall_local = 1'b0;
assign local_bb4_notexitcond201206_pop13_c0_ene5_valid_out_0 = 1'b1;
assign local_bb4_notexitcond201206_pop13_c0_ene5_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_3 = 1'b0;
assign rnode_9to10_bb4_c0_ene1209_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_keep_going_acl_pipeline_1_stall_in = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_NO_SHIFT_REG = rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_var__u23_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u23_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_7to8_bb4_var__u23_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u23_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_7to8_bb4_var__u23_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u23_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u23_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u23_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_var__u23_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_var__u23_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_var__u23_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_var__u23_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_var__u23_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_bb4_var__u23),
	.data_out(rnode_7to8_bb4_var__u23_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_var__u23_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_var__u23_0_reg_8_fifo.DATA_WIDTH = 64;
defparam rnode_7to8_bb4_var__u23_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_var__u23_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_var__u23_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u23_stall_in = 1'b0;
assign rnode_7to8_bb4_var__u23_0_NO_SHIFT_REG = rnode_7to8_bb4_var__u23_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_var__u23_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_var__u23_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_7to9_bb4_indvars_iv_next_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to9_bb4_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_7to9_bb4_indvars_iv_next_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_indvars_iv_next_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_7to9_bb4_indvars_iv_next_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_indvars_iv_next_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_indvars_iv_next_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_indvars_iv_next_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_7to9_bb4_indvars_iv_next_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to9_bb4_indvars_iv_next_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to9_bb4_indvars_iv_next_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_7to9_bb4_indvars_iv_next_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_7to9_bb4_indvars_iv_next_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(local_bb4_indvars_iv_next),
	.data_out(rnode_7to9_bb4_indvars_iv_next_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_7to9_bb4_indvars_iv_next_0_reg_9_fifo.DEPTH = 2;
defparam rnode_7to9_bb4_indvars_iv_next_0_reg_9_fifo.DATA_WIDTH = 64;
defparam rnode_7to9_bb4_indvars_iv_next_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to9_bb4_indvars_iv_next_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_7to9_bb4_indvars_iv_next_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_indvars_iv_next_stall_in_1 = 1'b0;
assign rnode_7to9_bb4_indvars_iv_next_0_NO_SHIFT_REG = rnode_7to9_bb4_indvars_iv_next_0_reg_9_NO_SHIFT_REG;
assign rnode_7to9_bb4_indvars_iv_next_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_7to9_bb4_indvars_iv_next_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_add18_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add18_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add18_1_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add18_2_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add18_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_valid_out_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_stall_in_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add18_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_add18_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_add18_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_add18_0_stall_in_0_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_add18_0_valid_out_0_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_add18_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_bb4_add18),
	.data_out(rnode_7to8_bb4_add18_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_add18_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_add18_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_7to8_bb4_add18_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_add18_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_add18_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add18_stall_in = 1'b0;
assign rnode_7to8_bb4_add18_0_stall_in_0_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_add18_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add18_0_NO_SHIFT_REG = rnode_7to8_bb4_add18_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_add18_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add18_1_NO_SHIFT_REG = rnode_7to8_bb4_add18_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_add18_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add18_2_NO_SHIFT_REG = rnode_7to8_bb4_add18_0_reg_8_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_var__u24_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u24_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_var__u24_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u24_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_var__u24_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u24_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u24_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u24_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_var__u24_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_var__u24_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_var__u24_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_var__u24_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_var__u24_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_bb4_var__u24),
	.data_out(rnode_7to8_bb4_var__u24_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_var__u24_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_var__u24_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_7to8_bb4_var__u24_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_var__u24_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_var__u24_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u24_stall_in = 1'b0;
assign rnode_7to8_bb4_var__u24_0_NO_SHIFT_REG = rnode_7to8_bb4_var__u24_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_var__u24_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_var__u24_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_arrayidx32205_pop11_c0_ene3),
	.data_out(rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_arrayidx32205_pop11_c0_ene3_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_NO_SHIFT_REG = rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4__pop12_c0_ene4_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4__pop12_c0_ene4),
	.data_out(rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__pop12_c0_ene4_stall_in_1 = 1'b0;
assign rnode_10to11_bb4__pop12_c0_ene4_0_NO_SHIFT_REG = rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond201206_pop13_c0_ene5),
	.data_out(rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond201206_pop13_c0_ene5_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_NO_SHIFT_REG = rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_arrayidx35_valid_out;
wire local_bb4_arrayidx35_stall_in;
wire local_bb4_arrayidx35_inputs_ready;
wire local_bb4_arrayidx35_stall_local;
wire [63:0] local_bb4_arrayidx35;

assign local_bb4_arrayidx35_inputs_ready = rnode_7to8_bb4_var__u23_0_valid_out_NO_SHIFT_REG;
assign local_bb4_arrayidx35 = ((input_gaussian & 64'hFFFFFFFFFFFFFC00) + (rnode_7to8_bb4_var__u23_0_NO_SHIFT_REG << 6'h2));
assign local_bb4_arrayidx35_valid_out = 1'b1;
assign rnode_7to8_bb4_var__u23_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp1_i3_stall_local;
wire local_bb4_cmp1_i3;

assign local_bb4_cmp1_i3 = (rnode_7to8_bb4_add18_0_NO_SHIFT_REG > 32'hEF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u25_stall_local;
wire [31:0] local_bb4_var__u25;

assign local_bb4_var__u25 = (rnode_7to8_bb4_add18_1_NO_SHIFT_REG << 32'h6);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u26_stall_local;
wire [31:0] local_bb4_var__u26;

assign local_bb4_var__u26 = (rnode_7to8_bb4_add18_2_NO_SHIFT_REG << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp14_valid_out;
wire local_bb4_cmp14_stall_in;
wire local_bb4_cmp14_inputs_ready;
wire local_bb4_cmp14_stall_local;
wire local_bb4_cmp14;

assign local_bb4_cmp14_inputs_ready = rnode_7to8_bb4_var__u24_0_valid_out_NO_SHIFT_REG;
assign local_bb4_cmp14 = ($signed(rnode_7to8_bb4_var__u24_0_NO_SHIFT_REG) > $signed(input_r));
assign local_bb4_cmp14_valid_out = 1'b1;
assign rnode_7to8_bb4_var__u24_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_arrayidx35_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_arrayidx35_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_8to9_bb4_arrayidx35_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_arrayidx35_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_8to9_bb4_arrayidx35_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_arrayidx35_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_arrayidx35_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_arrayidx35_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_arrayidx35_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_arrayidx35_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_arrayidx35_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_arrayidx35_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_arrayidx35_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in((local_bb4_arrayidx35 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_8to9_bb4_arrayidx35_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_arrayidx35_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_arrayidx35_0_reg_9_fifo.DATA_WIDTH = 64;
defparam rnode_8to9_bb4_arrayidx35_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_arrayidx35_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_arrayidx35_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_arrayidx35_stall_in = 1'b0;
assign rnode_8to9_bb4_arrayidx35_0_NO_SHIFT_REG = rnode_8to9_bb4_arrayidx35_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_arrayidx35_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_arrayidx35_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_add18_op_add188_stall_local;
wire [31:0] local_bb4_add18_op_add188;

assign local_bb4_add18_op_add188 = ((local_bb4_var__u25 & 32'hFFFFFFC0) + (local_bb4_var__u26 & 32'hFFFFFF00));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_cmp14_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_cmp14_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_cmp14_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_cmp14_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_cmp14_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_cmp14_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(local_bb4_cmp14),
	.data_out(rnode_8to9_bb4_cmp14_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_cmp14_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp14_stall_in = 1'b0;
assign rnode_8to9_bb4_cmp14_0_NO_SHIFT_REG = rnode_8to9_bb4_cmp14_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_cmp14_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_cmp14_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_arrayidx35_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_arrayidx35_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_9to10_bb4_arrayidx35_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_arrayidx35_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_9to10_bb4_arrayidx35_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_arrayidx35_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_arrayidx35_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_arrayidx35_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_arrayidx35_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_arrayidx35_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_arrayidx35_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_arrayidx35_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_arrayidx35_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in((rnode_8to9_bb4_arrayidx35_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_9to10_bb4_arrayidx35_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_arrayidx35_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_arrayidx35_0_reg_10_fifo.DATA_WIDTH = 64;
defparam rnode_9to10_bb4_arrayidx35_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_arrayidx35_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_arrayidx35_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_arrayidx35_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_arrayidx35_0_NO_SHIFT_REG = rnode_9to10_bb4_arrayidx35_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_arrayidx35_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_arrayidx35_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_phitmp_valid_out;
wire local_bb4_phitmp_stall_in;
wire local_bb4_phitmp_inputs_ready;
wire local_bb4_phitmp_stall_local;
wire [31:0] local_bb4_phitmp;

assign local_bb4_phitmp_inputs_ready = (rnode_7to8_bb4_add18_0_valid_out_0_NO_SHIFT_REG & rnode_7to8_bb4_add18_0_valid_out_1_NO_SHIFT_REG & rnode_7to8_bb4_add18_0_valid_out_2_NO_SHIFT_REG);
assign local_bb4_phitmp = (local_bb4_cmp1_i3 ? 32'h12AC0 : (local_bb4_add18_op_add188 & 32'hFFFFFFC0));
assign local_bb4_phitmp_valid_out = 1'b1;
assign rnode_7to8_bb4_add18_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_add18_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_add18_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u27_stall_local;
wire local_bb4_var__u27;

assign local_bb4_var__u27 = (local_bb4__acl_ffwd_dest_i1_10_u22 | rnode_8to9_bb4_cmp14_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_arrayidx35_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx35_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx35_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx35_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx35_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx35_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx35_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx35_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_arrayidx35_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_arrayidx35_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_arrayidx35_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_arrayidx35_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_arrayidx35_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in((rnode_9to10_bb4_arrayidx35_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_10to11_bb4_arrayidx35_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_arrayidx35_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_arrayidx35_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_arrayidx35_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_arrayidx35_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_arrayidx35_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_arrayidx35_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx35_0_NO_SHIFT_REG = rnode_10to11_bb4_arrayidx35_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_arrayidx35_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx35_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_phitmp_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_phitmp_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_phitmp_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_phitmp_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_phitmp_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_phitmp_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_phitmp_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_phitmp_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_phitmp_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_phitmp_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_phitmp_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_phitmp_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_phitmp_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in((local_bb4_phitmp & 32'hFFFFFFC0)),
	.data_out(rnode_8to9_bb4_phitmp_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_phitmp_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_phitmp_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4_phitmp_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_phitmp_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_phitmp_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_phitmp_stall_in = 1'b0;
assign rnode_8to9_bb4_phitmp_0_NO_SHIFT_REG = rnode_8to9_bb4_phitmp_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_phitmp_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_phitmp_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u27_valid_out_1;
wire local_bb4_var__u27_stall_in_1;
wire local_bb4_notexit_valid_out_0;
wire local_bb4_notexit_stall_in_0;
wire local_bb4_notexit_valid_out_1;
wire local_bb4_notexit_stall_in_1;
wire local_bb4_notexit_inputs_ready;
wire local_bb4_notexit_stall_local;
wire local_bb4_notexit;

assign local_bb4_notexit_inputs_ready = (rnode_7to9_bb4_c0_ene1209_0_valid_out_2_NO_SHIFT_REG & rnode_8to9_bb4_cmp14_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notexit = (local_bb4_var__u27 ^ 1'b1);
assign local_bb4_var__u27_valid_out_1 = 1'b1;
assign local_bb4_notexit_valid_out_0 = 1'b1;
assign local_bb4_notexit_valid_out_1 = 1'b1;
assign rnode_7to9_bb4_c0_ene1209_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_cmp14_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_sub17_add16204_pop10_c0_ene2_valid_out_1;
wire local_bb4_sub17_add16204_pop10_c0_ene2_stall_in_1;
wire local_bb4_add23_valid_out;
wire local_bb4_add23_stall_in;
wire local_bb4_add23_inputs_ready;
wire local_bb4_add23_stall_local;
wire [31:0] local_bb4_add23;

assign local_bb4_add23_inputs_ready = (SFC_2_VALID_8_9_0_valid_out_2_NO_SHIFT_REG & rnode_7to9_bb4_c0_ene1209_0_valid_out_1_NO_SHIFT_REG & rnode_8to9_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG & rnode_8to9_bb4_phitmp_0_valid_out_NO_SHIFT_REG);
assign local_bb4_add23 = ((rnode_8to9_bb4_phitmp_0_NO_SHIFT_REG & 32'hFFFFFFC0) + local_bb4_sub17_add16204_pop10_c0_ene2);
assign local_bb4_sub17_add16204_pop10_c0_ene2_valid_out_1 = 1'b1;
assign local_bb4_add23_valid_out = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in_2 = 1'b0;
assign rnode_7to9_bb4_c0_ene1209_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_phitmp_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_9to11_bb4_var__u27_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__u27_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__u27_0_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__u27_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__u27_0_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__u27_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__u27_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__u27_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_9to11_bb4_var__u27_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to11_bb4_var__u27_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to11_bb4_var__u27_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_9to11_bb4_var__u27_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_9to11_bb4_var__u27_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_var__u27),
	.data_out(rnode_9to11_bb4_var__u27_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_9to11_bb4_var__u27_0_reg_11_fifo.DEPTH = 2;
defparam rnode_9to11_bb4_var__u27_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_9to11_bb4_var__u27_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to11_bb4_var__u27_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_9to11_bb4_var__u27_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u27_stall_in_1 = 1'b0;
assign rnode_9to11_bb4_var__u27_0_NO_SHIFT_REG = rnode_9to11_bb4_var__u27_0_reg_11_NO_SHIFT_REG;
assign rnode_9to11_bb4_var__u27_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_var__u27_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_notexitcond_notexit_inputs_ready;
 reg local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_0;
 reg local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_1;
 reg local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_2;
 reg local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_3;
 reg local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_4;
wire local_bb4_notexitcond_notexit_output_regs_ready;
wire local_bb4_notexitcond_notexit_result;
wire local_bb4_notexitcond_notexit_fu_valid_out;
wire local_bb4_notexitcond_notexit_fu_stall_out;
 reg local_bb4_notexitcond_notexit_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_causedstall;

acl_push local_bb4_notexitcond_notexit_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(local_bb4_notexit),
	.stall_out(local_bb4_notexitcond_notexit_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond_notexit_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond_notexit_result),
	.feedback_out(feedback_data_out_1),
	.feedback_valid_out(feedback_valid_out_1),
	.feedback_stall_in(feedback_stall_in_1)
);

defparam local_bb4_notexitcond_notexit_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond_notexit_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond_notexit_feedback.FIFO_DEPTH = 8;
defparam local_bb4_notexitcond_notexit_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_notexitcond_notexit_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond_notexit_inputs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_output_regs_ready = 1'b1;
assign local_bb4_notexit_stall_in_0 = 1'b0;
assign SFC_2_VALID_8_9_0_stall_in_3 = 1'b0;
assign local_bb4_notexitcond_notexit_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond_notexit_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond_notexit_output_regs_ready)
		begin
			local_bb4_notexitcond_notexit_NO_SHIFT_REG <= local_bb4_notexitcond_notexit_result;
			local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond_notexit_stall_in_0))
			begin
				local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_1))
			begin
				local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_2))
			begin
				local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_3))
			begin
				local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_4))
			begin
				local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_indvars_iv_push7_indvars_iv_next_inputs_ready;
 reg local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG;
wire local_bb4_indvars_iv_push7_indvars_iv_next_stall_in;
wire local_bb4_indvars_iv_push7_indvars_iv_next_output_regs_ready;
wire [63:0] local_bb4_indvars_iv_push7_indvars_iv_next_result;
wire local_bb4_indvars_iv_push7_indvars_iv_next_fu_valid_out;
wire local_bb4_indvars_iv_push7_indvars_iv_next_fu_stall_out;
 reg [63:0] local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG;
wire local_bb4_indvars_iv_push7_indvars_iv_next_causedstall;

acl_push local_bb4_indvars_iv_push7_indvars_iv_next_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexit),
	.predicate(1'b0),
	.data_in(rnode_7to9_bb4_indvars_iv_next_0_NO_SHIFT_REG),
	.stall_out(local_bb4_indvars_iv_push7_indvars_iv_next_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_indvars_iv_push7_indvars_iv_next_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_indvars_iv_push7_indvars_iv_next_result),
	.feedback_out(feedback_data_out_7),
	.feedback_valid_out(feedback_valid_out_7),
	.feedback_stall_in(feedback_stall_in_7)
);

defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.STALLFREE = 1;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.DATA_WIDTH = 64;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.FIFO_DEPTH = 9;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.MIN_FIFO_LATENCY = 7;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.STYLE = "REGULAR";

assign local_bb4_indvars_iv_push7_indvars_iv_next_inputs_ready = 1'b1;
assign local_bb4_indvars_iv_push7_indvars_iv_next_output_regs_ready = 1'b1;
assign local_bb4_notexit_stall_in_1 = 1'b0;
assign SFC_2_VALID_8_9_0_stall_in_4 = 1'b0;
assign rnode_7to9_bb4_indvars_iv_next_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_indvars_iv_push7_indvars_iv_next_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG <= 'x;
		local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_indvars_iv_push7_indvars_iv_next_output_regs_ready)
		begin
			local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG <= local_bb4_indvars_iv_push7_indvars_iv_next_result;
			local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_indvars_iv_push7_indvars_iv_next_stall_in))
			begin
				local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(local_bb4_sub17_add16204_pop10_c0_ene2),
	.data_out(rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_sub17_add16204_pop10_c0_ene2_stall_in_1 = 1'b0;
assign rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_NO_SHIFT_REG = rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_add23_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add23_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_add23_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add23_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_add23_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add23_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add23_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add23_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_add23_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_add23_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_add23_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_add23_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_add23_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(local_bb4_add23),
	.data_out(rnode_9to10_bb4_add23_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_add23_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_add23_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_add23_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_add23_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_add23_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add23_stall_in = 1'b0;
assign rnode_9to10_bb4_add23_0_NO_SHIFT_REG = rnode_9to10_bb4_add23_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_add23_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_add23_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_arrayidx32205_push11_arrayidx32205_pop11_inputs_ready;
 reg local_bb4_arrayidx32205_push11_arrayidx32205_pop11_valid_out_NO_SHIFT_REG;
wire local_bb4_arrayidx32205_push11_arrayidx32205_pop11_stall_in;
wire local_bb4_arrayidx32205_push11_arrayidx32205_pop11_output_regs_ready;
wire [63:0] local_bb4_arrayidx32205_push11_arrayidx32205_pop11_result;
wire local_bb4_arrayidx32205_push11_arrayidx32205_pop11_fu_valid_out;
wire local_bb4_arrayidx32205_push11_arrayidx32205_pop11_fu_stall_out;
 reg [63:0] local_bb4_arrayidx32205_push11_arrayidx32205_pop11_NO_SHIFT_REG;
wire local_bb4_arrayidx32205_push11_arrayidx32205_pop11_causedstall;

acl_push local_bb4_arrayidx32205_push11_arrayidx32205_pop11_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_arrayidx32205_pop11_c0_ene3),
	.stall_out(local_bb4_arrayidx32205_push11_arrayidx32205_pop11_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_arrayidx32205_push11_arrayidx32205_pop11_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_arrayidx32205_push11_arrayidx32205_pop11_result),
	.feedback_out(feedback_data_out_11),
	.feedback_valid_out(feedback_valid_out_11),
	.feedback_stall_in(feedback_stall_in_11)
);

defparam local_bb4_arrayidx32205_push11_arrayidx32205_pop11_feedback.STALLFREE = 1;
defparam local_bb4_arrayidx32205_push11_arrayidx32205_pop11_feedback.DATA_WIDTH = 64;
defparam local_bb4_arrayidx32205_push11_arrayidx32205_pop11_feedback.FIFO_DEPTH = 9;
defparam local_bb4_arrayidx32205_push11_arrayidx32205_pop11_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_arrayidx32205_push11_arrayidx32205_pop11_feedback.STYLE = "REGULAR";

assign local_bb4_arrayidx32205_push11_arrayidx32205_pop11_inputs_ready = 1'b1;
assign local_bb4_arrayidx32205_push11_arrayidx32205_pop11_output_regs_ready = 1'b1;
assign local_bb4_arrayidx32205_pop11_c0_ene3_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_0 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_4 = 1'b0;
assign local_bb4_arrayidx32205_push11_arrayidx32205_pop11_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_arrayidx32205_push11_arrayidx32205_pop11_NO_SHIFT_REG <= 'x;
		local_bb4_arrayidx32205_push11_arrayidx32205_pop11_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_arrayidx32205_push11_arrayidx32205_pop11_output_regs_ready)
		begin
			local_bb4_arrayidx32205_push11_arrayidx32205_pop11_NO_SHIFT_REG <= local_bb4_arrayidx32205_push11_arrayidx32205_pop11_result;
			local_bb4_arrayidx32205_push11_arrayidx32205_pop11_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_arrayidx32205_push11_arrayidx32205_pop11_stall_in))
			begin
				local_bb4_arrayidx32205_push11_arrayidx32205_pop11_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4__push12__pop12_inputs_ready;
 reg local_bb4__push12__pop12_valid_out_NO_SHIFT_REG;
wire local_bb4__push12__pop12_stall_in;
wire local_bb4__push12__pop12_output_regs_ready;
wire local_bb4__push12__pop12_result;
wire local_bb4__push12__pop12_fu_valid_out;
wire local_bb4__push12__pop12_fu_stall_out;
 reg local_bb4__push12__pop12_NO_SHIFT_REG;
wire local_bb4__push12__pop12_causedstall;

acl_push local_bb4__push12__pop12_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4__pop12_c0_ene4),
	.stall_out(local_bb4__push12__pop12_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__push12__pop12_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4__push12__pop12_result),
	.feedback_out(feedback_data_out_12),
	.feedback_valid_out(feedback_valid_out_12),
	.feedback_stall_in(feedback_stall_in_12)
);

defparam local_bb4__push12__pop12_feedback.STALLFREE = 1;
defparam local_bb4__push12__pop12_feedback.DATA_WIDTH = 1;
defparam local_bb4__push12__pop12_feedback.FIFO_DEPTH = 9;
defparam local_bb4__push12__pop12_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4__push12__pop12_feedback.STYLE = "REGULAR";

assign local_bb4__push12__pop12_inputs_ready = 1'b1;
assign local_bb4__push12__pop12_output_regs_ready = 1'b1;
assign local_bb4__pop12_c0_ene4_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_2 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_6 = 1'b0;
assign local_bb4__push12__pop12_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4__push12__pop12_NO_SHIFT_REG <= 'x;
		local_bb4__push12__pop12_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4__push12__pop12_output_regs_ready)
		begin
			local_bb4__push12__pop12_NO_SHIFT_REG <= local_bb4__push12__pop12_result;
			local_bb4__push12__pop12_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4__push12__pop12_stall_in))
			begin
				local_bb4__push12__pop12_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_notexitcond201206_push13_notexitcond201206_pop13_inputs_ready;
 reg local_bb4_notexitcond201206_push13_notexitcond201206_pop13_valid_out_NO_SHIFT_REG;
wire local_bb4_notexitcond201206_push13_notexitcond201206_pop13_stall_in;
wire local_bb4_notexitcond201206_push13_notexitcond201206_pop13_output_regs_ready;
wire local_bb4_notexitcond201206_push13_notexitcond201206_pop13_result;
wire local_bb4_notexitcond201206_push13_notexitcond201206_pop13_fu_valid_out;
wire local_bb4_notexitcond201206_push13_notexitcond201206_pop13_fu_stall_out;
 reg local_bb4_notexitcond201206_push13_notexitcond201206_pop13_NO_SHIFT_REG;
wire local_bb4_notexitcond201206_push13_notexitcond201206_pop13_causedstall;

acl_push local_bb4_notexitcond201206_push13_notexitcond201206_pop13_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_notexitcond201206_pop13_c0_ene5),
	.stall_out(local_bb4_notexitcond201206_push13_notexitcond201206_pop13_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond201206_push13_notexitcond201206_pop13_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond201206_push13_notexitcond201206_pop13_result),
	.feedback_out(feedback_data_out_13),
	.feedback_valid_out(feedback_valid_out_13),
	.feedback_stall_in(feedback_stall_in_13)
);

defparam local_bb4_notexitcond201206_push13_notexitcond201206_pop13_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond201206_push13_notexitcond201206_pop13_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond201206_push13_notexitcond201206_pop13_feedback.FIFO_DEPTH = 9;
defparam local_bb4_notexitcond201206_push13_notexitcond201206_pop13_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_notexitcond201206_push13_notexitcond201206_pop13_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond201206_push13_notexitcond201206_pop13_inputs_ready = 1'b1;
assign local_bb4_notexitcond201206_push13_notexitcond201206_pop13_output_regs_ready = 1'b1;
assign local_bb4_notexitcond201206_pop13_c0_ene5_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_3 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_7 = 1'b0;
assign local_bb4_notexitcond201206_push13_notexitcond201206_pop13_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond201206_push13_notexitcond201206_pop13_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond201206_push13_notexitcond201206_pop13_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond201206_push13_notexitcond201206_pop13_output_regs_ready)
		begin
			local_bb4_notexitcond201206_push13_notexitcond201206_pop13_NO_SHIFT_REG <= local_bb4_notexitcond201206_push13_notexitcond201206_pop13_result;
			local_bb4_notexitcond201206_push13_notexitcond201206_pop13_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond201206_push13_notexitcond201206_pop13_stall_in))
			begin
				local_bb4_notexitcond201206_push13_notexitcond201206_pop13_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notexitcond_notexit_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notexitcond_notexit_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_4 = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG = rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_indvars_iv_push7_indvars_iv_next_stall_in = 1'b0;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG = rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_sub17_add16204_push10_sub17_add16204_pop10_inputs_ready;
 reg local_bb4_sub17_add16204_push10_sub17_add16204_pop10_valid_out_NO_SHIFT_REG;
wire local_bb4_sub17_add16204_push10_sub17_add16204_pop10_stall_in;
wire local_bb4_sub17_add16204_push10_sub17_add16204_pop10_output_regs_ready;
wire [31:0] local_bb4_sub17_add16204_push10_sub17_add16204_pop10_result;
wire local_bb4_sub17_add16204_push10_sub17_add16204_pop10_fu_valid_out;
wire local_bb4_sub17_add16204_push10_sub17_add16204_pop10_fu_stall_out;
 reg [31:0] local_bb4_sub17_add16204_push10_sub17_add16204_pop10_NO_SHIFT_REG;
wire local_bb4_sub17_add16204_push10_sub17_add16204_pop10_causedstall;

acl_push local_bb4_sub17_add16204_push10_sub17_add16204_pop10_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_NO_SHIFT_REG),
	.stall_out(local_bb4_sub17_add16204_push10_sub17_add16204_pop10_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sub17_add16204_push10_sub17_add16204_pop10_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_sub17_add16204_push10_sub17_add16204_pop10_result),
	.feedback_out(feedback_data_out_10),
	.feedback_valid_out(feedback_valid_out_10),
	.feedback_stall_in(feedback_stall_in_10)
);

defparam local_bb4_sub17_add16204_push10_sub17_add16204_pop10_feedback.STALLFREE = 1;
defparam local_bb4_sub17_add16204_push10_sub17_add16204_pop10_feedback.DATA_WIDTH = 32;
defparam local_bb4_sub17_add16204_push10_sub17_add16204_pop10_feedback.FIFO_DEPTH = 9;
defparam local_bb4_sub17_add16204_push10_sub17_add16204_pop10_feedback.MIN_FIFO_LATENCY = 8;
defparam local_bb4_sub17_add16204_push10_sub17_add16204_pop10_feedback.STYLE = "REGULAR";

assign local_bb4_sub17_add16204_push10_sub17_add16204_pop10_inputs_ready = 1'b1;
assign local_bb4_sub17_add16204_push10_sub17_add16204_pop10_output_regs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_1 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_5 = 1'b0;
assign rnode_9to10_bb4_sub17_add16204_pop10_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_sub17_add16204_push10_sub17_add16204_pop10_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_sub17_add16204_push10_sub17_add16204_pop10_NO_SHIFT_REG <= 'x;
		local_bb4_sub17_add16204_push10_sub17_add16204_pop10_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_sub17_add16204_push10_sub17_add16204_pop10_output_regs_ready)
		begin
			local_bb4_sub17_add16204_push10_sub17_add16204_pop10_NO_SHIFT_REG <= local_bb4_sub17_add16204_push10_sub17_add16204_pop10_result;
			local_bb4_sub17_add16204_push10_sub17_add16204_pop10_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_sub17_add16204_push10_sub17_add16204_pop10_stall_in))
			begin
				local_bb4_sub17_add16204_push10_sub17_add16204_pop10_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_idxprom24_stall_local;
wire [63:0] local_bb4_idxprom24;

assign local_bb4_idxprom24[63:32] = 32'h0;
assign local_bb4_idxprom24[31:0] = rnode_9to10_bb4_add23_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_arrayidx25_valid_out;
wire local_bb4_arrayidx25_stall_in;
wire local_bb4_arrayidx25_inputs_ready;
wire local_bb4_arrayidx25_stall_local;
wire [63:0] local_bb4_arrayidx25;

assign local_bb4_arrayidx25_inputs_ready = rnode_9to10_bb4_add23_0_valid_out_NO_SHIFT_REG;
assign local_bb4_arrayidx25 = ((input_in & 64'hFFFFFFFFFFFFFC00) + ((local_bb4_idxprom24 & 64'hFFFFFFFF) << 6'h2));
assign local_bb4_arrayidx25_valid_out = 1'b1;
assign rnode_9to10_bb4_add23_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_arrayidx25_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx25_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx25_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx25_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx25_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx25_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx25_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx25_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_arrayidx25_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_arrayidx25_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_arrayidx25_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_arrayidx25_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_arrayidx25_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in((local_bb4_arrayidx25 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_10to11_bb4_arrayidx25_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_arrayidx25_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_arrayidx25_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_arrayidx25_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_arrayidx25_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_arrayidx25_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_arrayidx25_stall_in = 1'b0;
assign rnode_10to11_bb4_arrayidx25_0_NO_SHIFT_REG = rnode_10to11_bb4_arrayidx25_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_arrayidx25_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx25_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi1210_stall_local;
wire [319:0] local_bb4_c0_exi1210;

assign local_bb4_c0_exi1210[63:0] = 64'bx;
assign local_bb4_c0_exi1210[127:64] = (rnode_10to11_bb4_arrayidx25_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign local_bb4_c0_exi1210[319:128] = 192'bx;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi2211_stall_local;
wire [319:0] local_bb4_c0_exi2211;

assign local_bb4_c0_exi2211[127:0] = local_bb4_c0_exi1210[127:0];
assign local_bb4_c0_exi2211[191:128] = rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_NO_SHIFT_REG;
assign local_bb4_c0_exi2211[319:192] = local_bb4_c0_exi1210[319:192];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi3212_stall_local;
wire [319:0] local_bb4_c0_exi3212;

assign local_bb4_c0_exi3212[191:0] = local_bb4_c0_exi2211[191:0];
assign local_bb4_c0_exi3212[255:192] = (rnode_10to11_bb4_arrayidx35_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign local_bb4_c0_exi3212[319:256] = local_bb4_c0_exi2211[319:256];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi4213_stall_local;
wire [319:0] local_bb4_c0_exi4213;

assign local_bb4_c0_exi4213[255:0] = local_bb4_c0_exi3212[255:0];
assign local_bb4_c0_exi4213[256] = rnode_9to11_bb4_var__u27_0_NO_SHIFT_REG;
assign local_bb4_c0_exi4213[319:257] = local_bb4_c0_exi3212[319:257];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi5_stall_local;
wire [319:0] local_bb4_c0_exi5;

assign local_bb4_c0_exi5[263:0] = local_bb4_c0_exi4213[263:0];
assign local_bb4_c0_exi5[264] = rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG;
assign local_bb4_c0_exi5[319:265] = local_bb4_c0_exi4213[319:265];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi6_stall_local;
wire [319:0] local_bb4_c0_exi6;

assign local_bb4_c0_exi6[271:0] = local_bb4_c0_exi5[271:0];
assign local_bb4_c0_exi6[272] = rnode_10to11_bb4__pop12_c0_ene4_0_NO_SHIFT_REG;
assign local_bb4_c0_exi6[319:273] = local_bb4_c0_exi5[319:273];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi7_valid_out;
wire local_bb4_c0_exi7_stall_in;
wire local_bb4_c0_exi7_inputs_ready;
wire local_bb4_c0_exi7_stall_local;
wire [319:0] local_bb4_c0_exi7;

assign local_bb4_c0_exi7_inputs_ready = (rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_arrayidx35_0_valid_out_NO_SHIFT_REG & rnode_9to11_bb4_var__u27_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_arrayidx25_0_valid_out_NO_SHIFT_REG);
assign local_bb4_c0_exi7[279:0] = local_bb4_c0_exi6[279:0];
assign local_bb4_c0_exi7[280] = rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_NO_SHIFT_REG;
assign local_bb4_c0_exi7[319:281] = local_bb4_c0_exi6[319:281];
assign local_bb4_c0_exi7_valid_out = 1'b1;
assign rnode_10to11_bb4_arrayidx32205_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx35_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_var__u27_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond201206_pop13_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx25_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_c0_exit214_c0_exi7_inputs_ready;
 reg local_bb4_c0_exit214_c0_exi7_valid_out_0_NO_SHIFT_REG;
wire local_bb4_c0_exit214_c0_exi7_stall_in_0;
 reg local_bb4_c0_exit214_c0_exi7_valid_out_1_NO_SHIFT_REG;
wire local_bb4_c0_exit214_c0_exi7_stall_in_1;
 reg [319:0] local_bb4_c0_exit214_c0_exi7_NO_SHIFT_REG;
wire [319:0] local_bb4_c0_exit214_c0_exi7_in;
wire local_bb4_c0_exit214_c0_exi7_valid;
wire local_bb4_c0_exit214_c0_exi7_causedstall;

acl_stall_free_sink local_bb4_c0_exit214_c0_exi7_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb4_c0_exi7),
	.data_out(local_bb4_c0_exit214_c0_exi7_in),
	.input_accepted(local_bb4_c0_enter208_c0_eni5_input_accepted),
	.valid_out(local_bb4_c0_exit214_c0_exi7_valid),
	.stall_in(~(local_bb4_c0_exit214_c0_exi7_output_regs_ready)),
	.stall_entry(local_bb4_c0_exit214_c0_exi7_entry_stall),
	.valid_in(local_bb4_c0_exit214_c0_exi7_valid_in),
	.IIphases(local_bb4_c0_exit214_c0_exi7_phases),
	.inc_pipelined_thread(local_bb4_c0_enter208_c0_eni5_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb4_c0_enter208_c0_eni5_dec_pipelined_thread)
);

defparam local_bb4_c0_exit214_c0_exi7_instance.DATA_WIDTH = 320;
defparam local_bb4_c0_exit214_c0_exi7_instance.PIPELINE_DEPTH = 15;
defparam local_bb4_c0_exit214_c0_exi7_instance.SHARINGII = 1;
defparam local_bb4_c0_exit214_c0_exi7_instance.SCHEDULEII = 1;
defparam local_bb4_c0_exit214_c0_exi7_instance.ALWAYS_THROTTLE = 0;

assign local_bb4_c0_exit214_c0_exi7_inputs_ready = 1'b1;
assign local_bb4_c0_exit214_c0_exi7_output_regs_ready = ((~(local_bb4_c0_exit214_c0_exi7_valid_out_0_NO_SHIFT_REG) | ~(local_bb4_c0_exit214_c0_exi7_stall_in_0)) & (~(local_bb4_c0_exit214_c0_exi7_valid_out_1_NO_SHIFT_REG) | ~(local_bb4_c0_exit214_c0_exi7_stall_in_1)));
assign local_bb4_c0_exit214_c0_exi7_valid_in = SFC_2_VALID_10_11_0_NO_SHIFT_REG;
assign local_bb4_c0_exi7_stall_in = 1'b0;
assign local_bb4_arrayidx32205_push11_arrayidx32205_pop11_stall_in = 1'b0;
assign local_bb4_sub17_add16204_push10_sub17_add16204_pop10_stall_in = 1'b0;
assign local_bb4__push12__pop12_stall_in = 1'b0;
assign local_bb4_notexitcond201206_push13_notexitcond201206_pop13_stall_in = 1'b0;
assign SFC_2_VALID_10_11_0_stall_in = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_c0_exit214_c0_exi7_causedstall = (1'b1 && (1'b0 && !(~(local_bb4_c0_exit214_c0_exi7_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c0_exit214_c0_exi7_NO_SHIFT_REG <= 'x;
		local_bb4_c0_exit214_c0_exi7_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_c0_exit214_c0_exi7_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c0_exit214_c0_exi7_output_regs_ready)
		begin
			local_bb4_c0_exit214_c0_exi7_NO_SHIFT_REG <= local_bb4_c0_exit214_c0_exi7_in;
			local_bb4_c0_exit214_c0_exi7_valid_out_0_NO_SHIFT_REG <= local_bb4_c0_exit214_c0_exi7_valid;
			local_bb4_c0_exit214_c0_exi7_valid_out_1_NO_SHIFT_REG <= local_bb4_c0_exit214_c0_exi7_valid;
		end
		else
		begin
			if (~(local_bb4_c0_exit214_c0_exi7_stall_in_0))
			begin
				local_bb4_c0_exit214_c0_exi7_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c0_exit214_c0_exi7_stall_in_1))
			begin
				local_bb4_c0_exit214_c0_exi7_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe1215_valid_out;
wire local_bb4_c0_exe1215_stall_in;
wire local_bb4_c0_exe1215_inputs_ready;
wire local_bb4_c0_exe1215_stall_local;
wire [63:0] local_bb4_c0_exe1215;

assign local_bb4_c0_exe1215_inputs_ready = local_bb4_c0_exit214_c0_exi7_valid_out_0_NO_SHIFT_REG;
assign local_bb4_c0_exe1215 = local_bb4_c0_exit214_c0_exi7_NO_SHIFT_REG[127:64];
assign local_bb4_c0_exe1215_valid_out = local_bb4_c0_exe1215_inputs_ready;
assign local_bb4_c0_exe1215_stall_local = local_bb4_c0_exe1215_stall_in;
assign local_bb4_c0_exit214_c0_exi7_stall_in_0 = (|local_bb4_c0_exe1215_stall_local);

// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_16to178_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG;
 logic rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG;
 logic [319:0] rnode_16to178_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG;
 logic rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [319:0] rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_NO_SHIFT_REG;
 logic rnode_16to178_bb4_c0_exit214_c0_exi7_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_16to178_bb4_c0_exit214_c0_exi7_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_c0_exit214_c0_exi7_NO_SHIFT_REG),
	.data_out(rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_fifo.DEPTH = 163;
defparam rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_fifo.DATA_WIDTH = 320;
defparam rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_fifo.IMPL = "ram";

assign rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_inputs_ready_NO_SHIFT_REG = local_bb4_c0_exit214_c0_exi7_valid_out_1_NO_SHIFT_REG;
assign local_bb4_c0_exit214_c0_exi7_stall_in_1 = rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_out_reg_178_NO_SHIFT_REG;
assign rnode_16to178_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG = rnode_16to178_bb4_c0_exit214_c0_exi7_0_reg_178_NO_SHIFT_REG;
assign rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_in_reg_178_NO_SHIFT_REG = rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG;
assign rnode_16to178_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG = rnode_16to178_bb4_c0_exit214_c0_exi7_0_valid_out_reg_178_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_ld__inputs_ready;
 reg local_bb4_ld__valid_out_NO_SHIFT_REG;
wire local_bb4_ld__stall_in;
wire local_bb4_ld__output_regs_ready;
wire local_bb4_ld__fu_stall_out;
wire local_bb4_ld__fu_valid_out;
wire [31:0] local_bb4_ld__lsu_dataout;
 reg [31:0] local_bb4_ld__NO_SHIFT_REG;
wire local_bb4_ld__causedstall;

lsu_top lsu_local_bb4_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb4_ld__fu_stall_out),
	.i_valid(local_bb4_ld__inputs_ready),
	.i_address((local_bb4_c0_exe1215 & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(local_bb4__acl_ffwd_dest_i1_10),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb4_ld__output_regs_ready)),
	.o_valid(local_bb4_ld__fu_valid_out),
	.o_readdata(local_bb4_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb4_ld__active),
	.avm_address(avm_local_bb4_ld__address),
	.avm_read(avm_local_bb4_ld__read),
	.avm_readdata(avm_local_bb4_ld__readdata),
	.avm_write(avm_local_bb4_ld__write),
	.avm_writeack(avm_local_bb4_ld__writeack),
	.avm_burstcount(avm_local_bb4_ld__burstcount),
	.avm_writedata(avm_local_bb4_ld__writedata),
	.avm_byteenable(avm_local_bb4_ld__byteenable),
	.avm_waitrequest(avm_local_bb4_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb4_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb4_ld_.AWIDTH = 33;
defparam lsu_local_bb4_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb4_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb4_ld_.READ = 1;
defparam lsu_local_bb4_ld_.ATOMIC = 0;
defparam lsu_local_bb4_ld_.WIDTH = 32;
defparam lsu_local_bb4_ld_.MWIDTH = 512;
defparam lsu_local_bb4_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb4_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb4_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb4_ld_.MEMORY_SIDE_MEM_LATENCY = 148;
defparam lsu_local_bb4_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb4_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb4_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb4_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb4_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb4_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb4_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb4_ld_.USECACHING = 0;
defparam lsu_local_bb4_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb4_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb4_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb4_ld_.ADDRSPACE = 1;
defparam lsu_local_bb4_ld_.STYLE = "BURST-COALESCED";

assign local_bb4_ld__inputs_ready = (local_bb4_c0_exe1215_valid_out & local_bb4__acl_ffwd_dest_i1_10_valid_out);
assign local_bb4_ld__output_regs_ready = (&(~(local_bb4_ld__valid_out_NO_SHIFT_REG) | ~(local_bb4_ld__stall_in)));
assign local_bb4_c0_exe1215_stall_in = (local_bb4_ld__fu_stall_out | ~(local_bb4_ld__inputs_ready));
assign local_bb4__acl_ffwd_dest_i1_10_stall_in = (local_bb4_ld__fu_stall_out | ~(local_bb4_ld__inputs_ready));
assign local_bb4_ld__causedstall = (local_bb4_ld__inputs_ready && (local_bb4_ld__fu_stall_out && !(~(local_bb4_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_ld__NO_SHIFT_REG <= 'x;
		local_bb4_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_ld__output_regs_ready)
		begin
			local_bb4_ld__NO_SHIFT_REG <= local_bb4_ld__lsu_dataout;
			local_bb4_ld__valid_out_NO_SHIFT_REG <= local_bb4_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb4_ld__stall_in))
			begin
				local_bb4_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG;
 logic [319:0] rnode_178to179_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG;
 logic [319:0] rnode_178to179_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_2_NO_SHIFT_REG;
 logic [319:0] rnode_178to179_bb4_c0_exit214_c0_exi7_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [319:0] rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_out_reg_179_NO_SHIFT_REG;
 reg rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG;
 reg rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG;
 reg rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_2_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(rnode_16to178_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG),
	.data_out(rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_fifo.DEPTH = 2;
defparam rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_fifo.DATA_WIDTH = 320;
defparam rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_fifo.IMPL = "ll_reg";

assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_inputs_ready_NO_SHIFT_REG = rnode_16to178_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG;
assign rnode_16to178_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG = rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_out_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_179_NO_SHIFT_REG = ((rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG & ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG)) | (rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG & ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG)) | (rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_2_NO_SHIFT_REG & ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_2_NO_SHIFT_REG)));
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG = (rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG & ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG));
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG = (rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG & ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG));
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_2_NO_SHIFT_REG = (rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG & ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_2_NO_SHIFT_REG));
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG = rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG = rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_c0_exit214_c0_exi7_2_NO_SHIFT_REG = rnode_178to179_bb4_c0_exit214_c0_exi7_0_reg_179_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG <= 1'b0;
		rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG <= (rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG & (rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG | ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG)) & rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_179_NO_SHIFT_REG);
		rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG <= (rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG & (rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG | ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG)) & rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_179_NO_SHIFT_REG);
		rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_2_NO_SHIFT_REG <= (rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_179_NO_SHIFT_REG & (rnode_178to179_bb4_c0_exit214_c0_exi7_0_consumed_2_NO_SHIFT_REG | ~(rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_2_NO_SHIFT_REG)) & rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_179_NO_SHIFT_REG);
	end
end


// This section implements a staging register.
// 
wire rstag_176to176_bb4_ld__valid_out_0;
wire rstag_176to176_bb4_ld__stall_in_0;
wire rstag_176to176_bb4_ld__valid_out_1;
wire rstag_176to176_bb4_ld__stall_in_1;
wire rstag_176to176_bb4_ld__inputs_ready;
wire rstag_176to176_bb4_ld__stall_local;
 reg rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG;
wire rstag_176to176_bb4_ld__combined_valid;
 reg [31:0] rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_176to176_bb4_ld_;
 reg rstag_176to176_bb4_ld__consumed_0_NO_SHIFT_REG;
 reg rstag_176to176_bb4_ld__consumed_1_NO_SHIFT_REG;

assign rstag_176to176_bb4_ld__inputs_ready = local_bb4_ld__valid_out_NO_SHIFT_REG;
assign rstag_176to176_bb4_ld_ = (rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG ? rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG : local_bb4_ld__NO_SHIFT_REG);
assign rstag_176to176_bb4_ld__combined_valid = (rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG | rstag_176to176_bb4_ld__inputs_ready);
assign rstag_176to176_bb4_ld__stall_local = ((rstag_176to176_bb4_ld__stall_in_0 & ~(rstag_176to176_bb4_ld__consumed_0_NO_SHIFT_REG)) | (rstag_176to176_bb4_ld__stall_in_1 & ~(rstag_176to176_bb4_ld__consumed_1_NO_SHIFT_REG)));
assign rstag_176to176_bb4_ld__valid_out_0 = (rstag_176to176_bb4_ld__combined_valid & ~(rstag_176to176_bb4_ld__consumed_0_NO_SHIFT_REG));
assign rstag_176to176_bb4_ld__valid_out_1 = (rstag_176to176_bb4_ld__combined_valid & ~(rstag_176to176_bb4_ld__consumed_1_NO_SHIFT_REG));
assign local_bb4_ld__stall_in = (|rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_176to176_bb4_ld__stall_local)
		begin
			if (~(rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= rstag_176to176_bb4_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG <= local_bb4_ld__NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_176to176_bb4_ld__consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_176to176_bb4_ld__consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_176to176_bb4_ld__consumed_0_NO_SHIFT_REG <= (rstag_176to176_bb4_ld__combined_valid & (rstag_176to176_bb4_ld__consumed_0_NO_SHIFT_REG | ~(rstag_176to176_bb4_ld__stall_in_0)) & rstag_176to176_bb4_ld__stall_local);
		rstag_176to176_bb4_ld__consumed_1_NO_SHIFT_REG <= (rstag_176to176_bb4_ld__combined_valid & (rstag_176to176_bb4_ld__consumed_1_NO_SHIFT_REG | ~(rstag_176to176_bb4_ld__stall_in_1)) & rstag_176to176_bb4_ld__stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe2216_valid_out;
wire local_bb4_c0_exe2216_stall_in;
wire local_bb4_c0_exe2216_inputs_ready;
wire local_bb4_c0_exe2216_stall_local;
wire [63:0] local_bb4_c0_exe2216;

assign local_bb4_c0_exe2216_inputs_ready = rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_c0_exe2216 = rnode_178to179_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG[191:128];
assign local_bb4_c0_exe2216_valid_out = local_bb4_c0_exe2216_inputs_ready;
assign local_bb4_c0_exe2216_stall_local = local_bb4_c0_exe2216_stall_in;
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG = (|local_bb4_c0_exe2216_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe3217_valid_out;
wire local_bb4_c0_exe3217_stall_in;
wire local_bb4_c0_exe3217_inputs_ready;
wire local_bb4_c0_exe3217_stall_local;
wire [63:0] local_bb4_c0_exe3217;

assign local_bb4_c0_exe3217_inputs_ready = rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_c0_exe3217 = rnode_178to179_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG[255:192];
assign local_bb4_c0_exe3217_valid_out = local_bb4_c0_exe3217_inputs_ready;
assign local_bb4_c0_exe3217_stall_local = local_bb4_c0_exe3217_stall_in;
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG = (|local_bb4_c0_exe3217_stall_local);

// Register node:
//  * latency = 159
//  * capacity = 159
 logic rnode_179to338_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG;
 logic [319:0] rnode_179to338_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG;
 logic rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [319:0] rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_NO_SHIFT_REG;
 logic rnode_179to338_bb4_c0_exit214_c0_exi7_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_179to338_bb4_c0_exit214_c0_exi7_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(rnode_178to179_bb4_c0_exit214_c0_exi7_2_NO_SHIFT_REG),
	.data_out(rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_fifo.DEPTH = 160;
defparam rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_fifo.DATA_WIDTH = 320;
defparam rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_fifo.IMPL = "ram";

assign rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_inputs_ready_NO_SHIFT_REG = rnode_178to179_bb4_c0_exit214_c0_exi7_0_valid_out_2_NO_SHIFT_REG;
assign rnode_178to179_bb4_c0_exit214_c0_exi7_0_stall_in_2_NO_SHIFT_REG = rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_out_reg_338_NO_SHIFT_REG;
assign rnode_179to338_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG = rnode_179to338_bb4_c0_exit214_c0_exi7_0_reg_338_NO_SHIFT_REG;
assign rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_in_reg_338_NO_SHIFT_REG = rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG;
assign rnode_179to338_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG = rnode_179to338_bb4_c0_exit214_c0_exi7_0_valid_out_reg_338_NO_SHIFT_REG;

// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_176to338_bb4_ld__0_valid_out_NO_SHIFT_REG;
 logic rnode_176to338_bb4_ld__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to338_bb4_ld__0_NO_SHIFT_REG;
 logic rnode_176to338_bb4_ld__0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to338_bb4_ld__0_reg_338_NO_SHIFT_REG;
 logic rnode_176to338_bb4_ld__0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_176to338_bb4_ld__0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_176to338_bb4_ld__0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_176to338_bb4_ld__0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to338_bb4_ld__0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to338_bb4_ld__0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_176to338_bb4_ld__0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_176to338_bb4_ld__0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(rstag_176to176_bb4_ld_),
	.data_out(rnode_176to338_bb4_ld__0_reg_338_NO_SHIFT_REG)
);

defparam rnode_176to338_bb4_ld__0_reg_338_fifo.DEPTH = 163;
defparam rnode_176to338_bb4_ld__0_reg_338_fifo.DATA_WIDTH = 32;
defparam rnode_176to338_bb4_ld__0_reg_338_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_176to338_bb4_ld__0_reg_338_fifo.IMPL = "ram";

assign rnode_176to338_bb4_ld__0_reg_338_inputs_ready_NO_SHIFT_REG = rstag_176to176_bb4_ld__valid_out_0;
assign rstag_176to176_bb4_ld__stall_in_0 = rnode_176to338_bb4_ld__0_stall_out_reg_338_NO_SHIFT_REG;
assign rnode_176to338_bb4_ld__0_NO_SHIFT_REG = rnode_176to338_bb4_ld__0_reg_338_NO_SHIFT_REG;
assign rnode_176to338_bb4_ld__0_stall_in_reg_338_NO_SHIFT_REG = rnode_176to338_bb4_ld__0_stall_in_NO_SHIFT_REG;
assign rnode_176to338_bb4_ld__0_valid_out_NO_SHIFT_REG = rnode_176to338_bb4_ld__0_valid_out_reg_338_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_cmp26_inputs_ready;
 reg local_bb4_cmp26_valid_out_NO_SHIFT_REG;
wire local_bb4_cmp26_stall_in;
wire local_bb4_cmp26_output_regs_ready;
wire local_bb4_cmp26;
 reg local_bb4_cmp26_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_cmp26_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_cmp26_causedstall;

acl_fp_cmp fp_module_local_bb4_cmp26 (
	.clock(clock),
	.dataa(rstag_176to176_bb4_ld_),
	.datab(32'h0),
	.enable(local_bb4_cmp26_output_regs_ready),
	.result(local_bb4_cmp26)
);

defparam fp_module_local_bb4_cmp26.COMPARISON_MODE = 3;

assign local_bb4_cmp26_inputs_ready = rstag_176to176_bb4_ld__valid_out_1;
assign local_bb4_cmp26_output_regs_ready = (&(~(local_bb4_cmp26_valid_out_NO_SHIFT_REG) | ~(local_bb4_cmp26_stall_in)));
assign rstag_176to176_bb4_ld__stall_in_1 = (~(local_bb4_cmp26_output_regs_ready) | ~(local_bb4_cmp26_inputs_ready));
assign local_bb4_cmp26_causedstall = (local_bb4_cmp26_inputs_ready && (~(local_bb4_cmp26_output_regs_ready) && !(~(local_bb4_cmp26_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_cmp26_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_cmp26_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_cmp26_output_regs_ready)
		begin
			local_bb4_cmp26_valid_pipe_0_NO_SHIFT_REG <= local_bb4_cmp26_inputs_ready;
			local_bb4_cmp26_valid_pipe_1_NO_SHIFT_REG <= local_bb4_cmp26_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_cmp26_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_cmp26_output_regs_ready)
		begin
			local_bb4_cmp26_valid_out_NO_SHIFT_REG <= local_bb4_cmp26_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb4_cmp26_stall_in))
			begin
				local_bb4_cmp26_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG;
 logic [319:0] rnode_338to339_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG;
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG;
 logic [319:0] rnode_338to339_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG;
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic [319:0] rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_339_NO_SHIFT_REG;
 logic rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_out_reg_339_NO_SHIFT_REG;
 reg rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG;
 reg rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_339_NO_SHIFT_REG),
	.valid_out(rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_339_NO_SHIFT_REG),
	.stall_out(rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_out_reg_339_NO_SHIFT_REG),
	.data_in(rnode_179to338_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG),
	.data_out(rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_NO_SHIFT_REG)
);

defparam rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_fifo.DEPTH = 1;
defparam rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_fifo.DATA_WIDTH = 320;
defparam rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_fifo.IMPL = "ll_reg";

assign rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_inputs_ready_NO_SHIFT_REG = rnode_179to338_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG;
assign rnode_179to338_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG = rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_out_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_339_NO_SHIFT_REG = ((rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG & ~(rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG)) | (rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG & ~(rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG)));
assign rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG = (rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_339_NO_SHIFT_REG & ~(rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG));
assign rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG = (rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_339_NO_SHIFT_REG & ~(rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG));
assign rnode_338to339_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG = rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_NO_SHIFT_REG;
assign rnode_338to339_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG = rnode_338to339_bb4_c0_exit214_c0_exi7_0_reg_339_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG <= (rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_339_NO_SHIFT_REG & (rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_0_NO_SHIFT_REG | ~(rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG)) & rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_339_NO_SHIFT_REG);
		rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG <= (rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_339_NO_SHIFT_REG & (rnode_338to339_bb4_c0_exit214_c0_exi7_0_consumed_1_NO_SHIFT_REG | ~(rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG)) & rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_339_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_179to179_bb4_cmp26_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_1_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_reg_179_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_179to179_bb4_cmp26_0_stall_out_reg_179_NO_SHIFT_REG;
 reg rnode_179to179_bb4_cmp26_0_consumed_0_NO_SHIFT_REG;
 reg rnode_179to179_bb4_cmp26_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_179to179_bb4_cmp26_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to179_bb4_cmp26_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to179_bb4_cmp26_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_179to179_bb4_cmp26_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_179to179_bb4_cmp26_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4_cmp26),
	.data_out(rnode_179to179_bb4_cmp26_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_179to179_bb4_cmp26_0_reg_179_fifo.DEPTH = 3;
defparam rnode_179to179_bb4_cmp26_0_reg_179_fifo.DATA_WIDTH = 1;
defparam rnode_179to179_bb4_cmp26_0_reg_179_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_179to179_bb4_cmp26_0_reg_179_fifo.IMPL = "zl_reg";

assign rnode_179to179_bb4_cmp26_0_reg_179_inputs_ready_NO_SHIFT_REG = local_bb4_cmp26_valid_out_NO_SHIFT_REG;
assign local_bb4_cmp26_stall_in = rnode_179to179_bb4_cmp26_0_stall_out_reg_179_NO_SHIFT_REG;
assign rnode_179to179_bb4_cmp26_0_stall_in_0_reg_179_NO_SHIFT_REG = ((rnode_179to179_bb4_cmp26_0_stall_in_0_NO_SHIFT_REG & ~(rnode_179to179_bb4_cmp26_0_consumed_0_NO_SHIFT_REG)) | (rnode_179to179_bb4_cmp26_0_stall_in_1_NO_SHIFT_REG & ~(rnode_179to179_bb4_cmp26_0_consumed_1_NO_SHIFT_REG)));
assign rnode_179to179_bb4_cmp26_0_valid_out_0_NO_SHIFT_REG = (rnode_179to179_bb4_cmp26_0_valid_out_0_reg_179_NO_SHIFT_REG & ~(rnode_179to179_bb4_cmp26_0_consumed_0_NO_SHIFT_REG));
assign rnode_179to179_bb4_cmp26_0_valid_out_1_NO_SHIFT_REG = (rnode_179to179_bb4_cmp26_0_valid_out_0_reg_179_NO_SHIFT_REG & ~(rnode_179to179_bb4_cmp26_0_consumed_1_NO_SHIFT_REG));
assign rnode_179to179_bb4_cmp26_0_NO_SHIFT_REG = rnode_179to179_bb4_cmp26_0_reg_179_NO_SHIFT_REG;
assign rnode_179to179_bb4_cmp26_1_NO_SHIFT_REG = rnode_179to179_bb4_cmp26_0_reg_179_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_179to179_bb4_cmp26_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_179to179_bb4_cmp26_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_179to179_bb4_cmp26_0_consumed_0_NO_SHIFT_REG <= (rnode_179to179_bb4_cmp26_0_valid_out_0_reg_179_NO_SHIFT_REG & (rnode_179to179_bb4_cmp26_0_consumed_0_NO_SHIFT_REG | ~(rnode_179to179_bb4_cmp26_0_stall_in_0_NO_SHIFT_REG)) & rnode_179to179_bb4_cmp26_0_stall_in_0_reg_179_NO_SHIFT_REG);
		rnode_179to179_bb4_cmp26_0_consumed_1_NO_SHIFT_REG <= (rnode_179to179_bb4_cmp26_0_valid_out_0_reg_179_NO_SHIFT_REG & (rnode_179to179_bb4_cmp26_0_consumed_1_NO_SHIFT_REG | ~(rnode_179to179_bb4_cmp26_0_stall_in_1_NO_SHIFT_REG)) & rnode_179to179_bb4_cmp26_0_stall_in_0_reg_179_NO_SHIFT_REG);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe5_stall_local;
wire local_bb4_c0_exe5;

assign local_bb4_c0_exe5 = rnode_338to339_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG[264];

// Register node:
//  * latency = 68
//  * capacity = 68
 logic rnode_339to407_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG;
 logic rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG;
 logic [319:0] rnode_339to407_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG;
 logic rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_inputs_ready_NO_SHIFT_REG;
 logic [319:0] rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_NO_SHIFT_REG;
 logic rnode_339to407_bb4_c0_exit214_c0_exi7_0_valid_out_reg_407_NO_SHIFT_REG;
 logic rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_in_reg_407_NO_SHIFT_REG;
 logic rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_out_reg_407_NO_SHIFT_REG;

acl_data_fifo rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_in_reg_407_NO_SHIFT_REG),
	.valid_out(rnode_339to407_bb4_c0_exit214_c0_exi7_0_valid_out_reg_407_NO_SHIFT_REG),
	.stall_out(rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_out_reg_407_NO_SHIFT_REG),
	.data_in(rnode_338to339_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG),
	.data_out(rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_NO_SHIFT_REG)
);

defparam rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_fifo.DEPTH = 69;
defparam rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_fifo.DATA_WIDTH = 320;
defparam rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_fifo.IMPL = "ram";

assign rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_inputs_ready_NO_SHIFT_REG = rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG;
assign rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG = rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_out_reg_407_NO_SHIFT_REG;
assign rnode_339to407_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG = rnode_339to407_bb4_c0_exit214_c0_exi7_0_reg_407_NO_SHIFT_REG;
assign rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_in_reg_407_NO_SHIFT_REG = rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG;
assign rnode_339to407_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG = rnode_339to407_bb4_c0_exit214_c0_exi7_0_valid_out_reg_407_NO_SHIFT_REG;

// Register node:
//  * latency = 159
//  * capacity = 159
 logic rnode_179to338_bb4_cmp26_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to338_bb4_cmp26_0_stall_in_NO_SHIFT_REG;
 logic rnode_179to338_bb4_cmp26_0_NO_SHIFT_REG;
 logic rnode_179to338_bb4_cmp26_0_reg_338_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to338_bb4_cmp26_0_reg_338_NO_SHIFT_REG;
 logic rnode_179to338_bb4_cmp26_0_valid_out_reg_338_NO_SHIFT_REG;
 logic rnode_179to338_bb4_cmp26_0_stall_in_reg_338_NO_SHIFT_REG;
 logic rnode_179to338_bb4_cmp26_0_stall_out_reg_338_NO_SHIFT_REG;

acl_data_fifo rnode_179to338_bb4_cmp26_0_reg_338_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to338_bb4_cmp26_0_reg_338_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to338_bb4_cmp26_0_stall_in_reg_338_NO_SHIFT_REG),
	.valid_out(rnode_179to338_bb4_cmp26_0_valid_out_reg_338_NO_SHIFT_REG),
	.stall_out(rnode_179to338_bb4_cmp26_0_stall_out_reg_338_NO_SHIFT_REG),
	.data_in(rnode_179to179_bb4_cmp26_0_NO_SHIFT_REG),
	.data_out(rnode_179to338_bb4_cmp26_0_reg_338_NO_SHIFT_REG)
);

defparam rnode_179to338_bb4_cmp26_0_reg_338_fifo.DEPTH = 160;
defparam rnode_179to338_bb4_cmp26_0_reg_338_fifo.DATA_WIDTH = 1;
defparam rnode_179to338_bb4_cmp26_0_reg_338_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_179to338_bb4_cmp26_0_reg_338_fifo.IMPL = "ram";

assign rnode_179to338_bb4_cmp26_0_reg_338_inputs_ready_NO_SHIFT_REG = rnode_179to179_bb4_cmp26_0_valid_out_0_NO_SHIFT_REG;
assign rnode_179to179_bb4_cmp26_0_stall_in_0_NO_SHIFT_REG = rnode_179to338_bb4_cmp26_0_stall_out_reg_338_NO_SHIFT_REG;
assign rnode_179to338_bb4_cmp26_0_NO_SHIFT_REG = rnode_179to338_bb4_cmp26_0_reg_338_NO_SHIFT_REG;
assign rnode_179to338_bb4_cmp26_0_stall_in_reg_338_NO_SHIFT_REG = rnode_179to338_bb4_cmp26_0_stall_in_NO_SHIFT_REG;
assign rnode_179to338_bb4_cmp26_0_valid_out_NO_SHIFT_REG = rnode_179to338_bb4_cmp26_0_valid_out_reg_338_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp26_xor_stall_local;
wire local_bb4_cmp26_xor;

assign local_bb4_cmp26_xor = (rnode_179to179_bb4_cmp26_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG;
 logic [319:0] rnode_407to408_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG;
 logic [319:0] rnode_407to408_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_2_NO_SHIFT_REG;
 logic [319:0] rnode_407to408_bb4_c0_exit214_c0_exi7_2_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_inputs_ready_NO_SHIFT_REG;
 logic [319:0] rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_408_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_408_NO_SHIFT_REG;
 logic rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_out_reg_408_NO_SHIFT_REG;
wire [97:0] rci_rcnode_338to339_rc0_t_313_0_reg_338;

acl_data_fifo rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_408_NO_SHIFT_REG),
	.valid_out(rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_408_NO_SHIFT_REG),
	.stall_out(rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_out_reg_408_NO_SHIFT_REG),
	.data_in(rnode_339to407_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG),
	.data_out(rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_NO_SHIFT_REG)
);

defparam rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_fifo.DEPTH = 1;
defparam rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_fifo.DATA_WIDTH = 320;
defparam rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_fifo.IMPL = "ll_reg";

assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_inputs_ready_NO_SHIFT_REG = rnode_339to407_bb4_c0_exit214_c0_exi7_0_valid_out_NO_SHIFT_REG;
assign rnode_339to407_bb4_c0_exit214_c0_exi7_0_stall_in_NO_SHIFT_REG = rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_out_reg_408_NO_SHIFT_REG;
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_0_reg_408_NO_SHIFT_REG = (rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG | rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG | rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_2_NO_SHIFT_REG);
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG = rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_408_NO_SHIFT_REG;
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG = rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_408_NO_SHIFT_REG;
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_2_NO_SHIFT_REG = rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_reg_408_NO_SHIFT_REG;
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG = rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_NO_SHIFT_REG;
assign rnode_407to408_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG = rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_NO_SHIFT_REG;
assign rnode_407to408_bb4_c0_exit214_c0_exi7_2_NO_SHIFT_REG = rnode_407to408_bb4_c0_exit214_c0_exi7_0_reg_408_NO_SHIFT_REG;
assign rci_rcnode_338to339_rc0_t_313_0_reg_338[31:0] = rcnode_1to338_rc7_t_313_0_NO_SHIFT_REG[31:0];
assign rci_rcnode_338to339_rc0_t_313_0_reg_338[32] = rcnode_1to338_rc7_t_313_0_NO_SHIFT_REG[32];
assign rci_rcnode_338to339_rc0_t_313_0_reg_338[64:33] = rcnode_1to338_rc7_t_313_0_NO_SHIFT_REG[64:33];
assign rci_rcnode_338to339_rc0_t_313_0_reg_338[65] = rnode_179to338_bb4_cmp26_0_NO_SHIFT_REG;
assign rci_rcnode_338to339_rc0_t_313_0_reg_338[97:66] = rnode_176to338_bb4_ld__0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_338to339_rc0_t_313_0_valid_out_0_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_in_0_NO_SHIFT_REG;
 logic [97:0] rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_valid_out_1_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_in_1_NO_SHIFT_REG;
 logic [97:0] rcnode_338to339_rc0_t_313_1_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_valid_out_2_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_in_2_NO_SHIFT_REG;
 logic [97:0] rcnode_338to339_rc0_t_313_2_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_valid_out_3_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_in_3_NO_SHIFT_REG;
 logic [97:0] rcnode_338to339_rc0_t_313_3_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_valid_out_4_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_in_4_NO_SHIFT_REG;
 logic [97:0] rcnode_338to339_rc0_t_313_4_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_valid_out_5_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_in_5_NO_SHIFT_REG;
 logic [97:0] rcnode_338to339_rc0_t_313_5_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_reg_339_inputs_ready_NO_SHIFT_REG;
 logic [97:0] rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_in_0_reg_339_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_IP_NO_SHIFT_REG;
 logic rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_NO_SHIFT_REG;

acl_data_fifo rcnode_338to339_rc0_t_313_0_reg_339_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_338to339_rc0_t_313_0_reg_339_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_338to339_rc0_t_313_0_stall_in_0_reg_339_NO_SHIFT_REG),
	.valid_out(rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG),
	.stall_out(rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_338to339_rc0_t_313_0_reg_338),
	.data_out(rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG)
);

defparam rcnode_338to339_rc0_t_313_0_reg_339_fifo.DEPTH = 1;
defparam rcnode_338to339_rc0_t_313_0_reg_339_fifo.DATA_WIDTH = 98;
defparam rcnode_338to339_rc0_t_313_0_reg_339_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_338to339_rc0_t_313_0_reg_339_fifo.IMPL = "ll_reg";

assign rcnode_338to339_rc0_t_313_0_reg_339_inputs_ready_NO_SHIFT_REG = (rnode_179to338_bb4_cmp26_0_valid_out_NO_SHIFT_REG & rnode_176to338_bb4_ld__0_valid_out_NO_SHIFT_REG & rcnode_1to338_rc7_t_313_0_valid_out_NO_SHIFT_REG);
assign rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_NO_SHIFT_REG = (~(rcnode_338to339_rc0_t_313_0_reg_339_inputs_ready_NO_SHIFT_REG) | rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_IP_NO_SHIFT_REG);
assign rnode_179to338_bb4_cmp26_0_stall_in_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_NO_SHIFT_REG;
assign rnode_176to338_bb4_ld__0_stall_in_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_1to338_rc7_t_313_0_stall_in_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_stall_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_0_stall_in_0_reg_339_NO_SHIFT_REG = (rcnode_338to339_rc0_t_313_0_stall_in_0_NO_SHIFT_REG | rcnode_338to339_rc0_t_313_0_stall_in_1_NO_SHIFT_REG | rcnode_338to339_rc0_t_313_0_stall_in_2_NO_SHIFT_REG | rcnode_338to339_rc0_t_313_0_stall_in_3_NO_SHIFT_REG | rcnode_338to339_rc0_t_313_0_stall_in_4_NO_SHIFT_REG | rcnode_338to339_rc0_t_313_0_stall_in_5_NO_SHIFT_REG);
assign rcnode_338to339_rc0_t_313_0_valid_out_0_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_0_valid_out_1_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_0_valid_out_2_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_0_valid_out_3_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_0_valid_out_4_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_0_valid_out_5_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_valid_out_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_1_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_2_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_3_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_4_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG;
assign rcnode_338to339_rc0_t_313_5_NO_SHIFT_REG = rcnode_338to339_rc0_t_313_0_reg_339_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__phi_decision101_or102_valid_out;
wire local_bb4__phi_decision101_or102_stall_in;
wire local_bb4__phi_decision101_or102_inputs_ready;
wire local_bb4__phi_decision101_or102_stall_local;
wire local_bb4__phi_decision101_or102;

assign local_bb4__phi_decision101_or102_inputs_ready = (rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_valid_out_NO_SHIFT_REG & rnode_179to179_bb4_cmp26_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4__phi_decision101_or102 = (local_bb4__acl_ffwd_dest_i1_10_u21 | local_bb4_cmp26_xor);
assign local_bb4__phi_decision101_or102_valid_out = local_bb4__phi_decision101_or102_inputs_ready;
assign local_bb4__phi_decision101_or102_stall_local = local_bb4__phi_decision101_or102_stall_in;
assign rnode_178to179_bb4__acl_ffwd_dest_i1_10_u21_0_stall_in_NO_SHIFT_REG = (local_bb4__phi_decision101_or102_stall_local | ~(local_bb4__phi_decision101_or102_inputs_ready));
assign rnode_179to179_bb4_cmp26_0_stall_in_1_NO_SHIFT_REG = (local_bb4__phi_decision101_or102_stall_local | ~(local_bb4__phi_decision101_or102_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe4218_stall_local;
wire local_bb4_c0_exe4218;

assign local_bb4_c0_exe4218 = rnode_407to408_bb4_c0_exit214_c0_exi7_0_NO_SHIFT_REG[256];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe7_valid_out;
wire local_bb4_c0_exe7_stall_in;
wire local_bb4_c0_exe4218_valid_out;
wire local_bb4_c0_exe4218_stall_in;
wire local_bb4_c0_exe7_inputs_ready;
wire local_bb4_c0_exe7_stall_local;
wire local_bb4_c0_exe7;

assign local_bb4_c0_exe7_inputs_ready = (rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_1_NO_SHIFT_REG & rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_c0_exe7 = rnode_407to408_bb4_c0_exit214_c0_exi7_1_NO_SHIFT_REG[280];
assign local_bb4_c0_exe7_stall_local = (local_bb4_c0_exe7_stall_in | local_bb4_c0_exe4218_stall_in);
assign local_bb4_c0_exe7_valid_out = local_bb4_c0_exe7_inputs_ready;
assign local_bb4_c0_exe4218_valid_out = local_bb4_c0_exe7_inputs_ready;
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_1_NO_SHIFT_REG = (local_bb4_c0_exe7_stall_local | ~(local_bb4_c0_exe7_inputs_ready));
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c0_exe7_stall_local | ~(local_bb4_c0_exe7_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni1_stall_local;
wire [255:0] local_bb4_c1_eni1;

assign local_bb4_c1_eni1[31:0] = 32'bx;
assign local_bb4_c1_eni1[63:32] = rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG[97:66];
assign local_bb4_c1_eni1[255:64] = 192'bx;

// This section implements a staging register.
// 
wire rstag_179to179_bb4__phi_decision101_or102_valid_out_0;
wire rstag_179to179_bb4__phi_decision101_or102_stall_in_0;
wire rstag_179to179_bb4__phi_decision101_or102_valid_out_1;
wire rstag_179to179_bb4__phi_decision101_or102_stall_in_1;
wire rstag_179to179_bb4__phi_decision101_or102_inputs_ready;
wire rstag_179to179_bb4__phi_decision101_or102_stall_local;
 reg rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG;
wire rstag_179to179_bb4__phi_decision101_or102_combined_valid;
 reg rstag_179to179_bb4__phi_decision101_or102_staging_reg_NO_SHIFT_REG;
wire rstag_179to179_bb4__phi_decision101_or102;
 reg rstag_179to179_bb4__phi_decision101_or102_consumed_0_NO_SHIFT_REG;
 reg rstag_179to179_bb4__phi_decision101_or102_consumed_1_NO_SHIFT_REG;

assign rstag_179to179_bb4__phi_decision101_or102_inputs_ready = local_bb4__phi_decision101_or102_valid_out;
assign rstag_179to179_bb4__phi_decision101_or102 = (rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG ? rstag_179to179_bb4__phi_decision101_or102_staging_reg_NO_SHIFT_REG : local_bb4__phi_decision101_or102);
assign rstag_179to179_bb4__phi_decision101_or102_combined_valid = (rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG | rstag_179to179_bb4__phi_decision101_or102_inputs_ready);
assign rstag_179to179_bb4__phi_decision101_or102_stall_local = ((rstag_179to179_bb4__phi_decision101_or102_stall_in_0 & ~(rstag_179to179_bb4__phi_decision101_or102_consumed_0_NO_SHIFT_REG)) | (rstag_179to179_bb4__phi_decision101_or102_stall_in_1 & ~(rstag_179to179_bb4__phi_decision101_or102_consumed_1_NO_SHIFT_REG)));
assign rstag_179to179_bb4__phi_decision101_or102_valid_out_0 = (rstag_179to179_bb4__phi_decision101_or102_combined_valid & ~(rstag_179to179_bb4__phi_decision101_or102_consumed_0_NO_SHIFT_REG));
assign rstag_179to179_bb4__phi_decision101_or102_valid_out_1 = (rstag_179to179_bb4__phi_decision101_or102_combined_valid & ~(rstag_179to179_bb4__phi_decision101_or102_consumed_1_NO_SHIFT_REG));
assign local_bb4__phi_decision101_or102_stall_in = (|rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_179to179_bb4__phi_decision101_or102_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_179to179_bb4__phi_decision101_or102_stall_local)
		begin
			if (~(rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG))
			begin
				rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG <= rstag_179to179_bb4__phi_decision101_or102_inputs_ready;
			end
		end
		else
		begin
			rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_179to179_bb4__phi_decision101_or102_staging_valid_NO_SHIFT_REG))
		begin
			rstag_179to179_bb4__phi_decision101_or102_staging_reg_NO_SHIFT_REG <= local_bb4__phi_decision101_or102;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_179to179_bb4__phi_decision101_or102_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_179to179_bb4__phi_decision101_or102_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_179to179_bb4__phi_decision101_or102_consumed_0_NO_SHIFT_REG <= (rstag_179to179_bb4__phi_decision101_or102_combined_valid & (rstag_179to179_bb4__phi_decision101_or102_consumed_0_NO_SHIFT_REG | ~(rstag_179to179_bb4__phi_decision101_or102_stall_in_0)) & rstag_179to179_bb4__phi_decision101_or102_stall_local);
		rstag_179to179_bb4__phi_decision101_or102_consumed_1_NO_SHIFT_REG <= (rstag_179to179_bb4__phi_decision101_or102_combined_valid & (rstag_179to179_bb4__phi_decision101_or102_consumed_1_NO_SHIFT_REG | ~(rstag_179to179_bb4__phi_decision101_or102_stall_in_1)) & rstag_179to179_bb4__phi_decision101_or102_stall_local);
	end
end


// This section implements a registered operation.
// 
wire local_bb4_ld__u28_inputs_ready;
 reg local_bb4_ld__u28_valid_out_NO_SHIFT_REG;
wire local_bb4_ld__u28_stall_in;
wire local_bb4_ld__u28_output_regs_ready;
wire local_bb4_ld__u28_fu_stall_out;
wire local_bb4_ld__u28_fu_valid_out;
wire [31:0] local_bb4_ld__u28_lsu_dataout;
 reg [31:0] local_bb4_ld__u28_NO_SHIFT_REG;
wire local_bb4_ld__u28_causedstall;

lsu_top lsu_local_bb4_ld__u28 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb4_ld__u28_fu_stall_out),
	.i_valid(local_bb4_ld__u28_inputs_ready),
	.i_address((local_bb4_c0_exe3217 & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_179to179_bb4__phi_decision101_or102),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb4_ld__u28_output_regs_ready)),
	.o_valid(local_bb4_ld__u28_fu_valid_out),
	.o_readdata(local_bb4_ld__u28_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb4_ld__u28_active),
	.avm_address(avm_local_bb4_ld__u28_address),
	.avm_read(avm_local_bb4_ld__u28_read),
	.avm_readdata(avm_local_bb4_ld__u28_readdata),
	.avm_write(avm_local_bb4_ld__u28_write),
	.avm_writeack(avm_local_bb4_ld__u28_writeack),
	.avm_burstcount(avm_local_bb4_ld__u28_burstcount),
	.avm_writedata(avm_local_bb4_ld__u28_writedata),
	.avm_byteenable(avm_local_bb4_ld__u28_byteenable),
	.avm_waitrequest(avm_local_bb4_ld__u28_waitrequest),
	.avm_readdatavalid(avm_local_bb4_ld__u28_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb4_ld__u28.AWIDTH = 33;
defparam lsu_local_bb4_ld__u28.WIDTH_BYTES = 4;
defparam lsu_local_bb4_ld__u28.MWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld__u28.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld__u28.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb4_ld__u28.READ = 1;
defparam lsu_local_bb4_ld__u28.ATOMIC = 0;
defparam lsu_local_bb4_ld__u28.WIDTH = 32;
defparam lsu_local_bb4_ld__u28.MWIDTH = 512;
defparam lsu_local_bb4_ld__u28.ATOMIC_WIDTH = 3;
defparam lsu_local_bb4_ld__u28.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb4_ld__u28.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb4_ld__u28.MEMORY_SIDE_MEM_LATENCY = 148;
defparam lsu_local_bb4_ld__u28.USE_WRITE_ACK = 0;
defparam lsu_local_bb4_ld__u28.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb4_ld__u28.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb4_ld__u28.NUMBER_BANKS = 1;
defparam lsu_local_bb4_ld__u28.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb4_ld__u28.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb4_ld__u28.USEINPUTFIFO = 0;
defparam lsu_local_bb4_ld__u28.USECACHING = 0;
defparam lsu_local_bb4_ld__u28.USEOUTPUTFIFO = 1;
defparam lsu_local_bb4_ld__u28.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb4_ld__u28.HIGH_FMAX = 1;
defparam lsu_local_bb4_ld__u28.ADDRSPACE = 1;
defparam lsu_local_bb4_ld__u28.STYLE = "BURST-COALESCED";

assign local_bb4_ld__u28_inputs_ready = (local_bb4_c0_exe3217_valid_out & rstag_179to179_bb4__phi_decision101_or102_valid_out_0);
assign local_bb4_ld__u28_output_regs_ready = (&(~(local_bb4_ld__u28_valid_out_NO_SHIFT_REG) | ~(local_bb4_ld__u28_stall_in)));
assign local_bb4_c0_exe3217_stall_in = (local_bb4_ld__u28_fu_stall_out | ~(local_bb4_ld__u28_inputs_ready));
assign rstag_179to179_bb4__phi_decision101_or102_stall_in_0 = (local_bb4_ld__u28_fu_stall_out | ~(local_bb4_ld__u28_inputs_ready));
assign local_bb4_ld__u28_causedstall = (local_bb4_ld__u28_inputs_ready && (local_bb4_ld__u28_fu_stall_out && !(~(local_bb4_ld__u28_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_ld__u28_NO_SHIFT_REG <= 'x;
		local_bb4_ld__u28_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_ld__u28_output_regs_ready)
		begin
			local_bb4_ld__u28_NO_SHIFT_REG <= local_bb4_ld__u28_lsu_dataout;
			local_bb4_ld__u28_valid_out_NO_SHIFT_REG <= local_bb4_ld__u28_fu_valid_out;
		end
		else
		begin
			if (~(local_bb4_ld__u28_stall_in))
			begin
				local_bb4_ld__u28_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_ld__u29_inputs_ready;
 reg local_bb4_ld__u29_valid_out_NO_SHIFT_REG;
wire local_bb4_ld__u29_stall_in;
wire local_bb4_ld__u29_output_regs_ready;
wire local_bb4_ld__u29_fu_stall_out;
wire local_bb4_ld__u29_fu_valid_out;
wire [31:0] local_bb4_ld__u29_lsu_dataout;
 reg [31:0] local_bb4_ld__u29_NO_SHIFT_REG;
wire local_bb4_ld__u29_causedstall;

lsu_top lsu_local_bb4_ld__u29 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb4_ld__u29_fu_stall_out),
	.i_valid(local_bb4_ld__u29_inputs_ready),
	.i_address(local_bb4_c0_exe2216),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_179to179_bb4__phi_decision101_or102),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb4_ld__u29_output_regs_ready)),
	.o_valid(local_bb4_ld__u29_fu_valid_out),
	.o_readdata(local_bb4_ld__u29_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb4_ld__u29_active),
	.avm_address(avm_local_bb4_ld__u29_address),
	.avm_read(avm_local_bb4_ld__u29_read),
	.avm_readdata(avm_local_bb4_ld__u29_readdata),
	.avm_write(avm_local_bb4_ld__u29_write),
	.avm_writeack(avm_local_bb4_ld__u29_writeack),
	.avm_burstcount(avm_local_bb4_ld__u29_burstcount),
	.avm_writedata(avm_local_bb4_ld__u29_writedata),
	.avm_byteenable(avm_local_bb4_ld__u29_byteenable),
	.avm_waitrequest(avm_local_bb4_ld__u29_waitrequest),
	.avm_readdatavalid(avm_local_bb4_ld__u29_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb4_ld__u29.AWIDTH = 33;
defparam lsu_local_bb4_ld__u29.WIDTH_BYTES = 4;
defparam lsu_local_bb4_ld__u29.MWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld__u29.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld__u29.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb4_ld__u29.READ = 1;
defparam lsu_local_bb4_ld__u29.ATOMIC = 0;
defparam lsu_local_bb4_ld__u29.WIDTH = 32;
defparam lsu_local_bb4_ld__u29.MWIDTH = 512;
defparam lsu_local_bb4_ld__u29.ATOMIC_WIDTH = 3;
defparam lsu_local_bb4_ld__u29.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb4_ld__u29.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb4_ld__u29.MEMORY_SIDE_MEM_LATENCY = 148;
defparam lsu_local_bb4_ld__u29.USE_WRITE_ACK = 0;
defparam lsu_local_bb4_ld__u29.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb4_ld__u29.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb4_ld__u29.NUMBER_BANKS = 1;
defparam lsu_local_bb4_ld__u29.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb4_ld__u29.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb4_ld__u29.USEINPUTFIFO = 0;
defparam lsu_local_bb4_ld__u29.USECACHING = 0;
defparam lsu_local_bb4_ld__u29.USEOUTPUTFIFO = 1;
defparam lsu_local_bb4_ld__u29.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb4_ld__u29.HIGH_FMAX = 1;
defparam lsu_local_bb4_ld__u29.ADDRSPACE = 1;
defparam lsu_local_bb4_ld__u29.STYLE = "BURST-COALESCED";

assign local_bb4_ld__u29_inputs_ready = (local_bb4_c0_exe2216_valid_out & rstag_179to179_bb4__phi_decision101_or102_valid_out_1);
assign local_bb4_ld__u29_output_regs_ready = (&(~(local_bb4_ld__u29_valid_out_NO_SHIFT_REG) | ~(local_bb4_ld__u29_stall_in)));
assign local_bb4_c0_exe2216_stall_in = (local_bb4_ld__u29_fu_stall_out | ~(local_bb4_ld__u29_inputs_ready));
assign rstag_179to179_bb4__phi_decision101_or102_stall_in_1 = (local_bb4_ld__u29_fu_stall_out | ~(local_bb4_ld__u29_inputs_ready));
assign local_bb4_ld__u29_causedstall = (local_bb4_ld__u29_inputs_ready && (local_bb4_ld__u29_fu_stall_out && !(~(local_bb4_ld__u29_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_ld__u29_NO_SHIFT_REG <= 'x;
		local_bb4_ld__u29_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_ld__u29_output_regs_ready)
		begin
			local_bb4_ld__u29_NO_SHIFT_REG <= local_bb4_ld__u29_lsu_dataout;
			local_bb4_ld__u29_valid_out_NO_SHIFT_REG <= local_bb4_ld__u29_fu_valid_out;
		end
		else
		begin
			if (~(local_bb4_ld__u29_stall_in))
			begin
				local_bb4_ld__u29_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_339to339_bb4_ld__u28_valid_out;
wire rstag_339to339_bb4_ld__u28_stall_in;
wire rstag_339to339_bb4_ld__u28_inputs_ready;
wire rstag_339to339_bb4_ld__u28_stall_local;
 reg rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG;
wire rstag_339to339_bb4_ld__u28_combined_valid;
 reg [31:0] rstag_339to339_bb4_ld__u28_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_339to339_bb4_ld__u28;

assign rstag_339to339_bb4_ld__u28_inputs_ready = local_bb4_ld__u28_valid_out_NO_SHIFT_REG;
assign rstag_339to339_bb4_ld__u28 = (rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG ? rstag_339to339_bb4_ld__u28_staging_reg_NO_SHIFT_REG : local_bb4_ld__u28_NO_SHIFT_REG);
assign rstag_339to339_bb4_ld__u28_combined_valid = (rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG | rstag_339to339_bb4_ld__u28_inputs_ready);
assign rstag_339to339_bb4_ld__u28_valid_out = rstag_339to339_bb4_ld__u28_combined_valid;
assign rstag_339to339_bb4_ld__u28_stall_local = rstag_339to339_bb4_ld__u28_stall_in;
assign local_bb4_ld__u28_stall_in = (|rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_339to339_bb4_ld__u28_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_339to339_bb4_ld__u28_stall_local)
		begin
			if (~(rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG))
			begin
				rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG <= rstag_339to339_bb4_ld__u28_inputs_ready;
			end
		end
		else
		begin
			rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_339to339_bb4_ld__u28_staging_valid_NO_SHIFT_REG))
		begin
			rstag_339to339_bb4_ld__u28_staging_reg_NO_SHIFT_REG <= local_bb4_ld__u28_NO_SHIFT_REG;
		end
	end
end


// This section implements a staging register.
// 
wire rstag_339to339_bb4_ld__u29_valid_out;
wire rstag_339to339_bb4_ld__u29_stall_in;
wire rstag_339to339_bb4_ld__u29_inputs_ready;
wire rstag_339to339_bb4_ld__u29_stall_local;
 reg rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG;
wire rstag_339to339_bb4_ld__u29_combined_valid;
 reg [31:0] rstag_339to339_bb4_ld__u29_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_339to339_bb4_ld__u29;

assign rstag_339to339_bb4_ld__u29_inputs_ready = local_bb4_ld__u29_valid_out_NO_SHIFT_REG;
assign rstag_339to339_bb4_ld__u29 = (rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG ? rstag_339to339_bb4_ld__u29_staging_reg_NO_SHIFT_REG : local_bb4_ld__u29_NO_SHIFT_REG);
assign rstag_339to339_bb4_ld__u29_combined_valid = (rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG | rstag_339to339_bb4_ld__u29_inputs_ready);
assign rstag_339to339_bb4_ld__u29_valid_out = rstag_339to339_bb4_ld__u29_combined_valid;
assign rstag_339to339_bb4_ld__u29_stall_local = rstag_339to339_bb4_ld__u29_stall_in;
assign local_bb4_ld__u29_stall_in = (|rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_339to339_bb4_ld__u29_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_339to339_bb4_ld__u29_stall_local)
		begin
			if (~(rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG))
			begin
				rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG <= rstag_339to339_bb4_ld__u29_inputs_ready;
			end
		end
		else
		begin
			rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_339to339_bb4_ld__u29_staging_valid_NO_SHIFT_REG))
		begin
			rstag_339to339_bb4_ld__u29_staging_reg_NO_SHIFT_REG <= local_bb4_ld__u29_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni2_stall_local;
wire [255:0] local_bb4_c1_eni2;

assign local_bb4_c1_eni2[63:0] = local_bb4_c1_eni1[63:0];
assign local_bb4_c1_eni2[95:64] = rstag_339to339_bb4_ld__u29;
assign local_bb4_c1_eni2[255:96] = local_bb4_c1_eni1[255:96];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni3_stall_local;
wire [255:0] local_bb4_c1_eni3;

assign local_bb4_c1_eni3[95:0] = local_bb4_c1_eni2[95:0];
assign local_bb4_c1_eni3[127:96] = rstag_339to339_bb4_ld__u28;
assign local_bb4_c1_eni3[255:128] = local_bb4_c1_eni2[255:128];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni4_stall_local;
wire [255:0] local_bb4_c1_eni4;

assign local_bb4_c1_eni4[127:0] = local_bb4_c1_eni3[127:0];
assign local_bb4_c1_eni4[159:128] = rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG[31:0];
assign local_bb4_c1_eni4[255:160] = local_bb4_c1_eni3[255:160];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni5_stall_local;
wire [255:0] local_bb4_c1_eni5;

assign local_bb4_c1_eni5[159:0] = local_bb4_c1_eni4[159:0];
assign local_bb4_c1_eni5[160] = rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG[32];
assign local_bb4_c1_eni5[255:161] = local_bb4_c1_eni4[255:161];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni6_stall_local;
wire [255:0] local_bb4_c1_eni6;

assign local_bb4_c1_eni6[191:0] = local_bb4_c1_eni5[191:0];
assign local_bb4_c1_eni6[223:192] = rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG[64:33];
assign local_bb4_c1_eni6[255:224] = local_bb4_c1_eni5[255:224];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni7_stall_local;
wire [255:0] local_bb4_c1_eni7;

assign local_bb4_c1_eni7[223:0] = local_bb4_c1_eni6[223:0];
assign local_bb4_c1_eni7[224] = rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG[65];
assign local_bb4_c1_eni7[255:225] = local_bb4_c1_eni6[255:225];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni8_valid_out;
wire local_bb4_c1_eni8_stall_in;
wire local_bb4_c0_exe5_valid_out_1;
wire local_bb4_c0_exe5_stall_in_1;
wire local_bb4_c1_eni8_inputs_ready;
wire local_bb4_c1_eni8_stall_local;
wire [255:0] local_bb4_c1_eni8;

assign local_bb4_c1_eni8_inputs_ready = (rcnode_338to339_rc0_t_313_0_valid_out_0_NO_SHIFT_REG & rcnode_338to339_rc0_t_313_0_valid_out_1_NO_SHIFT_REG & rcnode_338to339_rc0_t_313_0_valid_out_3_NO_SHIFT_REG & rcnode_338to339_rc0_t_313_0_valid_out_4_NO_SHIFT_REG & rcnode_338to339_rc0_t_313_0_valid_out_5_NO_SHIFT_REG & rstag_339to339_bb4_ld__u29_valid_out & rstag_339to339_bb4_ld__u28_valid_out & rnode_338to339_bb4_c0_exit214_c0_exi7_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_c1_eni8[231:0] = local_bb4_c1_eni7[231:0];
assign local_bb4_c1_eni8[232] = local_bb4_c0_exe5;
assign local_bb4_c1_eni8[255:233] = local_bb4_c1_eni7[255:233];
assign local_bb4_c1_eni8_stall_local = (local_bb4_c1_eni8_stall_in | local_bb4_c0_exe5_stall_in_1);
assign local_bb4_c1_eni8_valid_out = local_bb4_c1_eni8_inputs_ready;
assign local_bb4_c0_exe5_valid_out_1 = local_bb4_c1_eni8_inputs_ready;
assign rcnode_338to339_rc0_t_313_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));
assign rcnode_338to339_rc0_t_313_0_stall_in_1_NO_SHIFT_REG = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));
assign rcnode_338to339_rc0_t_313_0_stall_in_3_NO_SHIFT_REG = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));
assign rcnode_338to339_rc0_t_313_0_stall_in_4_NO_SHIFT_REG = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));
assign rcnode_338to339_rc0_t_313_0_stall_in_5_NO_SHIFT_REG = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));
assign rstag_339to339_bb4_ld__u29_stall_in = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));
assign rstag_339to339_bb4_ld__u28_stall_in = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));
assign rnode_338to339_bb4_c0_exit214_c0_exi7_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c1_eni8_stall_local | ~(local_bb4_c1_eni8_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb4_c1_enter_c1_eni8_inputs_ready;
 reg local_bb4_c1_enter_c1_eni8_valid_out_0_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_0;
 reg local_bb4_c1_enter_c1_eni8_valid_out_1_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_1;
 reg local_bb4_c1_enter_c1_eni8_valid_out_2_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_2;
 reg local_bb4_c1_enter_c1_eni8_valid_out_3_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_3;
 reg local_bb4_c1_enter_c1_eni8_valid_out_4_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_4;
 reg local_bb4_c1_enter_c1_eni8_valid_out_5_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_5;
 reg local_bb4_c1_enter_c1_eni8_valid_out_6_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_6;
 reg local_bb4_c1_enter_c1_eni8_valid_out_7_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_7;
 reg local_bb4_c1_enter_c1_eni8_valid_out_8_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_stall_in_8;
wire local_bb4_c1_enter_c1_eni8_output_regs_ready;
 reg [255:0] local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni8_input_accepted;
 reg local_bb4_c1_enter_c1_eni8_valid_bit_NO_SHIFT_REG;
wire local_bb4_c1_exit_c1_exi2_entry_stall;
wire local_bb4_c1_exit_c1_exi2_output_regs_ready;
wire [64:0] local_bb4_c1_exit_c1_exi2_valid_bits;
wire local_bb4_c1_exit_c1_exi2_valid_in;
wire local_bb4_c1_exit_c1_exi2_phases;
wire local_bb4_c1_enter_c1_eni8_inc_pipelined_thread;
wire local_bb4_c1_enter_c1_eni8_dec_pipelined_thread;
wire local_bb4_c1_enter_c1_eni8_causedstall;

assign local_bb4_c1_enter_c1_eni8_inputs_ready = (local_bb4_c1_eni8_valid_out & local_bb4_c0_exe5_valid_out_1 & rcnode_338to339_rc0_t_313_0_valid_out_2_NO_SHIFT_REG);
assign local_bb4_c1_enter_c1_eni8_output_regs_ready = 1'b1;
assign local_bb4_c1_enter_c1_eni8_input_accepted = (local_bb4_c1_enter_c1_eni8_inputs_ready && !(local_bb4_c1_exit_c1_exi2_entry_stall));
assign local_bb4_c1_enter_c1_eni8_inc_pipelined_thread = rcnode_338to339_rc0_t_313_0_NO_SHIFT_REG[32];
assign local_bb4_c1_enter_c1_eni8_dec_pipelined_thread = ~(local_bb4_c0_exe5);
assign local_bb4_c1_eni8_stall_in = ((~(local_bb4_c1_enter_c1_eni8_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign local_bb4_c0_exe5_stall_in_1 = ((~(local_bb4_c1_enter_c1_eni8_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign rcnode_338to339_rc0_t_313_0_stall_in_2_NO_SHIFT_REG = ((~(local_bb4_c1_enter_c1_eni8_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign local_bb4_c1_enter_c1_eni8_causedstall = (1'b1 && ((~(local_bb4_c1_enter_c1_eni8_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_enter_c1_eni8_valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb4_c1_enter_c1_eni8_valid_bit_NO_SHIFT_REG <= local_bb4_c1_enter_c1_eni8_input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG <= 'x;
		local_bb4_c1_enter_c1_eni8_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_7_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni8_valid_out_8_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c1_enter_c1_eni8_output_regs_ready)
		begin
			local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG <= local_bb4_c1_eni8;
			local_bb4_c1_enter_c1_eni8_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_6_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_7_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni8_valid_out_8_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_0))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_1))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_2))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_3))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_4))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_5))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_6))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_7))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni8_stall_in_8))
			begin
				local_bb4_c1_enter_c1_eni8_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene1_stall_local;
wire [31:0] local_bb4_c1_ene1;

assign local_bb4_c1_ene1 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene2_stall_local;
wire [31:0] local_bb4_c1_ene2;

assign local_bb4_c1_ene2 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[95:64];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene3_stall_local;
wire [31:0] local_bb4_c1_ene3;

assign local_bb4_c1_ene3 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[127:96];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene4_valid_out;
wire local_bb4_c1_ene4_stall_in;
wire local_bb4_c1_ene4_inputs_ready;
wire local_bb4_c1_ene4_stall_local;
wire [31:0] local_bb4_c1_ene4;

assign local_bb4_c1_ene4_inputs_ready = local_bb4_c1_enter_c1_eni8_valid_out_3_NO_SHIFT_REG;
assign local_bb4_c1_ene4 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[159:128];
assign local_bb4_c1_ene4_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni8_stall_in_3 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene5_stall_local;
wire local_bb4_c1_ene5;

assign local_bb4_c1_ene5 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[160];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene6_valid_out;
wire local_bb4_c1_ene6_stall_in;
wire local_bb4_c1_ene6_inputs_ready;
wire local_bb4_c1_ene6_stall_local;
wire [31:0] local_bb4_c1_ene6;

assign local_bb4_c1_ene6_inputs_ready = local_bb4_c1_enter_c1_eni8_valid_out_5_NO_SHIFT_REG;
assign local_bb4_c1_ene6 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[223:192];
assign local_bb4_c1_ene6_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni8_stall_in_5 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene7_valid_out;
wire local_bb4_c1_ene7_stall_in;
wire local_bb4_c1_ene7_inputs_ready;
wire local_bb4_c1_ene7_stall_local;
wire local_bb4_c1_ene7;

assign local_bb4_c1_ene7_inputs_ready = local_bb4_c1_enter_c1_eni8_valid_out_6_NO_SHIFT_REG;
assign local_bb4_c1_ene7 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[224];
assign local_bb4_c1_ene7_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni8_stall_in_6 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene8_valid_out;
wire local_bb4_c1_ene8_stall_in;
wire local_bb4_c1_ene8_inputs_ready;
wire local_bb4_c1_ene8_stall_local;
wire local_bb4_c1_ene8;

assign local_bb4_c1_ene8_inputs_ready = local_bb4_c1_enter_c1_eni8_valid_out_7_NO_SHIFT_REG;
assign local_bb4_c1_ene8 = local_bb4_c1_enter_c1_eni8_NO_SHIFT_REG[232];
assign local_bb4_c1_ene8_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni8_stall_in_7 = 1'b0;

// This section implements an unregistered operation.
// 
wire SFC_3_VALID_340_340_0_valid_out;
wire SFC_3_VALID_340_340_0_stall_in;
wire SFC_3_VALID_340_340_0_inputs_ready;
wire SFC_3_VALID_340_340_0_stall_local;
wire SFC_3_VALID_340_340_0;

assign SFC_3_VALID_340_340_0_inputs_ready = local_bb4_c1_enter_c1_eni8_valid_out_8_NO_SHIFT_REG;
assign SFC_3_VALID_340_340_0 = local_bb4_c1_enter_c1_eni8_valid_bit_NO_SHIFT_REG;
assign SFC_3_VALID_340_340_0_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni8_stall_in_8 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u30_stall_local;
wire [31:0] local_bb4_var__u30;

assign local_bb4_var__u30 = local_bb4_c1_ene1;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u31_stall_local;
wire [31:0] local_bb4_var__u31;

assign local_bb4_var__u31 = local_bb4_c1_ene2;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u32_stall_local;
wire [31:0] local_bb4_var__u32;

assign local_bb4_var__u32 = local_bb4_c1_ene3;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene4_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_c1_ene4_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene4_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene4_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene4_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_c1_ene4_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_c1_ene4_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_c1_ene4_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_c1_ene4_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_c1_ene4_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene4),
	.data_out(rnode_340to341_bb4_c1_ene4_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_c1_ene4_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_c1_ene4_0_reg_341_fifo.DATA_WIDTH = 32;
defparam rnode_340to341_bb4_c1_ene4_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_c1_ene4_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_c1_ene4_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene4_stall_in = 1'b0;
assign rnode_340to341_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_340to341_bb4_c1_ene4_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_c1_ene4_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_f_8_stall_local;
wire [31:0] local_bb4__acl_ffwd_dest_f_8;

assign local_bb4__acl_ffwd_dest_f_8 = ffwd_8_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene6_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_c1_ene6_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene6_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene6_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene6_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_c1_ene6_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_c1_ene6_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_c1_ene6_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_c1_ene6_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_c1_ene6_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene6),
	.data_out(rnode_340to341_bb4_c1_ene6_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_c1_ene6_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_c1_ene6_0_reg_341_fifo.DATA_WIDTH = 32;
defparam rnode_340to341_bb4_c1_ene6_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_c1_ene6_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_c1_ene6_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene6_stall_in = 1'b0;
assign rnode_340to341_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_340to341_bb4_c1_ene6_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_c1_ene6_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene7_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene7_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene7_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene7_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene7_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene7_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_c1_ene7_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_c1_ene7_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_c1_ene7_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_c1_ene7_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_c1_ene7_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene7),
	.data_out(rnode_340to341_bb4_c1_ene7_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_c1_ene7_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_c1_ene7_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb4_c1_ene7_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_c1_ene7_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_c1_ene7_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene7_stall_in = 1'b0;
assign rnode_340to341_bb4_c1_ene7_0_NO_SHIFT_REG = rnode_340to341_bb4_c1_ene7_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_c1_ene7_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene8_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene8_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene8_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene8_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene8_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene8_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_c1_ene8_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_c1_ene8_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_c1_ene8_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_c1_ene8_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_c1_ene8_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene8),
	.data_out(rnode_340to341_bb4_c1_ene8_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_c1_ene8_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_c1_ene8_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb4_c1_ene8_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_c1_ene8_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_c1_ene8_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene8_stall_in = 1'b0;
assign rnode_340to341_bb4_c1_ene8_0_NO_SHIFT_REG = rnode_340to341_bb4_c1_ene8_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_c1_ene8_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_340_341_0_inputs_ready;
 reg SFC_3_VALID_340_341_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_340_341_0_stall_in;
wire SFC_3_VALID_340_341_0_output_regs_ready;
 reg SFC_3_VALID_340_341_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_340_341_0_causedstall;

assign SFC_3_VALID_340_341_0_inputs_ready = 1'b1;
assign SFC_3_VALID_340_341_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_340_340_0_stall_in = 1'b0;
assign SFC_3_VALID_340_341_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_340_341_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_340_341_0_output_regs_ready)
		begin
			SFC_3_VALID_340_341_0_NO_SHIFT_REG <= SFC_3_VALID_340_340_0;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and2_i499_stall_local;
wire [31:0] local_bb4_and2_i499;

assign local_bb4_and2_i499 = (local_bb4_var__u30 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i504_stall_local;
wire [31:0] local_bb4_and12_i504;

assign local_bb4_and12_i504 = (local_bb4_var__u30 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i312_stall_local;
wire [31:0] local_bb4_shr_i312;

assign local_bb4_shr_i312 = (local_bb4_var__u31 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and5_i318_stall_local;
wire [31:0] local_bb4_and5_i318;

assign local_bb4_and5_i318 = (local_bb4_var__u31 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i314_stall_local;
wire [31:0] local_bb4_shr2_i314;

assign local_bb4_shr2_i314 = (local_bb4_var__u32 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i316_stall_local;
wire [31:0] local_bb4_xor_i316;

assign local_bb4_xor_i316 = (local_bb4_var__u32 ^ local_bb4_var__u31);

// This section implements an unregistered operation.
// 
wire local_bb4_and6_i319_stall_local;
wire [31:0] local_bb4_and6_i319;

assign local_bb4_and6_i319 = (local_bb4_var__u32 & 32'h7FFFFF);

// Register node:
//  * latency = 51
//  * capacity = 51
 logic rnode_341to392_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to392_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_341to392_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_341to392_bb4_c1_ene4_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to392_bb4_c1_ene4_0_reg_392_NO_SHIFT_REG;
 logic rnode_341to392_bb4_c1_ene4_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_341to392_bb4_c1_ene4_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_341to392_bb4_c1_ene4_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_341to392_bb4_c1_ene4_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to392_bb4_c1_ene4_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to392_bb4_c1_ene4_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_341to392_bb4_c1_ene4_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_341to392_bb4_c1_ene4_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_341to392_bb4_c1_ene4_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_341to392_bb4_c1_ene4_0_reg_392_fifo.DEPTH = 51;
defparam rnode_341to392_bb4_c1_ene4_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_341to392_bb4_c1_ene4_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to392_bb4_c1_ene4_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_341to392_bb4_c1_ene4_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to392_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_341to392_bb4_c1_ene4_0_reg_392_NO_SHIFT_REG;
assign rnode_341to392_bb4_c1_ene4_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_341to392_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u33_stall_local;
wire [31:0] local_bb4_var__u33;

assign local_bb4_var__u33 = local_bb4__acl_ffwd_dest_f_8;

// Register node:
//  * latency = 46
//  * capacity = 46
 logic rnode_341to387_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_341to387_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene6_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to387_bb4_c1_ene6_0_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene6_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene6_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene6_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_341to387_bb4_c1_ene6_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to387_bb4_c1_ene6_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to387_bb4_c1_ene6_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_341to387_bb4_c1_ene6_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_341to387_bb4_c1_ene6_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_341to387_bb4_c1_ene6_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_341to387_bb4_c1_ene6_0_reg_387_fifo.DEPTH = 46;
defparam rnode_341to387_bb4_c1_ene6_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_341to387_bb4_c1_ene6_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to387_bb4_c1_ene6_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_341to387_bb4_c1_ene6_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to387_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_341to387_bb4_c1_ene6_0_reg_387_NO_SHIFT_REG;
assign rnode_341to387_bb4_c1_ene6_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_341to387_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 54
//  * capacity = 54
 logic rnode_341to395_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to395_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to395_bb4_c1_ene7_0_NO_SHIFT_REG;
 logic rnode_341to395_bb4_c1_ene7_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to395_bb4_c1_ene7_0_reg_395_NO_SHIFT_REG;
 logic rnode_341to395_bb4_c1_ene7_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_341to395_bb4_c1_ene7_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_341to395_bb4_c1_ene7_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_341to395_bb4_c1_ene7_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to395_bb4_c1_ene7_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to395_bb4_c1_ene7_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_341to395_bb4_c1_ene7_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_341to395_bb4_c1_ene7_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_c1_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_341to395_bb4_c1_ene7_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_341to395_bb4_c1_ene7_0_reg_395_fifo.DEPTH = 54;
defparam rnode_341to395_bb4_c1_ene7_0_reg_395_fifo.DATA_WIDTH = 1;
defparam rnode_341to395_bb4_c1_ene7_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to395_bb4_c1_ene7_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_341to395_bb4_c1_ene7_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to395_bb4_c1_ene7_0_NO_SHIFT_REG = rnode_341to395_bb4_c1_ene7_0_reg_395_NO_SHIFT_REG;
assign rnode_341to395_bb4_c1_ene7_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_341to395_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 55
//  * capacity = 55
 logic rnode_341to396_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to396_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to396_bb4_c1_ene8_0_NO_SHIFT_REG;
 logic rnode_341to396_bb4_c1_ene8_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to396_bb4_c1_ene8_0_reg_396_NO_SHIFT_REG;
 logic rnode_341to396_bb4_c1_ene8_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_341to396_bb4_c1_ene8_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_341to396_bb4_c1_ene8_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_341to396_bb4_c1_ene8_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to396_bb4_c1_ene8_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to396_bb4_c1_ene8_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_341to396_bb4_c1_ene8_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_341to396_bb4_c1_ene8_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_c1_ene8_0_NO_SHIFT_REG),
	.data_out(rnode_341to396_bb4_c1_ene8_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_341to396_bb4_c1_ene8_0_reg_396_fifo.DEPTH = 55;
defparam rnode_341to396_bb4_c1_ene8_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_341to396_bb4_c1_ene8_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to396_bb4_c1_ene8_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_341to396_bb4_c1_ene8_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to396_bb4_c1_ene8_0_NO_SHIFT_REG = rnode_341to396_bb4_c1_ene8_0_reg_396_NO_SHIFT_REG;
assign rnode_341to396_bb4_c1_ene8_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_341to396_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_341_342_0_inputs_ready;
 reg SFC_3_VALID_341_342_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_341_342_0_stall_in;
wire SFC_3_VALID_341_342_0_output_regs_ready;
 reg SFC_3_VALID_341_342_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_341_342_0_causedstall;

assign SFC_3_VALID_341_342_0_inputs_ready = 1'b1;
assign SFC_3_VALID_341_342_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_340_341_0_stall_in = 1'b0;
assign SFC_3_VALID_341_342_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_341_342_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_341_342_0_output_regs_ready)
		begin
			SFC_3_VALID_341_342_0_NO_SHIFT_REG <= SFC_3_VALID_340_341_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i500_stall_local;
wire [31:0] local_bb4_shr3_i500;

assign local_bb4_shr3_i500 = ((local_bb4_and2_i499 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i313_stall_local;
wire [31:0] local_bb4_and_i313;

assign local_bb4_and_i313 = ((local_bb4_shr_i312 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i324_stall_local;
wire local_bb4_lnot14_i324;

assign local_bb4_lnot14_i324 = ((local_bb4_and5_i318 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i346_stall_local;
wire [31:0] local_bb4_or_i346;

assign local_bb4_or_i346 = ((local_bb4_and5_i318 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and3_i315_stall_local;
wire [31:0] local_bb4_and3_i315;

assign local_bb4_and3_i315 = ((local_bb4_shr2_i314 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_i325_stall_local;
wire local_bb4_lnot17_i325;

assign local_bb4_lnot17_i325 = ((local_bb4_and6_i319 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or47_i347_stall_local;
wire [31:0] local_bb4_or47_i347;

assign local_bb4_or47_i347 = ((local_bb4_and6_i319 & 32'h7FFFFF) | 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene4_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_c1_ene4_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene4_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene4_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene4_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_c1_ene4_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_c1_ene4_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_c1_ene4_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_c1_ene4_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_c1_ene4_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_341to392_bb4_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb4_c1_ene4_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_c1_ene4_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_c1_ene4_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_392to393_bb4_c1_ene4_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_c1_ene4_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_c1_ene4_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to392_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_392to393_bb4_c1_ene4_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_c1_ene4_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i496_stall_local;
wire [31:0] local_bb4_xor_i496;

assign local_bb4_xor_i496 = (local_bb4_var__u33 ^ 32'h80000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene6_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_c1_ene6_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene6_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene6_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene6_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_c1_ene6_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_c1_ene6_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_c1_ene6_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_c1_ene6_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_c1_ene6_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_341to387_bb4_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb4_c1_ene6_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_c1_ene6_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_c1_ene6_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb4_c1_ene6_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_c1_ene6_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_c1_ene6_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to387_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_387to388_bb4_c1_ene6_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_c1_ene6_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_c1_ene7_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_valid_out_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_stall_in_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_c1_ene7_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_c1_ene7_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_c1_ene7_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_c1_ene7_0_stall_in_0_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_c1_ene7_0_valid_out_0_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_c1_ene7_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(rnode_341to395_bb4_c1_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_395to396_bb4_c1_ene7_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_c1_ene7_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_c1_ene7_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_395to396_bb4_c1_ene7_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_c1_ene7_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_c1_ene7_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to395_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_c1_ene7_0_stall_in_0_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_c1_ene7_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_c1_ene7_0_NO_SHIFT_REG = rnode_395to396_bb4_c1_ene7_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_c1_ene7_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_c1_ene7_1_NO_SHIFT_REG = rnode_395to396_bb4_c1_ene7_0_reg_396_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_c1_ene8_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_valid_out_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_stall_in_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene8_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_c1_ene8_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_c1_ene8_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_c1_ene8_0_stall_in_0_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_c1_ene8_0_valid_out_0_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_c1_ene8_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(rnode_341to396_bb4_c1_ene8_0_NO_SHIFT_REG),
	.data_out(rnode_396to397_bb4_c1_ene8_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_c1_ene8_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_c1_ene8_0_reg_397_fifo.DATA_WIDTH = 1;
defparam rnode_396to397_bb4_c1_ene8_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_c1_ene8_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_c1_ene8_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to396_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_c1_ene8_0_stall_in_0_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_c1_ene8_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_c1_ene8_0_NO_SHIFT_REG = rnode_396to397_bb4_c1_ene8_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_c1_ene8_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_c1_ene8_1_NO_SHIFT_REG = rnode_396to397_bb4_c1_ene8_0_reg_397_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_342_343_0_inputs_ready;
 reg SFC_3_VALID_342_343_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_342_343_0_stall_in;
wire SFC_3_VALID_342_343_0_output_regs_ready;
 reg SFC_3_VALID_342_343_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_342_343_0_causedstall;

assign SFC_3_VALID_342_343_0_inputs_ready = 1'b1;
assign SFC_3_VALID_342_343_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_341_342_0_stall_in = 1'b0;
assign SFC_3_VALID_342_343_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_342_343_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_342_343_0_output_regs_ready)
		begin
			SFC_3_VALID_342_343_0_NO_SHIFT_REG <= SFC_3_VALID_341_342_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i320_stall_local;
wire local_bb4_lnot_i320;

assign local_bb4_lnot_i320 = ((local_bb4_and_i313 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i322_stall_local;
wire local_bb4_cmp_i322;

assign local_bb4_cmp_i322 = ((local_bb4_and_i313 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u34_stall_local;
wire [31:0] local_bb4_var__u34;

assign local_bb4_var__u34 = ((local_bb4_and6_i319 & 32'h7FFFFF) | (local_bb4_and_i313 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_not_i343_stall_local;
wire local_bb4_lnot14_not_i343;

assign local_bb4_lnot14_not_i343 = (local_bb4_lnot14_i324 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_conv_i_i348_stall_local;
wire [63:0] local_bb4_conv_i_i348;

assign local_bb4_conv_i_i348[63:32] = 32'h0;
assign local_bb4_conv_i_i348[31:0] = ((local_bb4_or_i346 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot8_i321_stall_local;
wire local_bb4_lnot8_i321;

assign local_bb4_lnot8_i321 = ((local_bb4_and3_i315 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_i323_stall_local;
wire local_bb4_cmp11_i323;

assign local_bb4_cmp11_i323 = ((local_bb4_and3_i315 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u35_stall_local;
wire [31:0] local_bb4_var__u35;

assign local_bb4_var__u35 = ((local_bb4_and3_i315 & 32'hFF) | (local_bb4_and6_i319 & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i357_stall_local;
wire [31:0] local_bb4_add_i357;

assign local_bb4_add_i357 = ((local_bb4_and3_i315 & 32'hFF) + (local_bb4_and_i313 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_not_i329_stall_local;
wire local_bb4_lnot17_not_i329;

assign local_bb4_lnot17_not_i329 = (local_bb4_lnot17_i325 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_conv1_i_i349_stall_local;
wire [63:0] local_bb4_conv1_i_i349;

assign local_bb4_conv1_i_i349[63:32] = 32'h0;
assign local_bb4_conv1_i_i349[31:0] = ((local_bb4_or47_i347 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i497_stall_local;
wire [31:0] local_bb4_and_i497;

assign local_bb4_and_i497 = (local_bb4_xor_i496 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i503_stall_local;
wire [31:0] local_bb4_and10_i503;

assign local_bb4_and10_i503 = (local_bb4_xor_i496 & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene7_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene7_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene7_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene7_0_valid_out_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene7_0_stall_in_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_c1_ene7_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_c1_ene7_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_c1_ene7_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_c1_ene7_0_stall_in_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_c1_ene7_0_valid_out_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_c1_ene7_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(rnode_395to396_bb4_c1_ene7_1_NO_SHIFT_REG),
	.data_out(rnode_396to397_bb4_c1_ene7_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_c1_ene7_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_c1_ene7_0_reg_397_fifo.DATA_WIDTH = 1;
defparam rnode_396to397_bb4_c1_ene7_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_c1_ene7_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_c1_ene7_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_c1_ene7_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_c1_ene7_0_NO_SHIFT_REG = rnode_396to397_bb4_c1_ene7_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_c1_ene7_0_stall_in_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_397to398_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to398_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG;
 logic rnode_397to398_bb4_c1_ene8_0_NO_SHIFT_REG;
 logic rnode_397to398_bb4_c1_ene8_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic rnode_397to398_bb4_c1_ene8_0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_c1_ene8_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_c1_ene8_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_c1_ene8_0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_397to398_bb4_c1_ene8_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to398_bb4_c1_ene8_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to398_bb4_c1_ene8_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_397to398_bb4_c1_ene8_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_397to398_bb4_c1_ene8_0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(rnode_396to397_bb4_c1_ene8_1_NO_SHIFT_REG),
	.data_out(rnode_397to398_bb4_c1_ene8_0_reg_398_NO_SHIFT_REG)
);

defparam rnode_397to398_bb4_c1_ene8_0_reg_398_fifo.DEPTH = 1;
defparam rnode_397to398_bb4_c1_ene8_0_reg_398_fifo.DATA_WIDTH = 1;
defparam rnode_397to398_bb4_c1_ene8_0_reg_398_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to398_bb4_c1_ene8_0_reg_398_fifo.IMPL = "shift_reg";

assign rnode_397to398_bb4_c1_ene8_0_reg_398_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_c1_ene8_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_397to398_bb4_c1_ene8_0_NO_SHIFT_REG = rnode_397to398_bb4_c1_ene8_0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb4_c1_ene8_0_stall_in_reg_398_NO_SHIFT_REG = 1'b0;
assign rnode_397to398_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_343_344_0_inputs_ready;
 reg SFC_3_VALID_343_344_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_343_344_0_stall_in;
wire SFC_3_VALID_343_344_0_output_regs_ready;
 reg SFC_3_VALID_343_344_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_343_344_0_causedstall;

assign SFC_3_VALID_343_344_0_inputs_ready = 1'b1;
assign SFC_3_VALID_343_344_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_342_343_0_stall_in = 1'b0;
assign SFC_3_VALID_343_344_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_343_344_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_343_344_0_output_regs_ready)
		begin
			SFC_3_VALID_343_344_0_NO_SHIFT_REG <= SFC_3_VALID_342_343_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u36_stall_local;
wire local_bb4_var__u36;

assign local_bb4_var__u36 = ((local_bb4_var__u34 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i344_stall_local;
wire local_bb4__28_i344;

assign local_bb4__28_i344 = (local_bb4_cmp_i322 & local_bb4_lnot14_not_i343);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i375_stall_local;
wire local_bb4_reduction_0_i375;

assign local_bb4_reduction_0_i375 = (local_bb4_lnot_i320 | local_bb4_lnot8_i321);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge8_demorgan_i326_stall_local;
wire local_bb4_brmerge8_demorgan_i326;

assign local_bb4_brmerge8_demorgan_i326 = (local_bb4_cmp11_i323 & local_bb4_lnot17_i325);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_not_i330_stall_local;
wire local_bb4_cmp11_not_i330;

assign local_bb4_cmp11_not_i330 = (local_bb4_cmp11_i323 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u37_stall_local;
wire local_bb4_var__u37;

assign local_bb4_var__u37 = (local_bb4_cmp_i322 | local_bb4_cmp11_i323);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u38_stall_local;
wire local_bb4_var__u38;

assign local_bb4_var__u38 = ((local_bb4_var__u35 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i498_stall_local;
wire [31:0] local_bb4_shr_i498;

assign local_bb4_shr_i498 = ((local_bb4_and_i497 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i505_stall_local;
wire local_bb4_cmp13_i505;

assign local_bb4_cmp13_i505 = ((local_bb4_and10_i503 & 32'hFFFF) > (local_bb4_and12_i504 & 32'hFFFF));

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_397to400_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to400_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_397to400_bb4_c1_ene7_0_NO_SHIFT_REG;
 logic rnode_397to400_bb4_c1_ene7_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic rnode_397to400_bb4_c1_ene7_0_reg_400_NO_SHIFT_REG;
 logic rnode_397to400_bb4_c1_ene7_0_valid_out_reg_400_NO_SHIFT_REG;
 logic rnode_397to400_bb4_c1_ene7_0_stall_in_reg_400_NO_SHIFT_REG;
 logic rnode_397to400_bb4_c1_ene7_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_397to400_bb4_c1_ene7_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to400_bb4_c1_ene7_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to400_bb4_c1_ene7_0_stall_in_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_397to400_bb4_c1_ene7_0_valid_out_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_397to400_bb4_c1_ene7_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in(rnode_396to397_bb4_c1_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_397to400_bb4_c1_ene7_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_397to400_bb4_c1_ene7_0_reg_400_fifo.DEPTH = 3;
defparam rnode_397to400_bb4_c1_ene7_0_reg_400_fifo.DATA_WIDTH = 1;
defparam rnode_397to400_bb4_c1_ene7_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to400_bb4_c1_ene7_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_397to400_bb4_c1_ene7_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_397to400_bb4_c1_ene7_0_NO_SHIFT_REG = rnode_397to400_bb4_c1_ene7_0_reg_400_NO_SHIFT_REG;
assign rnode_397to400_bb4_c1_ene7_0_stall_in_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_397to400_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_398to401_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_398to401_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG;
 logic rnode_398to401_bb4_c1_ene8_0_NO_SHIFT_REG;
 logic rnode_398to401_bb4_c1_ene8_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic rnode_398to401_bb4_c1_ene8_0_reg_401_NO_SHIFT_REG;
 logic rnode_398to401_bb4_c1_ene8_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_398to401_bb4_c1_ene8_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_398to401_bb4_c1_ene8_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_398to401_bb4_c1_ene8_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to401_bb4_c1_ene8_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to401_bb4_c1_ene8_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_398to401_bb4_c1_ene8_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_398to401_bb4_c1_ene8_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(rnode_397to398_bb4_c1_ene8_0_NO_SHIFT_REG),
	.data_out(rnode_398to401_bb4_c1_ene8_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_398to401_bb4_c1_ene8_0_reg_401_fifo.DEPTH = 3;
defparam rnode_398to401_bb4_c1_ene8_0_reg_401_fifo.DATA_WIDTH = 1;
defparam rnode_398to401_bb4_c1_ene8_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to401_bb4_c1_ene8_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_398to401_bb4_c1_ene8_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_398to401_bb4_c1_ene8_0_NO_SHIFT_REG = rnode_398to401_bb4_c1_ene8_0_reg_401_NO_SHIFT_REG;
assign rnode_398to401_bb4_c1_ene8_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_398to401_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_344_345_0_inputs_ready;
 reg SFC_3_VALID_344_345_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_344_345_0_stall_in;
wire SFC_3_VALID_344_345_0_output_regs_ready;
 reg SFC_3_VALID_344_345_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_344_345_0_causedstall;

assign SFC_3_VALID_344_345_0_inputs_ready = 1'b1;
assign SFC_3_VALID_344_345_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_343_344_0_stall_in = 1'b0;
assign SFC_3_VALID_344_345_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_344_345_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_344_345_0_output_regs_ready)
		begin
			SFC_3_VALID_344_345_0_NO_SHIFT_REG <= SFC_3_VALID_343_344_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_brmerge10_demorgan_i327_stall_local;
wire local_bb4_brmerge10_demorgan_i327;

assign local_bb4_brmerge10_demorgan_i327 = (local_bb4_brmerge8_demorgan_i326 & local_bb4_lnot_i320);

// This section implements an unregistered operation.
// 
wire local_bb4__mux9_mux_i328_stall_local;
wire local_bb4__mux9_mux_i328;

assign local_bb4__mux9_mux_i328 = (local_bb4_brmerge8_demorgan_i326 ^ local_bb4_cmp11_i323);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge3_i331_stall_local;
wire local_bb4_brmerge3_i331;

assign local_bb4_brmerge3_i331 = (local_bb4_var__u38 | local_bb4_cmp11_not_i330);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_i333_stall_local;
wire local_bb4__mux_mux_i333;

assign local_bb4__mux_mux_i333 = (local_bb4_var__u38 | local_bb4_cmp11_i323);

// This section implements an unregistered operation.
// 
wire local_bb4__not_i335_stall_local;
wire local_bb4__not_i335;

assign local_bb4__not_i335 = (local_bb4_var__u38 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i501_stall_local;
wire local_bb4_cmp_i501;

assign local_bb4_cmp_i501 = ((local_bb4_shr_i498 & 32'h7FFF) > (local_bb4_shr3_i500 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i502_stall_local;
wire local_bb4_cmp8_i502;

assign local_bb4_cmp8_i502 = ((local_bb4_shr_i498 & 32'h7FFF) == (local_bb4_shr3_i500 & 32'h7FFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_400to401_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_400to401_bb4_c1_ene7_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_c1_ene7_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic rnode_400to401_bb4_c1_ene7_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_c1_ene7_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_c1_ene7_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_c1_ene7_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4_c1_ene7_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4_c1_ene7_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4_c1_ene7_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4_c1_ene7_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4_c1_ene7_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(rnode_397to400_bb4_c1_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_400to401_bb4_c1_ene7_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4_c1_ene7_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4_c1_ene7_0_reg_401_fifo.DATA_WIDTH = 1;
defparam rnode_400to401_bb4_c1_ene7_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4_c1_ene7_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4_c1_ene7_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_397to400_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_c1_ene7_0_NO_SHIFT_REG = rnode_400to401_bb4_c1_ene7_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_c1_ene7_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_401to402_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_401to402_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG;
 logic rnode_401to402_bb4_c1_ene8_0_NO_SHIFT_REG;
 logic rnode_401to402_bb4_c1_ene8_0_reg_402_inputs_ready_NO_SHIFT_REG;
 logic rnode_401to402_bb4_c1_ene8_0_reg_402_NO_SHIFT_REG;
 logic rnode_401to402_bb4_c1_ene8_0_valid_out_reg_402_NO_SHIFT_REG;
 logic rnode_401to402_bb4_c1_ene8_0_stall_in_reg_402_NO_SHIFT_REG;
 logic rnode_401to402_bb4_c1_ene8_0_stall_out_reg_402_NO_SHIFT_REG;

acl_data_fifo rnode_401to402_bb4_c1_ene8_0_reg_402_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_401to402_bb4_c1_ene8_0_reg_402_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_401to402_bb4_c1_ene8_0_stall_in_reg_402_NO_SHIFT_REG),
	.valid_out(rnode_401to402_bb4_c1_ene8_0_valid_out_reg_402_NO_SHIFT_REG),
	.stall_out(rnode_401to402_bb4_c1_ene8_0_stall_out_reg_402_NO_SHIFT_REG),
	.data_in(rnode_398to401_bb4_c1_ene8_0_NO_SHIFT_REG),
	.data_out(rnode_401to402_bb4_c1_ene8_0_reg_402_NO_SHIFT_REG)
);

defparam rnode_401to402_bb4_c1_ene8_0_reg_402_fifo.DEPTH = 1;
defparam rnode_401to402_bb4_c1_ene8_0_reg_402_fifo.DATA_WIDTH = 1;
defparam rnode_401to402_bb4_c1_ene8_0_reg_402_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_401to402_bb4_c1_ene8_0_reg_402_fifo.IMPL = "shift_reg";

assign rnode_401to402_bb4_c1_ene8_0_reg_402_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_398to401_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_401to402_bb4_c1_ene8_0_NO_SHIFT_REG = rnode_401to402_bb4_c1_ene8_0_reg_402_NO_SHIFT_REG;
assign rnode_401to402_bb4_c1_ene8_0_stall_in_reg_402_NO_SHIFT_REG = 1'b0;
assign rnode_401to402_bb4_c1_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_345_346_0_inputs_ready;
 reg SFC_3_VALID_345_346_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_345_346_0_stall_in;
wire SFC_3_VALID_345_346_0_output_regs_ready;
 reg SFC_3_VALID_345_346_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_345_346_0_causedstall;

assign SFC_3_VALID_345_346_0_inputs_ready = 1'b1;
assign SFC_3_VALID_345_346_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_344_345_0_stall_in = 1'b0;
assign SFC_3_VALID_345_346_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_345_346_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_345_346_0_output_regs_ready)
		begin
			SFC_3_VALID_345_346_0_NO_SHIFT_REG <= SFC_3_VALID_344_345_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__26_demorgan_i341_stall_local;
wire local_bb4__26_demorgan_i341;

assign local_bb4__26_demorgan_i341 = (local_bb4_cmp_i322 | local_bb4_brmerge10_demorgan_i327);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge5_i332_stall_local;
wire local_bb4_brmerge5_i332;

assign local_bb4_brmerge5_i332 = (local_bb4_brmerge3_i331 | local_bb4_lnot17_not_i329);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i336_stall_local;
wire local_bb4_reduction_3_i336;

assign local_bb4_reduction_3_i336 = (local_bb4_cmp11_i323 & local_bb4__not_i335);

// This section implements an unregistered operation.
// 
wire local_bb4___i506_stall_local;
wire local_bb4___i506;

assign local_bb4___i506 = (local_bb4_cmp8_i502 & local_bb4_cmp13_i505);

// This section implements a registered operation.
// 
wire SFC_3_VALID_346_347_0_inputs_ready;
 reg SFC_3_VALID_346_347_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_346_347_0_stall_in;
wire SFC_3_VALID_346_347_0_output_regs_ready;
 reg SFC_3_VALID_346_347_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_346_347_0_causedstall;

assign SFC_3_VALID_346_347_0_inputs_ready = 1'b1;
assign SFC_3_VALID_346_347_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_345_346_0_stall_in = 1'b0;
assign SFC_3_VALID_346_347_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_346_347_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_346_347_0_output_regs_ready)
		begin
			SFC_3_VALID_346_347_0_NO_SHIFT_REG <= SFC_3_VALID_345_346_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_mux_i334_stall_local;
wire local_bb4__mux_mux_mux_i334;

assign local_bb4__mux_mux_mux_i334 = (local_bb4_brmerge5_i332 & local_bb4__mux_mux_i333);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i337_stall_local;
wire local_bb4_reduction_5_i337;

assign local_bb4_reduction_5_i337 = (local_bb4_lnot14_i324 & local_bb4_reduction_3_i336);

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene1_valid_out_1;
wire local_bb4_c1_ene1_stall_in_1;
wire local_bb4_var__u30_valid_out_2;
wire local_bb4_var__u30_stall_in_2;
wire local_bb4__21_i507_valid_out;
wire local_bb4__21_i507_stall_in;
wire local_bb4_c1_ene5_valid_out_1;
wire local_bb4_c1_ene5_stall_in_1;
wire local_bb4_xor_i496_valid_out_2;
wire local_bb4_xor_i496_stall_in_2;
wire local_bb4__21_i507_inputs_ready;
wire local_bb4__21_i507_stall_local;
wire local_bb4__21_i507;

assign local_bb4__21_i507_inputs_ready = (local_bb4_c1_enter_c1_eni8_valid_out_0_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni8_valid_out_4_NO_SHIFT_REG);
assign local_bb4__21_i507 = (local_bb4_cmp_i501 | local_bb4___i506);
assign local_bb4_c1_ene1_valid_out_1 = 1'b1;
assign local_bb4_var__u30_valid_out_2 = 1'b1;
assign local_bb4__21_i507_valid_out = 1'b1;
assign local_bb4_c1_ene5_valid_out_1 = 1'b1;
assign local_bb4_xor_i496_valid_out_2 = 1'b1;
assign local_bb4_c1_enter_c1_eni8_stall_in_0 = 1'b0;
assign local_bb4_c1_enter_c1_eni8_stall_in_4 = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_347_348_0_inputs_ready;
 reg SFC_3_VALID_347_348_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_347_348_0_stall_in;
wire SFC_3_VALID_347_348_0_output_regs_ready;
 reg SFC_3_VALID_347_348_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_347_348_0_causedstall;

assign SFC_3_VALID_347_348_0_inputs_ready = 1'b1;
assign SFC_3_VALID_347_348_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_346_347_0_stall_in = 1'b0;
assign SFC_3_VALID_347_348_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_347_348_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_347_348_0_output_regs_ready)
		begin
			SFC_3_VALID_347_348_0_NO_SHIFT_REG <= SFC_3_VALID_346_347_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i338_stall_local;
wire local_bb4_reduction_6_i338;

assign local_bb4_reduction_6_i338 = (local_bb4_var__u36 & local_bb4_reduction_5_i337);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_c1_ene1_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene1_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_c1_ene1_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene1_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene1_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene1_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_c1_ene1_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_c1_ene1_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_c1_ene1_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_c1_ene1_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_c1_ene1_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene1),
	.data_out(rnode_340to341_bb4_c1_ene1_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_c1_ene1_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_c1_ene1_0_reg_341_fifo.DATA_WIDTH = 32;
defparam rnode_340to341_bb4_c1_ene1_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_c1_ene1_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_c1_ene1_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene1_stall_in_1 = 1'b0;
assign rnode_340to341_bb4_c1_ene1_0_NO_SHIFT_REG = rnode_340to341_bb4_c1_ene1_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_c1_ene1_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_var__u30_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u30_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_var__u30_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u30_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u30_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_var__u30_1_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u30_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_var__u30_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u30_0_valid_out_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u30_0_stall_in_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u30_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_var__u30_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_var__u30_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_var__u30_0_stall_in_0_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_var__u30_0_valid_out_0_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_var__u30_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_var__u30),
	.data_out(rnode_340to341_bb4_var__u30_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_var__u30_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_var__u30_0_reg_341_fifo.DATA_WIDTH = 32;
defparam rnode_340to341_bb4_var__u30_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_var__u30_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_var__u30_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u30_stall_in_2 = 1'b0;
assign rnode_340to341_bb4_var__u30_0_stall_in_0_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_var__u30_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_var__u30_0_NO_SHIFT_REG = rnode_340to341_bb4_var__u30_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_var__u30_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_var__u30_1_NO_SHIFT_REG = rnode_340to341_bb4_var__u30_0_reg_341_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4__21_i507_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_1_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_valid_out_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_stall_in_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4__21_i507_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4__21_i507_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4__21_i507_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4__21_i507_0_stall_in_0_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4__21_i507_0_valid_out_0_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4__21_i507_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4__21_i507),
	.data_out(rnode_340to341_bb4__21_i507_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4__21_i507_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4__21_i507_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb4__21_i507_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4__21_i507_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4__21_i507_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i507_stall_in = 1'b0;
assign rnode_340to341_bb4__21_i507_0_stall_in_0_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4__21_i507_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4__21_i507_0_NO_SHIFT_REG = rnode_340to341_bb4__21_i507_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4__21_i507_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4__21_i507_1_NO_SHIFT_REG = rnode_340to341_bb4__21_i507_0_reg_341_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene5_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene5_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene5_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene5_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_c1_ene5_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_c1_ene5_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_c1_ene5_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_c1_ene5_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_c1_ene5_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_c1_ene5_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene5),
	.data_out(rnode_340to341_bb4_c1_ene5_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_c1_ene5_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_c1_ene5_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb4_c1_ene5_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_c1_ene5_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_c1_ene5_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene5_stall_in_1 = 1'b0;
assign rnode_340to341_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_340to341_bb4_c1_ene5_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_c1_ene5_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_xor_i496_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i496_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_xor_i496_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i496_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i496_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_xor_i496_1_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i496_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_xor_i496_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i496_0_valid_out_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i496_0_stall_in_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i496_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_xor_i496_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_xor_i496_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_xor_i496_0_stall_in_0_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_xor_i496_0_valid_out_0_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_xor_i496_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i496),
	.data_out(rnode_340to341_bb4_xor_i496_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_xor_i496_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_xor_i496_0_reg_341_fifo.DATA_WIDTH = 32;
defparam rnode_340to341_bb4_xor_i496_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_xor_i496_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_xor_i496_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i496_stall_in_2 = 1'b0;
assign rnode_340to341_bb4_xor_i496_0_stall_in_0_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_xor_i496_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_xor_i496_0_NO_SHIFT_REG = rnode_340to341_bb4_xor_i496_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_xor_i496_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_xor_i496_1_NO_SHIFT_REG = rnode_340to341_bb4_xor_i496_0_reg_341_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_348_349_0_inputs_ready;
 reg SFC_3_VALID_348_349_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_348_349_0_stall_in;
wire SFC_3_VALID_348_349_0_output_regs_ready;
 reg SFC_3_VALID_348_349_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_348_349_0_causedstall;

assign SFC_3_VALID_348_349_0_inputs_ready = 1'b1;
assign SFC_3_VALID_348_349_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_347_348_0_stall_in = 1'b0;
assign SFC_3_VALID_348_349_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_348_349_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_348_349_0_output_regs_ready)
		begin
			SFC_3_VALID_348_349_0_NO_SHIFT_REG <= SFC_3_VALID_347_348_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__24_i339_stall_local;
wire local_bb4__24_i339;

assign local_bb4__24_i339 = (local_bb4_cmp_i322 ? local_bb4_reduction_6_i338 : local_bb4_brmerge10_demorgan_i327);

// Register node:
//  * latency = 46
//  * capacity = 46
 logic rnode_341to387_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_341to387_bb4_c1_ene1_0_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene1_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to387_bb4_c1_ene1_0_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene1_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene1_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene1_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_341to387_bb4_c1_ene1_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to387_bb4_c1_ene1_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to387_bb4_c1_ene1_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_341to387_bb4_c1_ene1_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_341to387_bb4_c1_ene1_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_c1_ene1_0_NO_SHIFT_REG),
	.data_out(rnode_341to387_bb4_c1_ene1_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_341to387_bb4_c1_ene1_0_reg_387_fifo.DEPTH = 46;
defparam rnode_341to387_bb4_c1_ene1_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_341to387_bb4_c1_ene1_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to387_bb4_c1_ene1_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_341to387_bb4_c1_ene1_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to387_bb4_c1_ene1_0_NO_SHIFT_REG = rnode_341to387_bb4_c1_ene1_0_reg_387_NO_SHIFT_REG;
assign rnode_341to387_bb4_c1_ene1_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_341to387_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 46
//  * capacity = 46
 logic rnode_341to387_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene5_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene5_0_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene5_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene5_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_341to387_bb4_c1_ene5_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_341to387_bb4_c1_ene5_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to387_bb4_c1_ene5_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to387_bb4_c1_ene5_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_341to387_bb4_c1_ene5_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_341to387_bb4_c1_ene5_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_341to387_bb4_c1_ene5_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_341to387_bb4_c1_ene5_0_reg_387_fifo.DEPTH = 46;
defparam rnode_341to387_bb4_c1_ene5_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_341to387_bb4_c1_ene5_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to387_bb4_c1_ene5_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_341to387_bb4_c1_ene5_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to387_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_341to387_bb4_c1_ene5_0_reg_387_NO_SHIFT_REG;
assign rnode_341to387_bb4_c1_ene5_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_341to387_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__22_i508_stall_local;
wire [31:0] local_bb4__22_i508;

assign local_bb4__22_i508 = (rnode_340to341_bb4__21_i507_0_NO_SHIFT_REG ? rnode_340to341_bb4_var__u30_0_NO_SHIFT_REG : rnode_340to341_bb4_xor_i496_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i509_stall_local;
wire [31:0] local_bb4__23_i509;

assign local_bb4__23_i509 = (rnode_340to341_bb4__21_i507_1_NO_SHIFT_REG ? rnode_340to341_bb4_xor_i496_1_NO_SHIFT_REG : rnode_340to341_bb4_var__u30_1_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_3_VALID_349_350_0_inputs_ready;
 reg SFC_3_VALID_349_350_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_349_350_0_stall_in;
wire SFC_3_VALID_349_350_0_output_regs_ready;
 reg SFC_3_VALID_349_350_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_349_350_0_causedstall;

assign SFC_3_VALID_349_350_0_inputs_ready = 1'b1;
assign SFC_3_VALID_349_350_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_348_349_0_stall_in = 1'b0;
assign SFC_3_VALID_349_350_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_349_350_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_349_350_0_output_regs_ready)
		begin
			SFC_3_VALID_349_350_0_NO_SHIFT_REG <= SFC_3_VALID_348_349_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__25_i340_stall_local;
wire local_bb4__25_i340;

assign local_bb4__25_i340 = (local_bb4__24_i339 ? local_bb4_lnot14_i324 : local_bb4__mux_mux_mux_i334);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_c1_ene1_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene1_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_c1_ene1_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene1_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene1_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene1_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_c1_ene1_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_c1_ene1_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_c1_ene1_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_c1_ene1_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_c1_ene1_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_341to387_bb4_c1_ene1_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb4_c1_ene1_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_c1_ene1_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_c1_ene1_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb4_c1_ene1_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_c1_ene1_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_c1_ene1_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to387_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_c1_ene1_0_NO_SHIFT_REG = rnode_387to388_bb4_c1_ene1_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_c1_ene1_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_c1_ene5_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_1_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_c1_ene5_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_c1_ene5_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_c1_ene5_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_c1_ene5_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_c1_ene5_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_c1_ene5_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_341to387_bb4_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb4_c1_ene5_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_c1_ene5_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_c1_ene5_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb4_c1_ene5_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_c1_ene5_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_c1_ene5_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to387_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_c1_ene5_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_c1_ene5_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_387to388_bb4_c1_ene5_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_c1_ene5_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb4_c1_ene5_1_NO_SHIFT_REG = rnode_387to388_bb4_c1_ene5_0_reg_388_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i512_stall_local;
wire [31:0] local_bb4_shr18_i512;

assign local_bb4_shr18_i512 = (local_bb4__22_i508 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i510_stall_local;
wire [31:0] local_bb4_shr16_i510;

assign local_bb4_shr16_i510 = (local_bb4__23_i509 >> 32'h17);

// This section implements a registered operation.
// 
wire SFC_3_VALID_350_351_0_inputs_ready;
 reg SFC_3_VALID_350_351_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_350_351_0_stall_in;
wire SFC_3_VALID_350_351_0_output_regs_ready;
 reg SFC_3_VALID_350_351_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_350_351_0_causedstall;

assign SFC_3_VALID_350_351_0_inputs_ready = 1'b1;
assign SFC_3_VALID_350_351_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_349_350_0_stall_in = 1'b0;
assign SFC_3_VALID_350_351_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_350_351_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_350_351_0_output_regs_ready)
		begin
			SFC_3_VALID_350_351_0_NO_SHIFT_REG <= SFC_3_VALID_349_350_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__27_i342_stall_local;
wire local_bb4__27_i342;

assign local_bb4__27_i342 = (local_bb4__26_demorgan_i341 ? local_bb4__25_i340 : local_bb4__mux9_mux_i328);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u39_stall_local;
wire [31:0] local_bb4_var__u39;

assign local_bb4_var__u39 = rnode_387to388_bb4_c1_ene1_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_388to389_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_c1_ene5_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic rnode_388to389_bb4_c1_ene5_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_c1_ene5_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_c1_ene5_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_c1_ene5_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_c1_ene5_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_c1_ene5_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_c1_ene5_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_c1_ene5_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_c1_ene5_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(rnode_387to388_bb4_c1_ene5_1_NO_SHIFT_REG),
	.data_out(rnode_388to389_bb4_c1_ene5_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_c1_ene5_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_c1_ene5_0_reg_389_fifo.DATA_WIDTH = 1;
defparam rnode_388to389_bb4_c1_ene5_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_c1_ene5_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_c1_ene5_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_387to388_bb4_c1_ene5_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_388to389_bb4_c1_ene5_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_c1_ene5_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i513_stall_local;
wire [31:0] local_bb4_and19_i513;

assign local_bb4_and19_i513 = ((local_bb4_shr18_i512 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i538_stall_local;
wire [31:0] local_bb4_sub_i538;

assign local_bb4_sub_i538 = ((local_bb4_shr16_i510 & 32'h1FF) - (local_bb4_shr18_i512 & 32'h1FF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_351_352_0_inputs_ready;
 reg SFC_3_VALID_351_352_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_351_352_0_stall_in;
wire SFC_3_VALID_351_352_0_output_regs_ready;
 reg SFC_3_VALID_351_352_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_351_352_0_causedstall;

assign SFC_3_VALID_351_352_0_inputs_ready = 1'b1;
assign SFC_3_VALID_351_352_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_350_351_0_stall_in = 1'b0;
assign SFC_3_VALID_351_352_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_351_352_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_351_352_0_output_regs_ready)
		begin
			SFC_3_VALID_351_352_0_NO_SHIFT_REG <= SFC_3_VALID_350_351_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_xor_i316_valid_out;
wire local_bb4_xor_i316_stall_in;
wire local_bb4_add_i357_valid_out;
wire local_bb4_add_i357_stall_in;
wire local_bb4_conv_i_i348_valid_out;
wire local_bb4_conv_i_i348_stall_in;
wire local_bb4_conv1_i_i349_valid_out;
wire local_bb4_conv1_i_i349_stall_in;
wire local_bb4_reduction_0_i375_valid_out;
wire local_bb4_reduction_0_i375_stall_in;
wire local_bb4_var__u37_valid_out;
wire local_bb4_var__u37_stall_in;
wire local_bb4__29_i345_valid_out;
wire local_bb4__29_i345_stall_in;
wire local_bb4__29_i345_inputs_ready;
wire local_bb4__29_i345_stall_local;
wire local_bb4__29_i345;

assign local_bb4__29_i345_inputs_ready = (local_bb4_c1_enter_c1_eni8_valid_out_1_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni8_valid_out_2_NO_SHIFT_REG);
assign local_bb4__29_i345 = (local_bb4__28_i344 | local_bb4__27_i342);
assign local_bb4_xor_i316_valid_out = 1'b1;
assign local_bb4_add_i357_valid_out = 1'b1;
assign local_bb4_conv_i_i348_valid_out = 1'b1;
assign local_bb4_conv1_i_i349_valid_out = 1'b1;
assign local_bb4_reduction_0_i375_valid_out = 1'b1;
assign local_bb4_var__u37_valid_out = 1'b1;
assign local_bb4__29_i345_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni8_stall_in_1 = 1'b0;
assign local_bb4_c1_enter_c1_eni8_stall_in_2 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i_stall_local;
wire [31:0] local_bb4_shr2_i;

assign local_bb4_shr2_i = (local_bb4_var__u39 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and6_i_stall_local;
wire [31:0] local_bb4_and6_i;

assign local_bb4_and6_i = (local_bb4_var__u39 & 32'h7FFFFF);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_389to392_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to392_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_389to392_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_389to392_bb4_c1_ene5_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to392_bb4_c1_ene5_0_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb4_c1_ene5_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb4_c1_ene5_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb4_c1_ene5_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_389to392_bb4_c1_ene5_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to392_bb4_c1_ene5_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to392_bb4_c1_ene5_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_389to392_bb4_c1_ene5_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_389to392_bb4_c1_ene5_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_388to389_bb4_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_389to392_bb4_c1_ene5_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_389to392_bb4_c1_ene5_0_reg_392_fifo.DEPTH = 3;
defparam rnode_389to392_bb4_c1_ene5_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_389to392_bb4_c1_ene5_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to392_bb4_c1_ene5_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_389to392_bb4_c1_ene5_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_389to392_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_389to392_bb4_c1_ene5_0_reg_392_NO_SHIFT_REG;
assign rnode_389to392_bb4_c1_ene5_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_389to392_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i517_stall_local;
wire local_bb4_lnot23_i517;

assign local_bb4_lnot23_i517 = ((local_bb4_and19_i513 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i519_stall_local;
wire local_bb4_cmp27_i519;

assign local_bb4_cmp27_i519 = ((local_bb4_and19_i513 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and69_i_stall_local;
wire [31:0] local_bb4_and69_i;

assign local_bb4_and69_i = (local_bb4_sub_i538 & 32'hFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_352_353_0_inputs_ready;
 reg SFC_3_VALID_352_353_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_352_353_0_stall_in;
wire SFC_3_VALID_352_353_0_output_regs_ready;
 reg SFC_3_VALID_352_353_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_352_353_0_causedstall;

assign SFC_3_VALID_352_353_0_inputs_ready = 1'b1;
assign SFC_3_VALID_352_353_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_351_352_0_stall_in = 1'b0;
assign SFC_3_VALID_352_353_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_352_353_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_352_353_0_output_regs_ready)
		begin
			SFC_3_VALID_352_353_0_NO_SHIFT_REG <= SFC_3_VALID_351_352_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_xor_i316_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i316_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_xor_i316_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i316_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_xor_i316_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i316_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i316_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_xor_i316_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_xor_i316_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_xor_i316_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_xor_i316_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_xor_i316_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_xor_i316_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i316),
	.data_out(rnode_340to341_bb4_xor_i316_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_xor_i316_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_xor_i316_0_reg_341_fifo.DATA_WIDTH = 32;
defparam rnode_340to341_bb4_xor_i316_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_xor_i316_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_xor_i316_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i316_stall_in = 1'b0;
assign rnode_340to341_bb4_xor_i316_0_NO_SHIFT_REG = rnode_340to341_bb4_xor_i316_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_xor_i316_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_xor_i316_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_add_i357_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_add_i357_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_add_i357_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_add_i357_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_340to341_bb4_add_i357_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_add_i357_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_add_i357_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_add_i357_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_add_i357_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_add_i357_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_add_i357_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_add_i357_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_add_i357_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in((local_bb4_add_i357 & 32'h1FF)),
	.data_out(rnode_340to341_bb4_add_i357_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_add_i357_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_add_i357_0_reg_341_fifo.DATA_WIDTH = 32;
defparam rnode_340to341_bb4_add_i357_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_add_i357_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_add_i357_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add_i357_stall_in = 1'b0;
assign rnode_340to341_bb4_add_i357_0_NO_SHIFT_REG = rnode_340to341_bb4_add_i357_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_add_i357_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_add_i357_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_mul_i_i350_inputs_ready;
 reg local_bb4_mul_i_i350_valid_out_0_NO_SHIFT_REG;
wire local_bb4_mul_i_i350_stall_in_0;
 reg local_bb4_mul_i_i350_valid_out_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i350_stall_in_1;
wire local_bb4_mul_i_i350_output_regs_ready;
wire [63:0] local_bb4_mul_i_i350;
 reg local_bb4_mul_i_i350_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul_i_i350_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i350_causedstall;

acl_int_mult int_module_local_bb4_mul_i_i350 (
	.clock(clock),
	.dataa(((local_bb4_conv1_i_i349 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb4_conv_i_i348 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb4_mul_i_i350_output_regs_ready),
	.result(local_bb4_mul_i_i350)
);

defparam int_module_local_bb4_mul_i_i350.INPUT1_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i350.INPUT2_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i350.OUTPUT_WIDTH = 64;
defparam int_module_local_bb4_mul_i_i350.LATENCY = 3;
defparam int_module_local_bb4_mul_i_i350.SIGNED = 0;

assign local_bb4_mul_i_i350_inputs_ready = 1'b1;
assign local_bb4_mul_i_i350_output_regs_ready = 1'b1;
assign local_bb4_conv1_i_i349_stall_in = 1'b0;
assign local_bb4_conv_i_i348_stall_in = 1'b0;
assign local_bb4_mul_i_i350_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i350_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i350_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i350_output_regs_ready)
		begin
			local_bb4_mul_i_i350_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i350_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul_i_i350_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i350_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i350_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i350_output_regs_ready)
		begin
			local_bb4_mul_i_i350_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i350_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul_i_i350_stall_in_0))
			begin
				local_bb4_mul_i_i350_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_mul_i_i350_stall_in_1))
			begin
				local_bb4_mul_i_i350_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_reduction_0_i375_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_reduction_0_i375_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb4_reduction_0_i375_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_reduction_0_i375_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb4_reduction_0_i375_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_reduction_0_i375_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_reduction_0_i375_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_reduction_0_i375_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_reduction_0_i375_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_reduction_0_i375_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_reduction_0_i375_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_reduction_0_i375_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_reduction_0_i375_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_0_i375),
	.data_out(rnode_340to341_bb4_reduction_0_i375_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_reduction_0_i375_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_reduction_0_i375_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb4_reduction_0_i375_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_reduction_0_i375_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_reduction_0_i375_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_0_i375_stall_in = 1'b0;
assign rnode_340to341_bb4_reduction_0_i375_0_NO_SHIFT_REG = rnode_340to341_bb4_reduction_0_i375_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_reduction_0_i375_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_reduction_0_i375_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4_var__u37_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u37_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u37_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u37_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u37_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u37_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u37_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4_var__u37_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4_var__u37_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4_var__u37_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4_var__u37_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4_var__u37_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4_var__u37_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4_var__u37),
	.data_out(rnode_340to341_bb4_var__u37_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4_var__u37_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4_var__u37_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb4_var__u37_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4_var__u37_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4_var__u37_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u37_stall_in = 1'b0;
assign rnode_340to341_bb4_var__u37_0_NO_SHIFT_REG = rnode_340to341_bb4_var__u37_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4_var__u37_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_var__u37_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_340to341_bb4__29_i345_0_valid_out_NO_SHIFT_REG;
 logic rnode_340to341_bb4__29_i345_0_stall_in_NO_SHIFT_REG;
 logic rnode_340to341_bb4__29_i345_0_NO_SHIFT_REG;
 logic rnode_340to341_bb4__29_i345_0_reg_341_inputs_ready_NO_SHIFT_REG;
 logic rnode_340to341_bb4__29_i345_0_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4__29_i345_0_valid_out_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4__29_i345_0_stall_in_reg_341_NO_SHIFT_REG;
 logic rnode_340to341_bb4__29_i345_0_stall_out_reg_341_NO_SHIFT_REG;

acl_data_fifo rnode_340to341_bb4__29_i345_0_reg_341_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_340to341_bb4__29_i345_0_reg_341_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_340to341_bb4__29_i345_0_stall_in_reg_341_NO_SHIFT_REG),
	.valid_out(rnode_340to341_bb4__29_i345_0_valid_out_reg_341_NO_SHIFT_REG),
	.stall_out(rnode_340to341_bb4__29_i345_0_stall_out_reg_341_NO_SHIFT_REG),
	.data_in(local_bb4__29_i345),
	.data_out(rnode_340to341_bb4__29_i345_0_reg_341_NO_SHIFT_REG)
);

defparam rnode_340to341_bb4__29_i345_0_reg_341_fifo.DEPTH = 1;
defparam rnode_340to341_bb4__29_i345_0_reg_341_fifo.DATA_WIDTH = 1;
defparam rnode_340to341_bb4__29_i345_0_reg_341_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_340to341_bb4__29_i345_0_reg_341_fifo.IMPL = "shift_reg";

assign rnode_340to341_bb4__29_i345_0_reg_341_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__29_i345_stall_in = 1'b0;
assign rnode_340to341_bb4__29_i345_0_NO_SHIFT_REG = rnode_340to341_bb4__29_i345_0_reg_341_NO_SHIFT_REG;
assign rnode_340to341_bb4__29_i345_0_stall_in_reg_341_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4__29_i345_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or47_i_stall_local;
wire [31:0] local_bb4_or47_i;

assign local_bb4_or47_i = ((local_bb4_and6_i & 32'h7FFFFF) | 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene5_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene5_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene5_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene5_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_c1_ene5_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_c1_ene5_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_c1_ene5_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_c1_ene5_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_c1_ene5_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_c1_ene5_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_389to392_bb4_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb4_c1_ene5_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_c1_ene5_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_c1_ene5_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4_c1_ene5_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_c1_ene5_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_c1_ene5_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to392_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_392to393_bb4_c1_ene5_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_c1_ene5_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp70_i_stall_local;
wire local_bb4_cmp70_i;

assign local_bb4_cmp70_i = ((local_bb4_and69_i & 32'hFF) > 32'h1F);

// This section implements a registered operation.
// 
wire SFC_3_VALID_353_354_0_inputs_ready;
 reg SFC_3_VALID_353_354_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_353_354_0_stall_in;
wire SFC_3_VALID_353_354_0_output_regs_ready;
 reg SFC_3_VALID_353_354_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_353_354_0_causedstall;

assign SFC_3_VALID_353_354_0_inputs_ready = 1'b1;
assign SFC_3_VALID_353_354_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_352_353_0_stall_in = 1'b0;
assign SFC_3_VALID_353_354_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_353_354_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_353_354_0_output_regs_ready)
		begin
			SFC_3_VALID_353_354_0_NO_SHIFT_REG <= SFC_3_VALID_352_353_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_341to344_bb4_xor_i316_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to344_bb4_xor_i316_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_341to344_bb4_xor_i316_0_NO_SHIFT_REG;
 logic rnode_341to344_bb4_xor_i316_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to344_bb4_xor_i316_0_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4_xor_i316_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4_xor_i316_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4_xor_i316_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_341to344_bb4_xor_i316_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to344_bb4_xor_i316_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to344_bb4_xor_i316_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_341to344_bb4_xor_i316_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_341to344_bb4_xor_i316_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_xor_i316_0_NO_SHIFT_REG),
	.data_out(rnode_341to344_bb4_xor_i316_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_341to344_bb4_xor_i316_0_reg_344_fifo.DEPTH = 3;
defparam rnode_341to344_bb4_xor_i316_0_reg_344_fifo.DATA_WIDTH = 32;
defparam rnode_341to344_bb4_xor_i316_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to344_bb4_xor_i316_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_341to344_bb4_xor_i316_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_xor_i316_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb4_xor_i316_0_NO_SHIFT_REG = rnode_341to344_bb4_xor_i316_0_reg_344_NO_SHIFT_REG;
assign rnode_341to344_bb4_xor_i316_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb4_xor_i316_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_341to342_bb4_add_i357_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to342_bb4_add_i357_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_add_i357_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4_add_i357_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_add_i357_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_add_i357_0_valid_out_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_add_i357_0_stall_in_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_add_i357_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_341to342_bb4_add_i357_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to342_bb4_add_i357_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to342_bb4_add_i357_0_stall_in_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_341to342_bb4_add_i357_0_valid_out_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_341to342_bb4_add_i357_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in((rnode_340to341_bb4_add_i357_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_341to342_bb4_add_i357_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_341to342_bb4_add_i357_0_reg_342_fifo.DEPTH = 1;
defparam rnode_341to342_bb4_add_i357_0_reg_342_fifo.DATA_WIDTH = 32;
defparam rnode_341to342_bb4_add_i357_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to342_bb4_add_i357_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_341to342_bb4_add_i357_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_add_i357_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_add_i357_0_NO_SHIFT_REG = rnode_341to342_bb4_add_i357_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4_add_i357_0_stall_in_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_add_i357_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_conv3_i_i351_stall_local;
wire [31:0] local_bb4_conv3_i_i351;
wire [63:0] local_bb4_conv3_i_i351$ps;

assign local_bb4_conv3_i_i351$ps = (local_bb4_mul_i_i350 & 64'hFFFFFFFFFFFF);
assign local_bb4_conv3_i_i351 = local_bb4_conv3_i_i351$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u40_stall_local;
wire [63:0] local_bb4_var__u40;

assign local_bb4_var__u40 = ((local_bb4_mul_i_i350 & 64'hFFFFFFFFFFFF) >> 64'h18);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_341to344_bb4_reduction_0_i375_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to344_bb4_reduction_0_i375_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to344_bb4_reduction_0_i375_0_NO_SHIFT_REG;
 logic rnode_341to344_bb4_reduction_0_i375_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to344_bb4_reduction_0_i375_0_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4_reduction_0_i375_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4_reduction_0_i375_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4_reduction_0_i375_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_341to344_bb4_reduction_0_i375_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to344_bb4_reduction_0_i375_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to344_bb4_reduction_0_i375_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_341to344_bb4_reduction_0_i375_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_341to344_bb4_reduction_0_i375_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_reduction_0_i375_0_NO_SHIFT_REG),
	.data_out(rnode_341to344_bb4_reduction_0_i375_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_341to344_bb4_reduction_0_i375_0_reg_344_fifo.DEPTH = 3;
defparam rnode_341to344_bb4_reduction_0_i375_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_341to344_bb4_reduction_0_i375_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to344_bb4_reduction_0_i375_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_341to344_bb4_reduction_0_i375_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_reduction_0_i375_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb4_reduction_0_i375_0_NO_SHIFT_REG = rnode_341to344_bb4_reduction_0_i375_0_reg_344_NO_SHIFT_REG;
assign rnode_341to344_bb4_reduction_0_i375_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb4_reduction_0_i375_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_341to342_bb4_var__u37_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to342_bb4_var__u37_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to342_bb4_var__u37_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4_var__u37_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to342_bb4_var__u37_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_var__u37_0_valid_out_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_var__u37_0_stall_in_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_var__u37_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_341to342_bb4_var__u37_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to342_bb4_var__u37_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to342_bb4_var__u37_0_stall_in_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_341to342_bb4_var__u37_0_valid_out_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_341to342_bb4_var__u37_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4_var__u37_0_NO_SHIFT_REG),
	.data_out(rnode_341to342_bb4_var__u37_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_341to342_bb4_var__u37_0_reg_342_fifo.DEPTH = 1;
defparam rnode_341to342_bb4_var__u37_0_reg_342_fifo.DATA_WIDTH = 1;
defparam rnode_341to342_bb4_var__u37_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to342_bb4_var__u37_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_341to342_bb4_var__u37_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4_var__u37_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_var__u37_0_NO_SHIFT_REG = rnode_341to342_bb4_var__u37_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4_var__u37_0_stall_in_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_var__u37_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_341to344_bb4__29_i345_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to344_bb4__29_i345_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to344_bb4__29_i345_0_NO_SHIFT_REG;
 logic rnode_341to344_bb4__29_i345_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to344_bb4__29_i345_0_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4__29_i345_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4__29_i345_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_341to344_bb4__29_i345_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_341to344_bb4__29_i345_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to344_bb4__29_i345_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to344_bb4__29_i345_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_341to344_bb4__29_i345_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_341to344_bb4__29_i345_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(rnode_340to341_bb4__29_i345_0_NO_SHIFT_REG),
	.data_out(rnode_341to344_bb4__29_i345_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_341to344_bb4__29_i345_0_reg_344_fifo.DEPTH = 3;
defparam rnode_341to344_bb4__29_i345_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_341to344_bb4__29_i345_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to344_bb4__29_i345_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_341to344_bb4__29_i345_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_340to341_bb4__29_i345_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb4__29_i345_0_NO_SHIFT_REG = rnode_341to344_bb4__29_i345_0_reg_344_NO_SHIFT_REG;
assign rnode_341to344_bb4__29_i345_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_341to344_bb4__29_i345_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_conv1_i_i_stall_local;
wire [63:0] local_bb4_conv1_i_i;

assign local_bb4_conv1_i_i[63:32] = 32'h0;
assign local_bb4_conv1_i_i[31:0] = ((local_bb4_or47_i & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i508_valid_out_1;
wire local_bb4__22_i508_stall_in_1;
wire local_bb4__23_i509_valid_out_1;
wire local_bb4__23_i509_stall_in_1;
wire local_bb4_shr16_i510_valid_out_1;
wire local_bb4_shr16_i510_stall_in_1;
wire local_bb4_lnot23_i517_valid_out;
wire local_bb4_lnot23_i517_stall_in;
wire local_bb4_cmp27_i519_valid_out;
wire local_bb4_cmp27_i519_stall_in;
wire local_bb4_align_0_i539_valid_out;
wire local_bb4_align_0_i539_stall_in;
wire local_bb4_align_0_i539_inputs_ready;
wire local_bb4_align_0_i539_stall_local;
wire [31:0] local_bb4_align_0_i539;

assign local_bb4_align_0_i539_inputs_ready = (rnode_340to341_bb4__21_i507_0_valid_out_0_NO_SHIFT_REG & rnode_340to341_bb4_var__u30_0_valid_out_0_NO_SHIFT_REG & rnode_340to341_bb4_xor_i496_0_valid_out_0_NO_SHIFT_REG & rnode_340to341_bb4__21_i507_0_valid_out_1_NO_SHIFT_REG & rnode_340to341_bb4_xor_i496_0_valid_out_1_NO_SHIFT_REG & rnode_340to341_bb4_var__u30_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_align_0_i539 = (local_bb4_cmp70_i ? 32'h1F : (local_bb4_and69_i & 32'hFF));
assign local_bb4__22_i508_valid_out_1 = 1'b1;
assign local_bb4__23_i509_valid_out_1 = 1'b1;
assign local_bb4_shr16_i510_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i517_valid_out = 1'b1;
assign local_bb4_cmp27_i519_valid_out = 1'b1;
assign local_bb4_align_0_i539_valid_out = 1'b1;
assign rnode_340to341_bb4__21_i507_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_var__u30_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_xor_i496_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4__21_i507_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_xor_i496_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_340to341_bb4_var__u30_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_354_355_0_inputs_ready;
 reg SFC_3_VALID_354_355_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_354_355_0_stall_in;
wire SFC_3_VALID_354_355_0_output_regs_ready;
 reg SFC_3_VALID_354_355_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_354_355_0_causedstall;

assign SFC_3_VALID_354_355_0_inputs_ready = 1'b1;
assign SFC_3_VALID_354_355_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_353_354_0_stall_in = 1'b0;
assign SFC_3_VALID_354_355_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_354_355_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_354_355_0_output_regs_ready)
		begin
			SFC_3_VALID_354_355_0_NO_SHIFT_REG <= SFC_3_VALID_353_354_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4_xor_i316_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb4_xor_i316_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_xor_i316_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4_xor_i316_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_xor_i316_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_xor_i316_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_xor_i316_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_xor_i316_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4_xor_i316_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4_xor_i316_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4_xor_i316_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4_xor_i316_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4_xor_i316_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(rnode_341to344_bb4_xor_i316_0_NO_SHIFT_REG),
	.data_out(rnode_344to345_bb4_xor_i316_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4_xor_i316_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4_xor_i316_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_344to345_bb4_xor_i316_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4_xor_i316_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4_xor_i316_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to344_bb4_xor_i316_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_xor_i316_0_NO_SHIFT_REG = rnode_344to345_bb4_xor_i316_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4_xor_i316_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_xor_i316_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_add_i357_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_add_i357_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_add_i357_1_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_add_i357_2_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_add_i357_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_valid_out_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_stall_in_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_add_i357_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_add_i357_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_add_i357_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_add_i357_0_stall_in_0_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_add_i357_0_valid_out_0_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_add_i357_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((rnode_341to342_bb4_add_i357_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_342to343_bb4_add_i357_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_add_i357_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_add_i357_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb4_add_i357_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_add_i357_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_add_i357_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4_add_i357_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_add_i357_0_stall_in_0_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_add_i357_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_add_i357_0_NO_SHIFT_REG = rnode_342to343_bb4_add_i357_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_add_i357_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_add_i357_1_NO_SHIFT_REG = rnode_342to343_bb4_add_i357_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_add_i357_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_add_i357_2_NO_SHIFT_REG = rnode_342to343_bb4_add_i357_0_reg_343_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i16_i354_stall_local;
wire [31:0] local_bb4_shr_i16_i354;

assign local_bb4_shr_i16_i354 = (local_bb4_conv3_i_i351 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i18_i356_stall_local;
wire [31:0] local_bb4_shl1_i18_i356;

assign local_bb4_shl1_i18_i356 = (local_bb4_conv3_i_i351 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u41_stall_local;
wire [31:0] local_bb4_var__u41;

assign local_bb4_var__u41 = (local_bb4_conv3_i_i351 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i_i364_stall_local;
wire [31:0] local_bb4_shl1_i_i364;

assign local_bb4_shl1_i_i364 = (local_bb4_conv3_i_i351 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb4__tr_i352_stall_local;
wire [31:0] local_bb4__tr_i352;
wire [63:0] local_bb4__tr_i352$ps;

assign local_bb4__tr_i352$ps = (local_bb4_var__u40 & 64'hFFFFFF);
assign local_bb4__tr_i352 = local_bb4__tr_i352$ps[31:0];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4_reduction_0_i375_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb4_reduction_0_i375_0_stall_in_NO_SHIFT_REG;
 logic rnode_344to345_bb4_reduction_0_i375_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4_reduction_0_i375_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_344to345_bb4_reduction_0_i375_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_reduction_0_i375_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_reduction_0_i375_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_reduction_0_i375_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4_reduction_0_i375_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4_reduction_0_i375_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4_reduction_0_i375_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4_reduction_0_i375_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4_reduction_0_i375_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(rnode_341to344_bb4_reduction_0_i375_0_NO_SHIFT_REG),
	.data_out(rnode_344to345_bb4_reduction_0_i375_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4_reduction_0_i375_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4_reduction_0_i375_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_344to345_bb4_reduction_0_i375_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4_reduction_0_i375_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4_reduction_0_i375_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to344_bb4_reduction_0_i375_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_reduction_0_i375_0_NO_SHIFT_REG = rnode_344to345_bb4_reduction_0_i375_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4_reduction_0_i375_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_reduction_0_i375_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_var__u37_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb4_var__u37_0_stall_in_NO_SHIFT_REG;
 logic rnode_342to343_bb4_var__u37_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_var__u37_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic rnode_342to343_bb4_var__u37_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_var__u37_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_var__u37_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_var__u37_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_var__u37_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_var__u37_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_var__u37_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_var__u37_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_var__u37_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in(rnode_341to342_bb4_var__u37_0_NO_SHIFT_REG),
	.data_out(rnode_342to343_bb4_var__u37_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_var__u37_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_var__u37_0_reg_343_fifo.DATA_WIDTH = 1;
defparam rnode_342to343_bb4_var__u37_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_var__u37_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_var__u37_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4_var__u37_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_var__u37_0_NO_SHIFT_REG = rnode_342to343_bb4_var__u37_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_var__u37_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_var__u37_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4__29_i345_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb4__29_i345_0_stall_in_NO_SHIFT_REG;
 logic rnode_344to345_bb4__29_i345_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4__29_i345_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_344to345_bb4__29_i345_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__29_i345_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__29_i345_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__29_i345_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4__29_i345_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4__29_i345_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4__29_i345_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4__29_i345_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4__29_i345_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(rnode_341to344_bb4__29_i345_0_NO_SHIFT_REG),
	.data_out(rnode_344to345_bb4__29_i345_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4__29_i345_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4__29_i345_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_344to345_bb4__29_i345_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4__29_i345_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4__29_i345_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to344_bb4__29_i345_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__29_i345_0_NO_SHIFT_REG = rnode_344to345_bb4__29_i345_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4__29_i345_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__29_i345_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_341to342_bb4__22_i508_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4__22_i508_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4__22_i508_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4__22_i508_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_341to342_bb4__22_i508_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4__22_i508_1_NO_SHIFT_REG;
 logic rnode_341to342_bb4__22_i508_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4__22_i508_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4__22_i508_0_valid_out_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4__22_i508_0_stall_in_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4__22_i508_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_341to342_bb4__22_i508_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to342_bb4__22_i508_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to342_bb4__22_i508_0_stall_in_0_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_341to342_bb4__22_i508_0_valid_out_0_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_341to342_bb4__22_i508_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in(local_bb4__22_i508),
	.data_out(rnode_341to342_bb4__22_i508_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_341to342_bb4__22_i508_0_reg_342_fifo.DEPTH = 1;
defparam rnode_341to342_bb4__22_i508_0_reg_342_fifo.DATA_WIDTH = 32;
defparam rnode_341to342_bb4__22_i508_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to342_bb4__22_i508_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_341to342_bb4__22_i508_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i508_stall_in_1 = 1'b0;
assign rnode_341to342_bb4__22_i508_0_stall_in_0_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4__22_i508_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4__22_i508_0_NO_SHIFT_REG = rnode_341to342_bb4__22_i508_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4__22_i508_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4__22_i508_1_NO_SHIFT_REG = rnode_341to342_bb4__22_i508_0_reg_342_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_341to342_bb4__23_i509_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4__23_i509_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4__23_i509_1_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4__23_i509_2_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4__23_i509_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_valid_out_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_stall_in_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4__23_i509_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_341to342_bb4__23_i509_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to342_bb4__23_i509_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to342_bb4__23_i509_0_stall_in_0_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_341to342_bb4__23_i509_0_valid_out_0_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_341to342_bb4__23_i509_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in(local_bb4__23_i509),
	.data_out(rnode_341to342_bb4__23_i509_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_341to342_bb4__23_i509_0_reg_342_fifo.DEPTH = 1;
defparam rnode_341to342_bb4__23_i509_0_reg_342_fifo.DATA_WIDTH = 32;
defparam rnode_341to342_bb4__23_i509_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to342_bb4__23_i509_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_341to342_bb4__23_i509_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i509_stall_in_1 = 1'b0;
assign rnode_341to342_bb4__23_i509_0_stall_in_0_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4__23_i509_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4__23_i509_0_NO_SHIFT_REG = rnode_341to342_bb4__23_i509_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4__23_i509_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4__23_i509_1_NO_SHIFT_REG = rnode_341to342_bb4__23_i509_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4__23_i509_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4__23_i509_2_NO_SHIFT_REG = rnode_341to342_bb4__23_i509_0_reg_342_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_341to343_bb4_shr16_i510_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_341to343_bb4_shr16_i510_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_341to343_bb4_shr16_i510_0_NO_SHIFT_REG;
 logic rnode_341to343_bb4_shr16_i510_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_341to343_bb4_shr16_i510_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_341to343_bb4_shr16_i510_1_NO_SHIFT_REG;
 logic rnode_341to343_bb4_shr16_i510_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to343_bb4_shr16_i510_0_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb4_shr16_i510_0_valid_out_0_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb4_shr16_i510_0_stall_in_0_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb4_shr16_i510_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_341to343_bb4_shr16_i510_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to343_bb4_shr16_i510_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to343_bb4_shr16_i510_0_stall_in_0_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_341to343_bb4_shr16_i510_0_valid_out_0_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_341to343_bb4_shr16_i510_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i510 & 32'h1FF)),
	.data_out(rnode_341to343_bb4_shr16_i510_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_341to343_bb4_shr16_i510_0_reg_343_fifo.DEPTH = 2;
defparam rnode_341to343_bb4_shr16_i510_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_341to343_bb4_shr16_i510_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to343_bb4_shr16_i510_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_341to343_bb4_shr16_i510_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i510_stall_in_1 = 1'b0;
assign rnode_341to343_bb4_shr16_i510_0_stall_in_0_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_341to343_bb4_shr16_i510_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_341to343_bb4_shr16_i510_0_NO_SHIFT_REG = rnode_341to343_bb4_shr16_i510_0_reg_343_NO_SHIFT_REG;
assign rnode_341to343_bb4_shr16_i510_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_341to343_bb4_shr16_i510_1_NO_SHIFT_REG = rnode_341to343_bb4_shr16_i510_0_reg_343_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_341to342_bb4_lnot23_i517_0_valid_out_NO_SHIFT_REG;
 logic rnode_341to342_bb4_lnot23_i517_0_stall_in_NO_SHIFT_REG;
 logic rnode_341to342_bb4_lnot23_i517_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4_lnot23_i517_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to342_bb4_lnot23_i517_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_lnot23_i517_0_valid_out_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_lnot23_i517_0_stall_in_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_lnot23_i517_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_341to342_bb4_lnot23_i517_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to342_bb4_lnot23_i517_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to342_bb4_lnot23_i517_0_stall_in_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_341to342_bb4_lnot23_i517_0_valid_out_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_341to342_bb4_lnot23_i517_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i517),
	.data_out(rnode_341to342_bb4_lnot23_i517_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_341to342_bb4_lnot23_i517_0_reg_342_fifo.DEPTH = 1;
defparam rnode_341to342_bb4_lnot23_i517_0_reg_342_fifo.DATA_WIDTH = 1;
defparam rnode_341to342_bb4_lnot23_i517_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to342_bb4_lnot23_i517_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_341to342_bb4_lnot23_i517_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i517_stall_in = 1'b0;
assign rnode_341to342_bb4_lnot23_i517_0_NO_SHIFT_REG = rnode_341to342_bb4_lnot23_i517_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4_lnot23_i517_0_stall_in_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_lnot23_i517_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_341to343_bb4_cmp27_i519_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_1_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_2_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_valid_out_0_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_stall_in_0_reg_343_NO_SHIFT_REG;
 logic rnode_341to343_bb4_cmp27_i519_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_341to343_bb4_cmp27_i519_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to343_bb4_cmp27_i519_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to343_bb4_cmp27_i519_0_stall_in_0_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_341to343_bb4_cmp27_i519_0_valid_out_0_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_341to343_bb4_cmp27_i519_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i519),
	.data_out(rnode_341to343_bb4_cmp27_i519_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_341to343_bb4_cmp27_i519_0_reg_343_fifo.DEPTH = 2;
defparam rnode_341to343_bb4_cmp27_i519_0_reg_343_fifo.DATA_WIDTH = 1;
defparam rnode_341to343_bb4_cmp27_i519_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to343_bb4_cmp27_i519_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_341to343_bb4_cmp27_i519_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i519_stall_in = 1'b0;
assign rnode_341to343_bb4_cmp27_i519_0_stall_in_0_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_341to343_bb4_cmp27_i519_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_341to343_bb4_cmp27_i519_0_NO_SHIFT_REG = rnode_341to343_bb4_cmp27_i519_0_reg_343_NO_SHIFT_REG;
assign rnode_341to343_bb4_cmp27_i519_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_341to343_bb4_cmp27_i519_1_NO_SHIFT_REG = rnode_341to343_bb4_cmp27_i519_0_reg_343_NO_SHIFT_REG;
assign rnode_341to343_bb4_cmp27_i519_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_341to343_bb4_cmp27_i519_2_NO_SHIFT_REG = rnode_341to343_bb4_cmp27_i519_0_reg_343_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_341to342_bb4_align_0_i539_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_align_0_i539_0_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_align_0_i539_1_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_align_0_i539_2_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_align_0_i539_3_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_align_0_i539_4_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_reg_342_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_341to342_bb4_align_0_i539_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_valid_out_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_stall_in_0_reg_342_NO_SHIFT_REG;
 logic rnode_341to342_bb4_align_0_i539_0_stall_out_reg_342_NO_SHIFT_REG;

acl_data_fifo rnode_341to342_bb4_align_0_i539_0_reg_342_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_341to342_bb4_align_0_i539_0_reg_342_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_341to342_bb4_align_0_i539_0_stall_in_0_reg_342_NO_SHIFT_REG),
	.valid_out(rnode_341to342_bb4_align_0_i539_0_valid_out_0_reg_342_NO_SHIFT_REG),
	.stall_out(rnode_341to342_bb4_align_0_i539_0_stall_out_reg_342_NO_SHIFT_REG),
	.data_in((local_bb4_align_0_i539 & 32'hFF)),
	.data_out(rnode_341to342_bb4_align_0_i539_0_reg_342_NO_SHIFT_REG)
);

defparam rnode_341to342_bb4_align_0_i539_0_reg_342_fifo.DEPTH = 1;
defparam rnode_341to342_bb4_align_0_i539_0_reg_342_fifo.DATA_WIDTH = 32;
defparam rnode_341to342_bb4_align_0_i539_0_reg_342_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_341to342_bb4_align_0_i539_0_reg_342_fifo.IMPL = "shift_reg";

assign rnode_341to342_bb4_align_0_i539_0_reg_342_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_align_0_i539_stall_in = 1'b0;
assign rnode_341to342_bb4_align_0_i539_0_stall_in_0_reg_342_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_align_0_i539_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4_align_0_i539_0_NO_SHIFT_REG = rnode_341to342_bb4_align_0_i539_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4_align_0_i539_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4_align_0_i539_1_NO_SHIFT_REG = rnode_341to342_bb4_align_0_i539_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4_align_0_i539_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4_align_0_i539_2_NO_SHIFT_REG = rnode_341to342_bb4_align_0_i539_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4_align_0_i539_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4_align_0_i539_3_NO_SHIFT_REG = rnode_341to342_bb4_align_0_i539_0_reg_342_NO_SHIFT_REG;
assign rnode_341to342_bb4_align_0_i539_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_341to342_bb4_align_0_i539_4_NO_SHIFT_REG = rnode_341to342_bb4_align_0_i539_0_reg_342_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_355_356_0_inputs_ready;
 reg SFC_3_VALID_355_356_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_355_356_0_stall_in;
wire SFC_3_VALID_355_356_0_output_regs_ready;
 reg SFC_3_VALID_355_356_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_355_356_0_causedstall;

assign SFC_3_VALID_355_356_0_inputs_ready = 1'b1;
assign SFC_3_VALID_355_356_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_354_355_0_stall_in = 1'b0;
assign SFC_3_VALID_355_356_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_355_356_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_355_356_0_output_regs_ready)
		begin
			SFC_3_VALID_355_356_0_NO_SHIFT_REG <= SFC_3_VALID_354_355_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and4_i317_stall_local;
wire [31:0] local_bb4_and4_i317;

assign local_bb4_and4_i317 = (rnode_344to345_bb4_xor_i316_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_inc_i360_stall_local;
wire [31:0] local_bb4_inc_i360;

assign local_bb4_inc_i360 = ((rnode_342to343_bb4_add_i357_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp50_not_i365_stall_local;
wire local_bb4_cmp50_not_i365;

assign local_bb4_cmp50_not_i365 = ((rnode_342to343_bb4_add_i357_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i362_stall_local;
wire [31:0] local_bb4_shr_i_i362;

assign local_bb4_shr_i_i362 = ((local_bb4_var__u41 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i15_i353_stall_local;
wire [31:0] local_bb4_shl_i15_i353;

assign local_bb4_shl_i15_i353 = ((local_bb4__tr_i352 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb4_and48_i358_stall_local;
wire [31:0] local_bb4_and48_i358;

assign local_bb4_and48_i358 = ((local_bb4__tr_i352 & 32'hFFFFFF) & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i515_stall_local;
wire [31:0] local_bb4_and21_i515;

assign local_bb4_and21_i515 = (rnode_341to342_bb4__22_i508_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i514_valid_out;
wire local_bb4_and20_i514_stall_in;
wire local_bb4_and20_i514_inputs_ready;
wire local_bb4_and20_i514_stall_local;
wire [31:0] local_bb4_and20_i514;

assign local_bb4_and20_i514_inputs_ready = rnode_341to342_bb4__23_i509_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i514 = (rnode_341to342_bb4__23_i509_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i514_valid_out = 1'b1;
assign rnode_341to342_bb4__23_i509_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i520_valid_out;
wire local_bb4_and35_i520_stall_in;
wire local_bb4_and35_i520_inputs_ready;
wire local_bb4_and35_i520_stall_local;
wire [31:0] local_bb4_and35_i520;

assign local_bb4_and35_i520_inputs_ready = rnode_341to342_bb4__23_i509_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i520 = (rnode_341to342_bb4__23_i509_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i520_valid_out = 1'b1;
assign rnode_341to342_bb4__23_i509_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor36_i_stall_local;
wire [31:0] local_bb4_xor36_i;

assign local_bb4_xor36_i = (rnode_341to342_bb4__23_i509_2_NO_SHIFT_REG ^ rnode_341to342_bb4__22_i508_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i511_stall_local;
wire [31:0] local_bb4_and17_i511;

assign local_bb4_and17_i511 = ((rnode_341to343_bb4_shr16_i510_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_shr16_i510_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shr16_i510_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_shr16_i510_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shr16_i510_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_shr16_i510_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shr16_i510_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shr16_i510_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shr16_i510_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_shr16_i510_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_shr16_i510_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_shr16_i510_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_shr16_i510_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_shr16_i510_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((rnode_341to343_bb4_shr16_i510_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_343to345_bb4_shr16_i510_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_shr16_i510_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_shr16_i510_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_343to345_bb4_shr16_i510_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_shr16_i510_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_shr16_i510_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_341to343_bb4_shr16_i510_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_shr16_i510_0_NO_SHIFT_REG = rnode_343to345_bb4_shr16_i510_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_shr16_i510_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_shr16_i510_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and94_i_stall_local;
wire [31:0] local_bb4_and94_i;

assign local_bb4_and94_i = ((rnode_341to342_bb4_align_0_i539_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and96_i_stall_local;
wire [31:0] local_bb4_and96_i;

assign local_bb4_and96_i = ((rnode_341to342_bb4_align_0_i539_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and116_i_stall_local;
wire [31:0] local_bb4_and116_i;

assign local_bb4_and116_i = ((rnode_341to342_bb4_align_0_i539_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and131_i_stall_local;
wire [31:0] local_bb4_and131_i;

assign local_bb4_and131_i = ((rnode_341to342_bb4_align_0_i539_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and150_i_stall_local;
wire [31:0] local_bb4_and150_i;

assign local_bb4_and150_i = ((rnode_341to342_bb4_align_0_i539_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements a registered operation.
// 
wire SFC_3_VALID_356_357_0_inputs_ready;
 reg SFC_3_VALID_356_357_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_356_357_0_stall_in;
wire SFC_3_VALID_356_357_0_output_regs_ready;
 reg SFC_3_VALID_356_357_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_356_357_0_causedstall;

assign SFC_3_VALID_356_357_0_inputs_ready = 1'b1;
assign SFC_3_VALID_356_357_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_355_356_0_stall_in = 1'b0;
assign SFC_3_VALID_356_357_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_356_357_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_356_357_0_output_regs_ready)
		begin
			SFC_3_VALID_356_357_0_NO_SHIFT_REG <= SFC_3_VALID_355_356_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or_i17_i355_stall_local;
wire [31:0] local_bb4_or_i17_i355;

assign local_bb4_or_i17_i355 = ((local_bb4_shl_i15_i353 & 32'hFFFF00) | (local_bb4_shr_i16_i354 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool49_i359_stall_local;
wire local_bb4_tobool49_i359;

assign local_bb4_tobool49_i359 = ((local_bb4_and48_i358 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i524_stall_local;
wire local_bb4_lnot33_not_i524;

assign local_bb4_lnot33_not_i524 = ((local_bb4_and21_i515 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or65_i_stall_local;
wire [31:0] local_bb4_or65_i;

assign local_bb4_or65_i = ((local_bb4_and21_i515 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_and20_i514_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and20_i514_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_and20_i514_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and20_i514_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and20_i514_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_and20_i514_1_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and20_i514_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_and20_i514_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and20_i514_0_valid_out_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and20_i514_0_stall_in_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and20_i514_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_and20_i514_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_and20_i514_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_and20_i514_0_stall_in_0_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_and20_i514_0_valid_out_0_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_and20_i514_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i514 & 32'h7FFFFF)),
	.data_out(rnode_342to343_bb4_and20_i514_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_and20_i514_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_and20_i514_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb4_and20_i514_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_and20_i514_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_and20_i514_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i514_stall_in = 1'b0;
assign rnode_342to343_bb4_and20_i514_0_stall_in_0_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_and20_i514_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_and20_i514_0_NO_SHIFT_REG = rnode_342to343_bb4_and20_i514_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_and20_i514_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_and20_i514_1_NO_SHIFT_REG = rnode_342to343_bb4_and20_i514_0_reg_343_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_and35_i520_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and35_i520_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_and35_i520_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and35_i520_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_and35_i520_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and35_i520_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and35_i520_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and35_i520_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_and35_i520_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_and35_i520_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_and35_i520_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_and35_i520_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_and35_i520_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i520 & 32'h80000000)),
	.data_out(rnode_342to343_bb4_and35_i520_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_and35_i520_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_and35_i520_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb4_and35_i520_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_and35_i520_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_and35_i520_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i520_stall_in = 1'b0;
assign rnode_342to343_bb4_and35_i520_0_NO_SHIFT_REG = rnode_342to343_bb4_and35_i520_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_and35_i520_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_and35_i520_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp38_i_stall_local;
wire local_bb4_cmp38_i;

assign local_bb4_cmp38_i = ($signed(local_bb4_xor36_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor36_lobit_i_stall_local;
wire [31:0] local_bb4_xor36_lobit_i;

assign local_bb4_xor36_lobit_i = ($signed(local_bb4_xor36_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and37_lobit_i_stall_local;
wire [31:0] local_bb4_and37_lobit_i;

assign local_bb4_and37_lobit_i = (local_bb4_xor36_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i516_stall_local;
wire local_bb4_lnot_i516;

assign local_bb4_lnot_i516 = ((local_bb4_and17_i511 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i518_stall_local;
wire local_bb4_cmp25_i518;

assign local_bb4_cmp25_i518 = ((local_bb4_and17_i511 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp97_i_stall_local;
wire local_bb4_cmp97_i;

assign local_bb4_cmp97_i = ((local_bb4_and96_i & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp117_i_stall_local;
wire local_bb4_cmp117_i;

assign local_bb4_cmp117_i = ((local_bb4_and116_i & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp132_not_i_stall_local;
wire local_bb4_cmp132_not_i;

assign local_bb4_cmp132_not_i = ((local_bb4_and131_i & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i550_stall_local;
wire local_bb4_Pivot20_i550;

assign local_bb4_Pivot20_i550 = ((local_bb4_and150_i & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i551_stall_local;
wire local_bb4_SwitchLeaf_i551;

assign local_bb4_SwitchLeaf_i551 = ((local_bb4_and150_i & 32'h3) == 32'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_357_358_0_inputs_ready;
 reg SFC_3_VALID_357_358_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_357_358_0_stall_in;
wire SFC_3_VALID_357_358_0_output_regs_ready;
 reg SFC_3_VALID_357_358_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_357_358_0_causedstall;

assign SFC_3_VALID_357_358_0_inputs_ready = 1'b1;
assign SFC_3_VALID_357_358_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_356_357_0_stall_in = 1'b0;
assign SFC_3_VALID_357_358_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_357_358_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_357_358_0_output_regs_ready)
		begin
			SFC_3_VALID_357_358_0_NO_SHIFT_REG <= SFC_3_VALID_356_357_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_i361_stall_local;
wire [31:0] local_bb4_shl_i_i361;

assign local_bb4_shl_i_i361 = ((local_bb4_or_i17_i355 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__31_i366_stall_local;
wire local_bb4__31_i366;

assign local_bb4__31_i366 = (local_bb4_tobool49_i359 & local_bb4_cmp50_not_i365);

// This section implements an unregistered operation.
// 
wire local_bb4_shl66_i_stall_local;
wire [31:0] local_bb4_shl66_i;

assign local_bb4_shl66_i = ((local_bb4_or65_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i522_stall_local;
wire local_bb4_lnot30_i522;

assign local_bb4_lnot30_i522 = ((rnode_342to343_bb4_and20_i514_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i534_stall_local;
wire [31:0] local_bb4_or_i534;

assign local_bb4_or_i534 = ((rnode_342to343_bb4_and20_i514_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_and35_i520_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and35_i520_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_and35_i520_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and35_i520_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_and35_i520_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and35_i520_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and35_i520_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and35_i520_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_and35_i520_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_and35_i520_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_and35_i520_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_and35_i520_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_and35_i520_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((rnode_342to343_bb4_and35_i520_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_343to345_bb4_and35_i520_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_and35_i520_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_and35_i520_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_343to345_bb4_and35_i520_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_and35_i520_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_and35_i520_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_and35_i520_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_and35_i520_0_NO_SHIFT_REG = rnode_343to345_bb4_and35_i520_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_and35_i520_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_and35_i520_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i521_stall_local;
wire local_bb4_cmp25_not_i521;

assign local_bb4_cmp25_not_i521 = (local_bb4_cmp25_i518 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u42_stall_local;
wire local_bb4_var__u42;

assign local_bb4_var__u42 = (local_bb4_cmp25_i518 | rnode_341to343_bb4_cmp27_i519_2_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_3_VALID_358_359_0_inputs_ready;
 reg SFC_3_VALID_358_359_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_358_359_0_stall_in;
wire SFC_3_VALID_358_359_0_output_regs_ready;
 reg SFC_3_VALID_358_359_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_358_359_0_causedstall;

assign SFC_3_VALID_358_359_0_inputs_ready = 1'b1;
assign SFC_3_VALID_358_359_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_357_358_0_stall_in = 1'b0;
assign SFC_3_VALID_358_359_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_358_359_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_358_359_0_output_regs_ready)
		begin
			SFC_3_VALID_358_359_0_NO_SHIFT_REG <= SFC_3_VALID_357_358_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i363_stall_local;
wire [31:0] local_bb4_or_i_i363;

assign local_bb4_or_i_i363 = ((local_bb4_shl_i_i361 & 32'h1FFFFFE) | (local_bb4_shr_i_i362 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i367_stall_local;
wire [31:0] local_bb4__32_i367;

assign local_bb4__32_i367 = (local_bb4__31_i366 ? (local_bb4_shl1_i_i364 & 32'hFFFFFE00) : (local_bb4_shl1_i18_i356 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__36_i371_stall_local;
wire [31:0] local_bb4__36_i371;

assign local_bb4__36_i371 = (local_bb4__31_i366 ? (rnode_342to343_bb4_add_i357_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i537_stall_local;
wire [31:0] local_bb4__28_i537;

assign local_bb4__28_i537 = (rnode_341to342_bb4_lnot23_i517_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl66_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i526_stall_local;
wire local_bb4_lnot30_not_i526;

assign local_bb4_lnot30_not_i526 = (local_bb4_lnot30_i522 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i535_stall_local;
wire [31:0] local_bb4_shl_i535;

assign local_bb4_shl_i535 = ((local_bb4_or_i534 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_345to346_bb4_and35_i520_0_valid_out_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and35_i520_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_and35_i520_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and35_i520_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_and35_i520_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and35_i520_0_valid_out_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and35_i520_0_stall_in_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and35_i520_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_345to346_bb4_and35_i520_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to346_bb4_and35_i520_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to346_bb4_and35_i520_0_stall_in_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_345to346_bb4_and35_i520_0_valid_out_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_345to346_bb4_and35_i520_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in((rnode_343to345_bb4_and35_i520_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_345to346_bb4_and35_i520_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_345to346_bb4_and35_i520_0_reg_346_fifo.DEPTH = 1;
defparam rnode_345to346_bb4_and35_i520_0_reg_346_fifo.DATA_WIDTH = 32;
defparam rnode_345to346_bb4_and35_i520_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to346_bb4_and35_i520_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_345to346_bb4_and35_i520_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_343to345_bb4_and35_i520_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_and35_i520_0_NO_SHIFT_REG = rnode_345to346_bb4_and35_i520_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4_and35_i520_0_stall_in_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_and35_i520_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i523_stall_local;
wire local_bb4_or_cond_i523;

assign local_bb4_or_cond_i523 = (local_bb4_lnot30_i522 | local_bb4_cmp25_not_i521);

// This section implements a registered operation.
// 
wire SFC_3_VALID_359_360_0_inputs_ready;
 reg SFC_3_VALID_359_360_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_359_360_0_stall_in;
wire SFC_3_VALID_359_360_0_output_regs_ready;
 reg SFC_3_VALID_359_360_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_359_360_0_causedstall;

assign SFC_3_VALID_359_360_0_inputs_ready = 1'b1;
assign SFC_3_VALID_359_360_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_358_359_0_stall_in = 1'b0;
assign SFC_3_VALID_359_360_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_359_360_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_359_360_0_output_regs_ready)
		begin
			SFC_3_VALID_359_360_0_NO_SHIFT_REG <= SFC_3_VALID_358_359_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__34_i369_stall_local;
wire [31:0] local_bb4__34_i369;

assign local_bb4__34_i369 = (local_bb4__31_i366 ? (local_bb4_or_i_i363 & 32'h1FFFFFF) : (local_bb4_or_i17_i355 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i368_stall_local;
wire [31:0] local_bb4__33_i368;

assign local_bb4__33_i368 = (local_bb4_tobool49_i359 ? (local_bb4__32_i367 & 32'hFFFFFF00) : (local_bb4_shl1_i18_i356 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__37_i372_stall_local;
wire [31:0] local_bb4__37_i372;

assign local_bb4__37_i372 = (local_bb4_tobool49_i359 ? (local_bb4__36_i371 & 32'h1FF) : (local_bb4_inc_i360 & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb4_and73_i_stall_local;
wire [31:0] local_bb4_and73_i;

assign local_bb4_and73_i = ((local_bb4__28_i537 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and76_i_stall_local;
wire [31:0] local_bb4_and76_i;

assign local_bb4_and76_i = ((local_bb4__28_i537 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and79_i_stall_local;
wire [31:0] local_bb4_and79_i;

assign local_bb4_and79_i = ((local_bb4__28_i537 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr95_i_stall_local;
wire [31:0] local_bb4_shr95_i;

assign local_bb4_shr95_i = ((local_bb4__28_i537 & 32'h7FFFFF8) >> (local_bb4_and94_i & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and91_i_stall_local;
wire [31:0] local_bb4_and91_i;

assign local_bb4_and91_i = ((local_bb4__28_i537 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i541_stall_local;
wire [31:0] local_bb4_and88_i541;

assign local_bb4_and88_i541 = ((local_bb4__28_i537 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and85_i_stall_local;
wire [31:0] local_bb4_and85_i;

assign local_bb4_and85_i = ((local_bb4__28_i537 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u43_stall_local;
wire [31:0] local_bb4_var__u43;

assign local_bb4_var__u43 = ((local_bb4__28_i537 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i527_stall_local;
wire local_bb4_or_cond_not_i527;

assign local_bb4_or_cond_not_i527 = (local_bb4_cmp25_i518 & local_bb4_lnot30_not_i526);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i536_stall_local;
wire [31:0] local_bb4__27_i536;

assign local_bb4__27_i536 = (local_bb4_lnot_i516 ? 32'h0 : ((local_bb4_shl_i535 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i531_stall_local;
wire local_bb4_reduction_8_i531;

assign local_bb4_reduction_8_i531 = (rnode_341to343_bb4_cmp27_i519_1_NO_SHIFT_REG & local_bb4_or_cond_i523);

// This section implements a registered operation.
// 
wire SFC_3_VALID_360_361_0_inputs_ready;
 reg SFC_3_VALID_360_361_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_360_361_0_stall_in;
wire SFC_3_VALID_360_361_0_output_regs_ready;
 reg SFC_3_VALID_360_361_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_360_361_0_causedstall;

assign SFC_3_VALID_360_361_0_inputs_ready = 1'b1;
assign SFC_3_VALID_360_361_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_359_360_0_stall_in = 1'b0;
assign SFC_3_VALID_360_361_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_360_361_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_360_361_0_output_regs_ready)
		begin
			SFC_3_VALID_360_361_0_NO_SHIFT_REG <= SFC_3_VALID_359_360_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__35_i370_stall_local;
wire [31:0] local_bb4__35_i370;

assign local_bb4__35_i370 = (local_bb4_tobool49_i359 ? (local_bb4__34_i369 & 32'h1FFFFFF) : (local_bb4_or_i17_i355 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp53_i373_stall_local;
wire local_bb4_cmp53_i373;

assign local_bb4_cmp53_i373 = ((local_bb4__37_i372 & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp68_i377_stall_local;
wire local_bb4_cmp68_i377;

assign local_bb4_cmp68_i377 = ((local_bb4__37_i372 & 32'h3FF) < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i379_stall_local;
wire [31:0] local_bb4_sub_i379;

assign local_bb4_sub_i379 = ((local_bb4__37_i372 & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp71_not_i394_stall_local;
wire local_bb4_cmp71_not_i394;

assign local_bb4_cmp71_not_i394 = ((local_bb4__37_i372 & 32'h3FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4_and73_tr_i_stall_local;
wire [7:0] local_bb4_and73_tr_i;
wire [31:0] local_bb4_and73_tr_i$ps;

assign local_bb4_and73_tr_i$ps = (local_bb4_and73_i & 32'hFFFFFF);
assign local_bb4_and73_tr_i = local_bb4_and73_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i540_stall_local;
wire local_bb4_cmp77_i540;

assign local_bb4_cmp77_i540 = ((local_bb4_and76_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp80_i_stall_local;
wire local_bb4_cmp80_i;

assign local_bb4_cmp80_i = ((local_bb4_and79_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and143_i_stall_local;
wire [31:0] local_bb4_and143_i;

assign local_bb4_and143_i = (local_bb4_shr95_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr151_i_stall_local;
wire [31:0] local_bb4_shr151_i;

assign local_bb4_shr151_i = (local_bb4_shr95_i >> (local_bb4_and150_i & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u44_stall_local;
wire [31:0] local_bb4_var__u44;

assign local_bb4_var__u44 = (local_bb4_shr95_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and147_i_stall_local;
wire [31:0] local_bb4_and147_i;

assign local_bb4_and147_i = (local_bb4_shr95_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp92_i_stall_local;
wire local_bb4_cmp92_i;

assign local_bb4_cmp92_i = ((local_bb4_and91_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp89_i_stall_local;
wire local_bb4_cmp89_i;

assign local_bb4_cmp89_i = ((local_bb4_and88_i541 & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp86_i_stall_local;
wire local_bb4_cmp86_i;

assign local_bb4_cmp86_i = ((local_bb4_and85_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u45_stall_local;
wire local_bb4_var__u45;

assign local_bb4_var__u45 = ((local_bb4_var__u43 & 32'hFFF8) != 32'h0);

// This section implements a registered operation.
// 
wire SFC_3_VALID_361_362_0_inputs_ready;
 reg SFC_3_VALID_361_362_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_361_362_0_stall_in;
wire SFC_3_VALID_361_362_0_output_regs_ready;
 reg SFC_3_VALID_361_362_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_361_362_0_causedstall;

assign SFC_3_VALID_361_362_0_inputs_ready = 1'b1;
assign SFC_3_VALID_361_362_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_360_361_0_stall_in = 1'b0;
assign SFC_3_VALID_361_362_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_361_362_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_361_362_0_output_regs_ready)
		begin
			SFC_3_VALID_361_362_0_NO_SHIFT_REG <= SFC_3_VALID_360_361_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and75_i378_stall_local;
wire [31:0] local_bb4_and75_i378;

assign local_bb4_and75_i378 = ((local_bb4__35_i370 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and83_i384_stall_local;
wire [31:0] local_bb4_and83_i384;

assign local_bb4_and83_i384 = ((local_bb4__35_i370 & 32'h1FFFFFF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or581_i374_stall_local;
wire local_bb4_or581_i374;

assign local_bb4_or581_i374 = (rnode_342to343_bb4_var__u37_0_NO_SHIFT_REG | local_bb4_cmp53_i373);

// This section implements an unregistered operation.
// 
wire local_bb4_and74_i380_stall_local;
wire [31:0] local_bb4_and74_i380;

assign local_bb4_and74_i380 = ((local_bb4_sub_i379 & 32'hFF800000) + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool75_i_stall_local;
wire [7:0] local_bb4_frombool75_i;

assign local_bb4_frombool75_i = (local_bb4_and73_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u46_stall_local;
wire [31:0] local_bb4_var__u46;

assign local_bb4_var__u46 = ((local_bb4_and147_i & 32'h3FFFFFFF) | local_bb4_shr95_i);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i545_stall_local;
wire local_bb4__31_v_i545;

assign local_bb4__31_v_i545 = (local_bb4_cmp97_i ? local_bb4_cmp80_i : local_bb4_cmp92_i);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i543_stall_local;
wire local_bb4__30_v_i543;

assign local_bb4__30_v_i543 = (local_bb4_cmp97_i ? local_bb4_cmp77_i540 : local_bb4_cmp89_i);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool110_i_stall_local;
wire [7:0] local_bb4_frombool110_i;

assign local_bb4_frombool110_i[7:1] = 7'h0;
assign local_bb4_frombool110_i[0] = local_bb4_cmp86_i;

// This section implements an unregistered operation.
// 
wire local_bb4_or108_i_stall_local;
wire [31:0] local_bb4_or108_i;

assign local_bb4_or108_i[31:1] = 31'h0;
assign local_bb4_or108_i[0] = local_bb4_var__u45;

// This section implements a registered operation.
// 
wire SFC_3_VALID_362_363_0_inputs_ready;
 reg SFC_3_VALID_362_363_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_362_363_0_stall_in;
wire SFC_3_VALID_362_363_0_output_regs_ready;
 reg SFC_3_VALID_362_363_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_362_363_0_causedstall;

assign SFC_3_VALID_362_363_0_inputs_ready = 1'b1;
assign SFC_3_VALID_362_363_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_361_362_0_stall_in = 1'b0;
assign SFC_3_VALID_362_363_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_362_363_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_362_363_0_output_regs_ready)
		begin
			SFC_3_VALID_362_363_0_NO_SHIFT_REG <= SFC_3_VALID_361_362_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__33_i368_valid_out;
wire local_bb4__33_i368_stall_in;
wire local_bb4_cmp68_i377_valid_out;
wire local_bb4_cmp68_i377_stall_in;
wire local_bb4_cmp71_not_i394_valid_out;
wire local_bb4_cmp71_not_i394_stall_in;
wire local_bb4_and75_i378_valid_out;
wire local_bb4_and75_i378_stall_in;
wire local_bb4_and83_i384_valid_out;
wire local_bb4_and83_i384_stall_in;
wire local_bb4_or581_i374_valid_out;
wire local_bb4_or581_i374_stall_in;
wire local_bb4_shl_i381_valid_out;
wire local_bb4_shl_i381_stall_in;
wire local_bb4_shl_i381_inputs_ready;
wire local_bb4_shl_i381_stall_local;
wire [31:0] local_bb4_shl_i381;

assign local_bb4_shl_i381_inputs_ready = (local_bb4_mul_i_i350_valid_out_0_NO_SHIFT_REG & local_bb4_mul_i_i350_valid_out_1_NO_SHIFT_REG & rnode_342to343_bb4_add_i357_0_valid_out_1_NO_SHIFT_REG & rnode_342to343_bb4_add_i357_0_valid_out_0_NO_SHIFT_REG & rnode_342to343_bb4_add_i357_0_valid_out_2_NO_SHIFT_REG & rnode_342to343_bb4_var__u37_0_valid_out_NO_SHIFT_REG);
assign local_bb4_shl_i381 = ((local_bb4_and74_i380 & 32'hFF800000) & 32'h7F800000);
assign local_bb4__33_i368_valid_out = 1'b1;
assign local_bb4_cmp68_i377_valid_out = 1'b1;
assign local_bb4_cmp71_not_i394_valid_out = 1'b1;
assign local_bb4_and75_i378_valid_out = 1'b1;
assign local_bb4_and83_i384_valid_out = 1'b1;
assign local_bb4_or581_i374_valid_out = 1'b1;
assign local_bb4_shl_i381_valid_out = 1'b1;
assign local_bb4_mul_i_i350_stall_in_0 = 1'b0;
assign local_bb4_mul_i_i350_stall_in_1 = 1'b0;
assign rnode_342to343_bb4_add_i357_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_add_i357_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_add_i357_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_var__u37_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or1606_i_stall_local;
wire [31:0] local_bb4_or1606_i;

assign local_bb4_or1606_i = (local_bb4_var__u46 | (local_bb4_and143_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i546_stall_local;
wire [7:0] local_bb4__31_i546;

assign local_bb4__31_i546[7:1] = 7'h0;
assign local_bb4__31_i546[0] = local_bb4__31_v_i545;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i544_stall_local;
wire [7:0] local_bb4__30_i544;

assign local_bb4__30_i544[7:1] = 7'h0;
assign local_bb4__30_i544[0] = local_bb4__30_v_i543;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i542_stall_local;
wire [7:0] local_bb4__29_i542;

assign local_bb4__29_i542 = (local_bb4_cmp97_i ? (local_bb4_frombool75_i & 8'h1) : (local_bb4_frombool110_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i547_stall_local;
wire [31:0] local_bb4__32_i547;

assign local_bb4__32_i547 = (local_bb4_cmp97_i ? 32'h0 : (local_bb4_or108_i & 32'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_363_364_0_inputs_ready;
 reg SFC_3_VALID_363_364_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_363_364_0_stall_in;
wire SFC_3_VALID_363_364_0_output_regs_ready;
 reg SFC_3_VALID_363_364_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_363_364_0_causedstall;

assign SFC_3_VALID_363_364_0_inputs_ready = 1'b1;
assign SFC_3_VALID_363_364_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_362_363_0_stall_in = 1'b0;
assign SFC_3_VALID_363_364_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_363_364_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_363_364_0_output_regs_ready)
		begin
			SFC_3_VALID_363_364_0_NO_SHIFT_REG <= SFC_3_VALID_362_363_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb4__33_i368_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_343to344_bb4__33_i368_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4__33_i368_0_NO_SHIFT_REG;
 logic rnode_343to344_bb4__33_i368_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_343to344_bb4__33_i368_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4__33_i368_1_NO_SHIFT_REG;
 logic rnode_343to344_bb4__33_i368_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4__33_i368_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4__33_i368_0_valid_out_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4__33_i368_0_stall_in_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4__33_i368_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb4__33_i368_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb4__33_i368_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb4__33_i368_0_stall_in_0_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb4__33_i368_0_valid_out_0_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb4__33_i368_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in((local_bb4__33_i368 & 32'hFFFFFF00)),
	.data_out(rnode_343to344_bb4__33_i368_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb4__33_i368_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb4__33_i368_0_reg_344_fifo.DATA_WIDTH = 32;
defparam rnode_343to344_bb4__33_i368_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb4__33_i368_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb4__33_i368_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__33_i368_stall_in = 1'b0;
assign rnode_343to344_bb4__33_i368_0_stall_in_0_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb4__33_i368_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4__33_i368_0_NO_SHIFT_REG = rnode_343to344_bb4__33_i368_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb4__33_i368_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4__33_i368_1_NO_SHIFT_REG = rnode_343to344_bb4__33_i368_0_reg_344_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_cmp68_i377_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp68_i377_0_stall_in_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp68_i377_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp68_i377_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp68_i377_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp68_i377_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp68_i377_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp68_i377_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_cmp68_i377_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_cmp68_i377_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_cmp68_i377_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_cmp68_i377_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_cmp68_i377_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(local_bb4_cmp68_i377),
	.data_out(rnode_343to345_bb4_cmp68_i377_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_cmp68_i377_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_cmp68_i377_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_343to345_bb4_cmp68_i377_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_cmp68_i377_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_cmp68_i377_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp68_i377_stall_in = 1'b0;
assign rnode_343to345_bb4_cmp68_i377_0_NO_SHIFT_REG = rnode_343to345_bb4_cmp68_i377_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_cmp68_i377_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp68_i377_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_cmp71_not_i394_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp71_not_i394_0_stall_in_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp71_not_i394_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp71_not_i394_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp71_not_i394_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp71_not_i394_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp71_not_i394_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp71_not_i394_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_cmp71_not_i394_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_cmp71_not_i394_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_cmp71_not_i394_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_cmp71_not_i394_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_cmp71_not_i394_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(local_bb4_cmp71_not_i394),
	.data_out(rnode_343to345_bb4_cmp71_not_i394_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_cmp71_not_i394_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_cmp71_not_i394_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_343to345_bb4_cmp71_not_i394_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_cmp71_not_i394_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_cmp71_not_i394_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp71_not_i394_stall_in = 1'b0;
assign rnode_343to345_bb4_cmp71_not_i394_0_NO_SHIFT_REG = rnode_343to345_bb4_cmp71_not_i394_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_cmp71_not_i394_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp71_not_i394_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_and75_i378_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and75_i378_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_and75_i378_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and75_i378_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_and75_i378_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and75_i378_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and75_i378_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and75_i378_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_and75_i378_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_and75_i378_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_and75_i378_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_and75_i378_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_and75_i378_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((local_bb4_and75_i378 & 32'h7FFFFF)),
	.data_out(rnode_343to345_bb4_and75_i378_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_and75_i378_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_and75_i378_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_343to345_bb4_and75_i378_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_and75_i378_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_and75_i378_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and75_i378_stall_in = 1'b0;
assign rnode_343to345_bb4_and75_i378_0_NO_SHIFT_REG = rnode_343to345_bb4_and75_i378_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_and75_i378_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_and75_i378_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb4_and83_i384_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to344_bb4_and83_i384_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4_and83_i384_0_NO_SHIFT_REG;
 logic rnode_343to344_bb4_and83_i384_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4_and83_i384_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_and83_i384_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_and83_i384_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_and83_i384_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb4_and83_i384_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb4_and83_i384_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb4_and83_i384_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb4_and83_i384_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb4_and83_i384_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in((local_bb4_and83_i384 & 32'h1)),
	.data_out(rnode_343to344_bb4_and83_i384_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb4_and83_i384_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb4_and83_i384_0_reg_344_fifo.DATA_WIDTH = 32;
defparam rnode_343to344_bb4_and83_i384_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb4_and83_i384_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb4_and83_i384_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and83_i384_stall_in = 1'b0;
assign rnode_343to344_bb4_and83_i384_0_NO_SHIFT_REG = rnode_343to344_bb4_and83_i384_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb4_and83_i384_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb4_and83_i384_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_or581_i374_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_1_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_valid_out_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_stall_in_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_or581_i374_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_or581_i374_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_or581_i374_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_or581_i374_0_stall_in_0_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_or581_i374_0_valid_out_0_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_or581_i374_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(local_bb4_or581_i374),
	.data_out(rnode_343to345_bb4_or581_i374_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_or581_i374_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_or581_i374_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_343to345_bb4_or581_i374_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_or581_i374_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_or581_i374_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or581_i374_stall_in = 1'b0;
assign rnode_343to345_bb4_or581_i374_0_stall_in_0_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_or581_i374_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_343to345_bb4_or581_i374_0_NO_SHIFT_REG = rnode_343to345_bb4_or581_i374_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_or581_i374_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_343to345_bb4_or581_i374_1_NO_SHIFT_REG = rnode_343to345_bb4_or581_i374_0_reg_345_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_shl_i381_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shl_i381_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_shl_i381_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shl_i381_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_shl_i381_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shl_i381_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shl_i381_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_shl_i381_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_shl_i381_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_shl_i381_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_shl_i381_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_shl_i381_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_shl_i381_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((local_bb4_shl_i381 & 32'h7F800000)),
	.data_out(rnode_343to345_bb4_shl_i381_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_shl_i381_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_shl_i381_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_343to345_bb4_shl_i381_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_shl_i381_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_shl_i381_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shl_i381_stall_in = 1'b0;
assign rnode_343to345_bb4_shl_i381_0_NO_SHIFT_REG = rnode_343to345_bb4_shl_i381_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_shl_i381_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_shl_i381_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or163_i_stall_local;
wire [31:0] local_bb4_or163_i;

assign local_bb4_or163_i = (local_bb4_or1606_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1247_i_stall_local;
wire [7:0] local_bb4_or1247_i;

assign local_bb4_or1247_i = ((local_bb4__30_i544 & 8'h1) | (local_bb4__29_i542 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i549_stall_local;
wire [7:0] local_bb4__33_i549;

assign local_bb4__33_i549 = (local_bb4_cmp117_i ? (local_bb4__29_i542 & 8'h1) : (local_bb4__31_i546 & 8'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_364_365_0_inputs_ready;
 reg SFC_3_VALID_364_365_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_364_365_0_stall_in;
wire SFC_3_VALID_364_365_0_output_regs_ready;
 reg SFC_3_VALID_364_365_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_364_365_0_causedstall;

assign SFC_3_VALID_364_365_0_inputs_ready = 1'b1;
assign SFC_3_VALID_364_365_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_363_364_0_stall_in = 1'b0;
assign SFC_3_VALID_364_365_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_364_365_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_364_365_0_output_regs_ready)
		begin
			SFC_3_VALID_364_365_0_NO_SHIFT_REG <= SFC_3_VALID_363_364_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i383_stall_local;
wire local_bb4_cmp77_i383;

assign local_bb4_cmp77_i383 = ((rnode_343to344_bb4__33_i368_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u47_stall_local;
wire local_bb4_var__u47;

assign local_bb4_var__u47 = ($signed((rnode_343to344_bb4__33_i368_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u48_stall_local;
wire [31:0] local_bb4_var__u48;

assign local_bb4_var__u48[31:1] = 31'h0;
assign local_bb4_var__u48[0] = rnode_343to345_bb4_cmp68_i377_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool84_i385_stall_local;
wire local_bb4_tobool84_i385;

assign local_bb4_tobool84_i385 = ((rnode_343to344_bb4_and83_i384_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i376_stall_local;
wire local_bb4_reduction_2_i376;

assign local_bb4_reduction_2_i376 = (rnode_344to345_bb4_reduction_0_i375_0_NO_SHIFT_REG | rnode_343to345_bb4_or581_i374_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cond111_i402_stall_local;
wire [31:0] local_bb4_cond111_i402;

assign local_bb4_cond111_i402 = (rnode_343to345_bb4_or581_i374_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or76_i382_stall_local;
wire [31:0] local_bb4_or76_i382;

assign local_bb4_or76_i382 = ((rnode_343to345_bb4_shl_i381_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_343to345_bb4_and75_i378_0_NO_SHIFT_REG & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i552_stall_local;
wire [31:0] local_bb4__37_v_i552;

assign local_bb4__37_v_i552 = (local_bb4_Pivot20_i550 ? 32'h0 : (local_bb4_or163_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i548_stall_local;
wire [31:0] local_bb4_or124_i548;

assign local_bb4_or124_i548[31:8] = 24'h0;
assign local_bb4_or124_i548[7:0] = (local_bb4_or1247_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u49_stall_local;
wire [7:0] local_bb4_var__u49;

assign local_bb4_var__u49 = ((local_bb4__33_i549 & 8'h1) & 8'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_365_366_0_inputs_ready;
 reg SFC_3_VALID_365_366_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_365_366_0_stall_in;
wire SFC_3_VALID_365_366_0_output_regs_ready;
 reg SFC_3_VALID_365_366_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_365_366_0_causedstall;

assign SFC_3_VALID_365_366_0_inputs_ready = 1'b1;
assign SFC_3_VALID_365_366_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_364_365_0_stall_in = 1'b0;
assign SFC_3_VALID_365_366_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_365_366_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_365_366_0_output_regs_ready)
		begin
			SFC_3_VALID_365_366_0_NO_SHIFT_REG <= SFC_3_VALID_364_365_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__39_i386_stall_local;
wire local_bb4__39_i386;

assign local_bb4__39_i386 = (local_bb4_tobool84_i385 & local_bb4_var__u47);

// This section implements an unregistered operation.
// 
wire local_bb4_conv101_i397_stall_local;
wire [31:0] local_bb4_conv101_i397;

assign local_bb4_conv101_i397[31:1] = 31'h0;
assign local_bb4_conv101_i397[0] = local_bb4_reduction_2_i376;

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i553_stall_local;
wire [31:0] local_bb4__39_v_i553;

assign local_bb4__39_v_i553 = (local_bb4_SwitchLeaf_i551 ? (local_bb4_var__u44 & 32'h1) : (local_bb4__37_v_i552 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or125_i_stall_local;
wire [31:0] local_bb4_or125_i;

assign local_bb4_or125_i = (local_bb4_cmp117_i ? 32'h0 : (local_bb4_or124_i548 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv136_i_stall_local;
wire [31:0] local_bb4_conv136_i;

assign local_bb4_conv136_i[31:8] = 24'h0;
assign local_bb4_conv136_i[7:0] = (local_bb4_var__u49 & 8'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_366_367_0_inputs_ready;
 reg SFC_3_VALID_366_367_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_366_367_0_stall_in;
wire SFC_3_VALID_366_367_0_output_regs_ready;
 reg SFC_3_VALID_366_367_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_366_367_0_causedstall;

assign SFC_3_VALID_366_367_0_inputs_ready = 1'b1;
assign SFC_3_VALID_366_367_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_365_366_0_stall_in = 1'b0;
assign SFC_3_VALID_366_367_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_366_367_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_366_367_0_output_regs_ready)
		begin
			SFC_3_VALID_366_367_0_NO_SHIFT_REG <= SFC_3_VALID_365_366_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__40_i387_valid_out;
wire local_bb4__40_i387_stall_in;
wire local_bb4__40_i387_inputs_ready;
wire local_bb4__40_i387_stall_local;
wire local_bb4__40_i387;

assign local_bb4__40_i387_inputs_ready = (rnode_343to344_bb4__33_i368_0_valid_out_0_NO_SHIFT_REG & rnode_343to344_bb4__33_i368_0_valid_out_1_NO_SHIFT_REG & rnode_343to344_bb4_and83_i384_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40_i387 = (local_bb4_cmp77_i383 | local_bb4__39_i386);
assign local_bb4__40_i387_valid_out = 1'b1;
assign rnode_343to344_bb4__33_i368_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb4__33_i368_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb4_and83_i384_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i554_stall_local;
wire [31:0] local_bb4_reduction_3_i554;

assign local_bb4_reduction_3_i554 = ((local_bb4__32_i547 & 32'h1) | (local_bb4_or125_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or137_i_stall_local;
wire [31:0] local_bb4_or137_i;

assign local_bb4_or137_i = (local_bb4_cmp132_not_i ? (local_bb4_conv136_i & 32'h1) : 32'h0);

// This section implements a registered operation.
// 
wire SFC_3_VALID_367_368_0_inputs_ready;
 reg SFC_3_VALID_367_368_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_367_368_0_stall_in;
wire SFC_3_VALID_367_368_0_output_regs_ready;
 reg SFC_3_VALID_367_368_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_367_368_0_causedstall;

assign SFC_3_VALID_367_368_0_inputs_ready = 1'b1;
assign SFC_3_VALID_367_368_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_366_367_0_stall_in = 1'b0;
assign SFC_3_VALID_367_368_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_367_368_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_367_368_0_output_regs_ready)
		begin
			SFC_3_VALID_367_368_0_NO_SHIFT_REG <= SFC_3_VALID_366_367_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4__40_i387_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb4__40_i387_0_stall_in_NO_SHIFT_REG;
 logic rnode_344to345_bb4__40_i387_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4__40_i387_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_344to345_bb4__40_i387_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__40_i387_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__40_i387_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__40_i387_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4__40_i387_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4__40_i387_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4__40_i387_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4__40_i387_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4__40_i387_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(local_bb4__40_i387),
	.data_out(rnode_344to345_bb4__40_i387_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4__40_i387_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4__40_i387_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_344to345_bb4__40_i387_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4__40_i387_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4__40_i387_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_i387_stall_in = 1'b0;
assign rnode_344to345_bb4__40_i387_0_NO_SHIFT_REG = rnode_344to345_bb4__40_i387_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4__40_i387_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__40_i387_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i556_stall_local;
wire [31:0] local_bb4_reduction_5_i556;

assign local_bb4_reduction_5_i556 = (local_bb4_shr151_i | (local_bb4_reduction_3_i554 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i555_stall_local;
wire [31:0] local_bb4_reduction_4_i555;

assign local_bb4_reduction_4_i555 = ((local_bb4_or137_i & 32'h1) | (local_bb4__39_v_i553 & 32'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_368_369_0_inputs_ready;
 reg SFC_3_VALID_368_369_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_368_369_0_stall_in;
wire SFC_3_VALID_368_369_0_output_regs_ready;
 reg SFC_3_VALID_368_369_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_368_369_0_causedstall;

assign SFC_3_VALID_368_369_0_inputs_ready = 1'b1;
assign SFC_3_VALID_368_369_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_367_368_0_stall_in = 1'b0;
assign SFC_3_VALID_368_369_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_368_369_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_368_369_0_output_regs_ready)
		begin
			SFC_3_VALID_368_369_0_NO_SHIFT_REG <= SFC_3_VALID_367_368_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_cond_i388_stall_local;
wire [31:0] local_bb4_cond_i388;

assign local_bb4_cond_i388[31:1] = 31'h0;
assign local_bb4_cond_i388[0] = rnode_344to345_bb4__40_i387_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i557_stall_local;
wire [31:0] local_bb4_reduction_6_i557;

assign local_bb4_reduction_6_i557 = ((local_bb4_reduction_4_i555 & 32'h1) | local_bb4_reduction_5_i556);

// This section implements a registered operation.
// 
wire SFC_3_VALID_369_370_0_inputs_ready;
 reg SFC_3_VALID_369_370_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_369_370_0_stall_in;
wire SFC_3_VALID_369_370_0_output_regs_ready;
 reg SFC_3_VALID_369_370_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_369_370_0_causedstall;

assign SFC_3_VALID_369_370_0_inputs_ready = 1'b1;
assign SFC_3_VALID_369_370_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_368_369_0_stall_in = 1'b0;
assign SFC_3_VALID_369_370_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_369_370_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_369_370_0_output_regs_ready)
		begin
			SFC_3_VALID_369_370_0_NO_SHIFT_REG <= SFC_3_VALID_368_369_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_add87_i389_stall_local;
wire [31:0] local_bb4_add87_i389;

assign local_bb4_add87_i389 = ((local_bb4_cond_i388 & 32'h1) + (local_bb4_or76_i382 & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i524_valid_out;
wire local_bb4_lnot33_not_i524_stall_in;
wire local_bb4_cmp38_i_valid_out;
wire local_bb4_cmp38_i_stall_in;
wire local_bb4_and37_lobit_i_valid_out;
wire local_bb4_and37_lobit_i_stall_in;
wire local_bb4_xor189_i_valid_out;
wire local_bb4_xor189_i_stall_in;
wire local_bb4_xor189_i_inputs_ready;
wire local_bb4_xor189_i_stall_local;
wire [31:0] local_bb4_xor189_i;

assign local_bb4_xor189_i_inputs_ready = (rnode_341to342_bb4__22_i508_0_valid_out_0_NO_SHIFT_REG & rnode_341to342_bb4_lnot23_i517_0_valid_out_NO_SHIFT_REG & rnode_341to342_bb4_align_0_i539_0_valid_out_0_NO_SHIFT_REG & rnode_341to342_bb4_align_0_i539_0_valid_out_4_NO_SHIFT_REG & rnode_341to342_bb4_align_0_i539_0_valid_out_1_NO_SHIFT_REG & rnode_341to342_bb4_align_0_i539_0_valid_out_2_NO_SHIFT_REG & rnode_341to342_bb4_align_0_i539_0_valid_out_3_NO_SHIFT_REG & rnode_341to342_bb4__23_i509_0_valid_out_2_NO_SHIFT_REG & rnode_341to342_bb4__22_i508_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor189_i = (local_bb4_reduction_6_i557 ^ local_bb4_xor36_lobit_i);
assign local_bb4_lnot33_not_i524_valid_out = 1'b1;
assign local_bb4_cmp38_i_valid_out = 1'b1;
assign local_bb4_and37_lobit_i_valid_out = 1'b1;
assign local_bb4_xor189_i_valid_out = 1'b1;
assign rnode_341to342_bb4__22_i508_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_lnot23_i517_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_align_0_i539_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_align_0_i539_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_align_0_i539_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_align_0_i539_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4_align_0_i539_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4__23_i509_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_341to342_bb4__22_i508_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_370_371_0_inputs_ready;
 reg SFC_3_VALID_370_371_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_370_371_0_stall_in;
wire SFC_3_VALID_370_371_0_output_regs_ready;
 reg SFC_3_VALID_370_371_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_370_371_0_causedstall;

assign SFC_3_VALID_370_371_0_inputs_ready = 1'b1;
assign SFC_3_VALID_370_371_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_369_370_0_stall_in = 1'b0;
assign SFC_3_VALID_370_371_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_370_371_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_370_371_0_output_regs_ready)
		begin
			SFC_3_VALID_370_371_0_NO_SHIFT_REG <= SFC_3_VALID_369_370_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and88_i390_stall_local;
wire [31:0] local_bb4_and88_i390;

assign local_bb4_and88_i390 = (local_bb4_add87_i389 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i392_stall_local;
wire [31:0] local_bb4_and90_i392;

assign local_bb4_and90_i392 = (local_bb4_add87_i389 & 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_lnot33_not_i524_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb4_lnot33_not_i524_0_stall_in_NO_SHIFT_REG;
 logic rnode_342to343_bb4_lnot33_not_i524_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_lnot33_not_i524_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic rnode_342to343_bb4_lnot33_not_i524_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_lnot33_not_i524_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_lnot33_not_i524_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_lnot33_not_i524_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_lnot33_not_i524_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_lnot33_not_i524_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_lnot33_not_i524_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_lnot33_not_i524_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_lnot33_not_i524_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i524),
	.data_out(rnode_342to343_bb4_lnot33_not_i524_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_lnot33_not_i524_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_lnot33_not_i524_0_reg_343_fifo.DATA_WIDTH = 1;
defparam rnode_342to343_bb4_lnot33_not_i524_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_lnot33_not_i524_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_lnot33_not_i524_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i524_stall_in = 1'b0;
assign rnode_342to343_bb4_lnot33_not_i524_0_NO_SHIFT_REG = rnode_342to343_bb4_lnot33_not_i524_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_lnot33_not_i524_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_lnot33_not_i524_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_valid_out_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_stall_in_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_cmp38_i_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_cmp38_i_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_cmp38_i_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_cmp38_i_0_stall_in_0_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_cmp38_i_0_valid_out_0_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_cmp38_i_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in(local_bb4_cmp38_i),
	.data_out(rnode_342to343_bb4_cmp38_i_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_cmp38_i_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_cmp38_i_0_reg_343_fifo.DATA_WIDTH = 1;
defparam rnode_342to343_bb4_cmp38_i_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_cmp38_i_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_cmp38_i_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp38_i_stall_in = 1'b0;
assign rnode_342to343_bb4_cmp38_i_0_stall_in_0_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_cmp38_i_0_NO_SHIFT_REG = rnode_342to343_bb4_cmp38_i_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_cmp38_i_1_NO_SHIFT_REG = rnode_342to343_bb4_cmp38_i_0_reg_343_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and37_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_and37_lobit_i_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and37_lobit_i_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_and37_lobit_i_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and37_lobit_i_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and37_lobit_i_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_and37_lobit_i_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_and37_lobit_i_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_and37_lobit_i_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_and37_lobit_i_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_and37_lobit_i_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_and37_lobit_i_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in((local_bb4_and37_lobit_i & 32'h1)),
	.data_out(rnode_342to343_bb4_and37_lobit_i_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_and37_lobit_i_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_and37_lobit_i_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb4_and37_lobit_i_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_and37_lobit_i_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_and37_lobit_i_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and37_lobit_i_stall_in = 1'b0;
assign rnode_342to343_bb4_and37_lobit_i_0_NO_SHIFT_REG = rnode_342to343_bb4_and37_lobit_i_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_and37_lobit_i_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_342to343_bb4_xor189_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_342to343_bb4_xor189_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_xor189_i_0_NO_SHIFT_REG;
 logic rnode_342to343_bb4_xor189_i_0_reg_343_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_342to343_bb4_xor189_i_0_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_xor189_i_0_valid_out_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_xor189_i_0_stall_in_reg_343_NO_SHIFT_REG;
 logic rnode_342to343_bb4_xor189_i_0_stall_out_reg_343_NO_SHIFT_REG;

acl_data_fifo rnode_342to343_bb4_xor189_i_0_reg_343_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_342to343_bb4_xor189_i_0_reg_343_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_342to343_bb4_xor189_i_0_stall_in_reg_343_NO_SHIFT_REG),
	.valid_out(rnode_342to343_bb4_xor189_i_0_valid_out_reg_343_NO_SHIFT_REG),
	.stall_out(rnode_342to343_bb4_xor189_i_0_stall_out_reg_343_NO_SHIFT_REG),
	.data_in(local_bb4_xor189_i),
	.data_out(rnode_342to343_bb4_xor189_i_0_reg_343_NO_SHIFT_REG)
);

defparam rnode_342to343_bb4_xor189_i_0_reg_343_fifo.DEPTH = 1;
defparam rnode_342to343_bb4_xor189_i_0_reg_343_fifo.DATA_WIDTH = 32;
defparam rnode_342to343_bb4_xor189_i_0_reg_343_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_342to343_bb4_xor189_i_0_reg_343_fifo.IMPL = "shift_reg";

assign rnode_342to343_bb4_xor189_i_0_reg_343_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor189_i_stall_in = 1'b0;
assign rnode_342to343_bb4_xor189_i_0_NO_SHIFT_REG = rnode_342to343_bb4_xor189_i_0_reg_343_NO_SHIFT_REG;
assign rnode_342to343_bb4_xor189_i_0_stall_in_reg_343_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_xor189_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_371_372_0_inputs_ready;
 reg SFC_3_VALID_371_372_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_371_372_0_stall_in;
wire SFC_3_VALID_371_372_0_output_regs_ready;
 reg SFC_3_VALID_371_372_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_371_372_0_causedstall;

assign SFC_3_VALID_371_372_0_inputs_ready = 1'b1;
assign SFC_3_VALID_371_372_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_370_371_0_stall_in = 1'b0;
assign SFC_3_VALID_371_372_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_371_372_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_371_372_0_output_regs_ready)
		begin
			SFC_3_VALID_371_372_0_NO_SHIFT_REG <= SFC_3_VALID_370_371_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or89_i391_stall_local;
wire [31:0] local_bb4_or89_i391;

assign local_bb4_or89_i391 = ((local_bb4_and88_i390 & 32'h7FFFFFFF) | (local_bb4_and4_i317 & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i393_stall_local;
wire local_bb4_cmp91_i393;

assign local_bb4_cmp91_i393 = ((local_bb4_and90_i392 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i525_stall_local;
wire local_bb4_brmerge_not_i525;

assign local_bb4_brmerge_not_i525 = (rnode_341to343_bb4_cmp27_i519_0_NO_SHIFT_REG & rnode_342to343_bb4_lnot33_not_i524_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_2_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_valid_out_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_stall_in_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_cmp38_i_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_cmp38_i_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_cmp38_i_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_cmp38_i_0_stall_in_0_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_cmp38_i_0_valid_out_0_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_cmp38_i_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(rnode_342to343_bb4_cmp38_i_1_NO_SHIFT_REG),
	.data_out(rnode_343to345_bb4_cmp38_i_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_cmp38_i_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_cmp38_i_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_343to345_bb4_cmp38_i_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_cmp38_i_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_cmp38_i_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_342to343_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp38_i_0_stall_in_0_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_343to345_bb4_cmp38_i_0_NO_SHIFT_REG = rnode_343to345_bb4_cmp38_i_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_343to345_bb4_cmp38_i_1_NO_SHIFT_REG = rnode_343to345_bb4_cmp38_i_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_343to345_bb4_cmp38_i_2_NO_SHIFT_REG = rnode_343to345_bb4_cmp38_i_0_reg_345_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i558_stall_local;
wire [31:0] local_bb4_add_i558;

assign local_bb4_add_i558 = ((local_bb4__27_i536 & 32'h7FFFFF8) | (rnode_342to343_bb4_and37_lobit_i_0_NO_SHIFT_REG & 32'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_372_373_0_inputs_ready;
 reg SFC_3_VALID_372_373_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_372_373_0_stall_in;
wire SFC_3_VALID_372_373_0_output_regs_ready;
 reg SFC_3_VALID_372_373_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_372_373_0_causedstall;

assign SFC_3_VALID_372_373_0_inputs_ready = 1'b1;
assign SFC_3_VALID_372_373_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_371_372_0_stall_in = 1'b0;
assign SFC_3_VALID_372_373_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_372_373_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_372_373_0_output_regs_ready)
		begin
			SFC_3_VALID_372_373_0_NO_SHIFT_REG <= SFC_3_VALID_371_372_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_brmerge14_i395_stall_local;
wire local_bb4_brmerge14_i395;

assign local_bb4_brmerge14_i395 = (local_bb4_cmp91_i393 | rnode_343to345_bb4_cmp71_not_i394_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i528_stall_local;
wire local_bb4__24_i528;

assign local_bb4__24_i528 = (local_bb4_or_cond_not_i527 | local_bb4_brmerge_not_i525);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i529_stall_local;
wire local_bb4_brmerge_not_not_i529;

assign local_bb4_brmerge_not_not_i529 = (local_bb4_brmerge_not_i525 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp38_i_stall_local;
wire local_bb4_not_cmp38_i;

assign local_bb4_not_cmp38_i = (rnode_343to345_bb4_cmp38_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add193_i_stall_local;
wire [31:0] local_bb4_add193_i;

assign local_bb4_add193_i = ((local_bb4_add_i558 & 32'h7FFFFF9) + rnode_342to343_bb4_xor189_i_0_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_3_VALID_373_374_0_inputs_ready;
 reg SFC_3_VALID_373_374_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_373_374_0_stall_in;
wire SFC_3_VALID_373_374_0_output_regs_ready;
 reg SFC_3_VALID_373_374_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_373_374_0_causedstall;

assign SFC_3_VALID_373_374_0_inputs_ready = 1'b1;
assign SFC_3_VALID_373_374_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_372_373_0_stall_in = 1'b0;
assign SFC_3_VALID_373_374_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_373_374_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_373_374_0_output_regs_ready)
		begin
			SFC_3_VALID_373_374_0_NO_SHIFT_REG <= SFC_3_VALID_372_373_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_conv99_i396_stall_local;
wire [31:0] local_bb4_conv99_i396;

assign local_bb4_conv99_i396 = (local_bb4_brmerge14_i395 ? (local_bb4_var__u48 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i530_stall_local;
wire local_bb4_reduction_7_i530;

assign local_bb4_reduction_7_i530 = (local_bb4_cmp25_i518 & local_bb4_brmerge_not_not_i529);

// This section implements a registered operation.
// 
wire SFC_3_VALID_374_375_0_inputs_ready;
 reg SFC_3_VALID_374_375_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_374_375_0_stall_in;
wire SFC_3_VALID_374_375_0_output_regs_ready;
 reg SFC_3_VALID_374_375_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_374_375_0_causedstall;

assign SFC_3_VALID_374_375_0_inputs_ready = 1'b1;
assign SFC_3_VALID_374_375_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_373_374_0_stall_in = 1'b0;
assign SFC_3_VALID_374_375_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_374_375_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_374_375_0_output_regs_ready)
		begin
			SFC_3_VALID_374_375_0_NO_SHIFT_REG <= SFC_3_VALID_373_374_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or102_i398_stall_local;
wire [31:0] local_bb4_or102_i398;

assign local_bb4_or102_i398 = ((local_bb4_conv99_i396 & 32'h1) | (local_bb4_conv101_i397 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i532_stall_local;
wire local_bb4_reduction_9_i532;

assign local_bb4_reduction_9_i532 = (local_bb4_reduction_7_i530 & local_bb4_reduction_8_i531);

// This section implements a registered operation.
// 
wire SFC_3_VALID_375_376_0_inputs_ready;
 reg SFC_3_VALID_375_376_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_375_376_0_stall_in;
wire SFC_3_VALID_375_376_0_output_regs_ready;
 reg SFC_3_VALID_375_376_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_375_376_0_causedstall;

assign SFC_3_VALID_375_376_0_inputs_ready = 1'b1;
assign SFC_3_VALID_375_376_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_374_375_0_stall_in = 1'b0;
assign SFC_3_VALID_375_376_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_375_376_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_375_376_0_output_regs_ready)
		begin
			SFC_3_VALID_375_376_0_NO_SHIFT_REG <= SFC_3_VALID_374_375_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_tobool103_i399_stall_local;
wire local_bb4_tobool103_i399;

assign local_bb4_tobool103_i399 = ((local_bb4_or102_i398 & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i511_valid_out_2;
wire local_bb4_and17_i511_stall_in_2;
wire local_bb4_var__u42_valid_out;
wire local_bb4_var__u42_stall_in;
wire local_bb4_add193_i_valid_out;
wire local_bb4_add193_i_stall_in;
wire local_bb4__26_i533_valid_out;
wire local_bb4__26_i533_stall_in;
wire local_bb4__26_i533_inputs_ready;
wire local_bb4__26_i533_stall_local;
wire local_bb4__26_i533;

assign local_bb4__26_i533_inputs_ready = (rnode_341to343_bb4_shr16_i510_0_valid_out_0_NO_SHIFT_REG & rnode_341to343_bb4_cmp27_i519_0_valid_out_2_NO_SHIFT_REG & rnode_342to343_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_342to343_bb4_xor189_i_0_valid_out_NO_SHIFT_REG & rnode_342to343_bb4_and20_i514_0_valid_out_0_NO_SHIFT_REG & rnode_341to343_bb4_cmp27_i519_0_valid_out_0_NO_SHIFT_REG & rnode_342to343_bb4_lnot33_not_i524_0_valid_out_NO_SHIFT_REG & rnode_341to343_bb4_cmp27_i519_0_valid_out_1_NO_SHIFT_REG & rnode_342to343_bb4_and20_i514_0_valid_out_1_NO_SHIFT_REG & rnode_342to343_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i533 = (local_bb4_reduction_9_i532 ? rnode_342to343_bb4_cmp38_i_0_NO_SHIFT_REG : local_bb4__24_i528);
assign local_bb4_and17_i511_valid_out_2 = 1'b1;
assign local_bb4_var__u42_valid_out = 1'b1;
assign local_bb4_add193_i_valid_out = 1'b1;
assign local_bb4__26_i533_valid_out = 1'b1;
assign rnode_341to343_bb4_shr16_i510_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_341to343_bb4_cmp27_i519_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_and37_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_xor189_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_and20_i514_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_341to343_bb4_cmp27_i519_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_lnot33_not_i524_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_341to343_bb4_cmp27_i519_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_and20_i514_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_342to343_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_376_377_0_inputs_ready;
 reg SFC_3_VALID_376_377_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_376_377_0_stall_in;
wire SFC_3_VALID_376_377_0_output_regs_ready;
 reg SFC_3_VALID_376_377_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_376_377_0_causedstall;

assign SFC_3_VALID_376_377_0_inputs_ready = 1'b1;
assign SFC_3_VALID_376_377_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_375_376_0_stall_in = 1'b0;
assign SFC_3_VALID_376_377_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_376_377_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_376_377_0_output_regs_ready)
		begin
			SFC_3_VALID_376_377_0_NO_SHIFT_REG <= SFC_3_VALID_375_376_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_cond107_i400_stall_local;
wire [31:0] local_bb4_cond107_i400;

assign local_bb4_cond107_i400 = (local_bb4_tobool103_i399 ? (local_bb4_and4_i317 & 32'h80000000) : 32'hFFFFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_343to345_bb4_and17_i511_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and17_i511_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_and17_i511_0_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and17_i511_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to345_bb4_and17_i511_0_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and17_i511_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and17_i511_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_343to345_bb4_and17_i511_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_343to345_bb4_and17_i511_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to345_bb4_and17_i511_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to345_bb4_and17_i511_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_343to345_bb4_and17_i511_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_343to345_bb4_and17_i511_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i511 & 32'hFF)),
	.data_out(rnode_343to345_bb4_and17_i511_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_343to345_bb4_and17_i511_0_reg_345_fifo.DEPTH = 2;
defparam rnode_343to345_bb4_and17_i511_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_343to345_bb4_and17_i511_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to345_bb4_and17_i511_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_343to345_bb4_and17_i511_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i511_stall_in_2 = 1'b0;
assign rnode_343to345_bb4_and17_i511_0_NO_SHIFT_REG = rnode_343to345_bb4_and17_i511_0_reg_345_NO_SHIFT_REG;
assign rnode_343to345_bb4_and17_i511_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_and17_i511_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb4_var__u42_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to344_bb4_var__u42_0_stall_in_NO_SHIFT_REG;
 logic rnode_343to344_bb4_var__u42_0_NO_SHIFT_REG;
 logic rnode_343to344_bb4_var__u42_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to344_bb4_var__u42_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_var__u42_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_var__u42_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_var__u42_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb4_var__u42_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb4_var__u42_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb4_var__u42_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb4_var__u42_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb4_var__u42_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(local_bb4_var__u42),
	.data_out(rnode_343to344_bb4_var__u42_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb4_var__u42_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb4_var__u42_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_343to344_bb4_var__u42_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb4_var__u42_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb4_var__u42_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u42_stall_in = 1'b0;
assign rnode_343to344_bb4_var__u42_0_NO_SHIFT_REG = rnode_343to344_bb4_var__u42_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb4_var__u42_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb4_var__u42_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4_add193_i_0_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4_add193_i_1_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4_add193_i_2_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4_add193_i_3_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_343to344_bb4_add193_i_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_valid_out_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_stall_in_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4_add193_i_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb4_add193_i_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb4_add193_i_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb4_add193_i_0_stall_in_0_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb4_add193_i_0_valid_out_0_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb4_add193_i_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(local_bb4_add193_i),
	.data_out(rnode_343to344_bb4_add193_i_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb4_add193_i_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb4_add193_i_0_reg_344_fifo.DATA_WIDTH = 32;
defparam rnode_343to344_bb4_add193_i_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb4_add193_i_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb4_add193_i_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add193_i_stall_in = 1'b0;
assign rnode_343to344_bb4_add193_i_0_stall_in_0_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4_add193_i_0_NO_SHIFT_REG = rnode_343to344_bb4_add193_i_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4_add193_i_1_NO_SHIFT_REG = rnode_343to344_bb4_add193_i_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4_add193_i_2_NO_SHIFT_REG = rnode_343to344_bb4_add193_i_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4_add193_i_3_NO_SHIFT_REG = rnode_343to344_bb4_add193_i_0_reg_344_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_343to344_bb4__26_i533_0_valid_out_NO_SHIFT_REG;
 logic rnode_343to344_bb4__26_i533_0_stall_in_NO_SHIFT_REG;
 logic rnode_343to344_bb4__26_i533_0_NO_SHIFT_REG;
 logic rnode_343to344_bb4__26_i533_0_reg_344_inputs_ready_NO_SHIFT_REG;
 logic rnode_343to344_bb4__26_i533_0_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4__26_i533_0_valid_out_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4__26_i533_0_stall_in_reg_344_NO_SHIFT_REG;
 logic rnode_343to344_bb4__26_i533_0_stall_out_reg_344_NO_SHIFT_REG;

acl_data_fifo rnode_343to344_bb4__26_i533_0_reg_344_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_343to344_bb4__26_i533_0_reg_344_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_343to344_bb4__26_i533_0_stall_in_reg_344_NO_SHIFT_REG),
	.valid_out(rnode_343to344_bb4__26_i533_0_valid_out_reg_344_NO_SHIFT_REG),
	.stall_out(rnode_343to344_bb4__26_i533_0_stall_out_reg_344_NO_SHIFT_REG),
	.data_in(local_bb4__26_i533),
	.data_out(rnode_343to344_bb4__26_i533_0_reg_344_NO_SHIFT_REG)
);

defparam rnode_343to344_bb4__26_i533_0_reg_344_fifo.DEPTH = 1;
defparam rnode_343to344_bb4__26_i533_0_reg_344_fifo.DATA_WIDTH = 1;
defparam rnode_343to344_bb4__26_i533_0_reg_344_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_343to344_bb4__26_i533_0_reg_344_fifo.IMPL = "shift_reg";

assign rnode_343to344_bb4__26_i533_0_reg_344_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i533_stall_in = 1'b0;
assign rnode_343to344_bb4__26_i533_0_NO_SHIFT_REG = rnode_343to344_bb4__26_i533_0_reg_344_NO_SHIFT_REG;
assign rnode_343to344_bb4__26_i533_0_stall_in_reg_344_NO_SHIFT_REG = 1'b0;
assign rnode_343to344_bb4__26_i533_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_377_378_0_inputs_ready;
 reg SFC_3_VALID_377_378_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_377_378_0_stall_in;
wire SFC_3_VALID_377_378_0_output_regs_ready;
 reg SFC_3_VALID_377_378_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_377_378_0_causedstall;

assign SFC_3_VALID_377_378_0_inputs_ready = 1'b1;
assign SFC_3_VALID_377_378_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_376_377_0_stall_in = 1'b0;
assign SFC_3_VALID_377_378_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_377_378_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_377_378_0_output_regs_ready)
		begin
			SFC_3_VALID_377_378_0_NO_SHIFT_REG <= SFC_3_VALID_376_377_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and108_i401_stall_local;
wire [31:0] local_bb4_and108_i401;

assign local_bb4_and108_i401 = (local_bb4_cond107_i400 & local_bb4_or89_i391);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4_var__u42_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb4_var__u42_0_stall_in_NO_SHIFT_REG;
 logic rnode_344to345_bb4_var__u42_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4_var__u42_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic rnode_344to345_bb4_var__u42_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_var__u42_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_var__u42_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_var__u42_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4_var__u42_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4_var__u42_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4_var__u42_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4_var__u42_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4_var__u42_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in(rnode_343to344_bb4_var__u42_0_NO_SHIFT_REG),
	.data_out(rnode_344to345_bb4_var__u42_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4_var__u42_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4_var__u42_0_reg_345_fifo.DATA_WIDTH = 1;
defparam rnode_344to345_bb4_var__u42_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4_var__u42_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4_var__u42_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4_var__u42_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_var__u42_0_NO_SHIFT_REG = rnode_344to345_bb4_var__u42_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4_var__u42_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_var__u42_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and194_i_valid_out;
wire local_bb4_and194_i_stall_in;
wire local_bb4_and194_i_inputs_ready;
wire local_bb4_and194_i_stall_local;
wire [31:0] local_bb4_and194_i;

assign local_bb4_and194_i_inputs_ready = rnode_343to344_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and194_i = (rnode_343to344_bb4_add193_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and194_i_valid_out = 1'b1;
assign rnode_343to344_bb4_add193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and196_i_valid_out;
wire local_bb4_and196_i_stall_in;
wire local_bb4_and196_i_inputs_ready;
wire local_bb4_and196_i_stall_local;
wire [31:0] local_bb4_and196_i;

assign local_bb4_and196_i_inputs_ready = rnode_343to344_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and196_i = (rnode_343to344_bb4_add193_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and196_i_valid_out = 1'b1;
assign rnode_343to344_bb4_add193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and199_i_valid_out;
wire local_bb4_and199_i_stall_in;
wire local_bb4_and199_i_inputs_ready;
wire local_bb4_and199_i_stall_local;
wire [31:0] local_bb4_and199_i;

assign local_bb4_and199_i_inputs_ready = rnode_343to344_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and199_i = (rnode_343to344_bb4_add193_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and199_i_valid_out = 1'b1;
assign rnode_343to344_bb4_add193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and202_i_stall_local;
wire [31:0] local_bb4_and202_i;

assign local_bb4_and202_i = (rnode_343to344_bb4_add193_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_344to346_bb4__26_i533_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to346_bb4__26_i533_0_stall_in_NO_SHIFT_REG;
 logic rnode_344to346_bb4__26_i533_0_NO_SHIFT_REG;
 logic rnode_344to346_bb4__26_i533_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic rnode_344to346_bb4__26_i533_0_reg_346_NO_SHIFT_REG;
 logic rnode_344to346_bb4__26_i533_0_valid_out_reg_346_NO_SHIFT_REG;
 logic rnode_344to346_bb4__26_i533_0_stall_in_reg_346_NO_SHIFT_REG;
 logic rnode_344to346_bb4__26_i533_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_344to346_bb4__26_i533_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to346_bb4__26_i533_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to346_bb4__26_i533_0_stall_in_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_344to346_bb4__26_i533_0_valid_out_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_344to346_bb4__26_i533_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in(rnode_343to344_bb4__26_i533_0_NO_SHIFT_REG),
	.data_out(rnode_344to346_bb4__26_i533_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_344to346_bb4__26_i533_0_reg_346_fifo.DEPTH = 2;
defparam rnode_344to346_bb4__26_i533_0_reg_346_fifo.DATA_WIDTH = 1;
defparam rnode_344to346_bb4__26_i533_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to346_bb4__26_i533_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_344to346_bb4__26_i533_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_343to344_bb4__26_i533_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to346_bb4__26_i533_0_NO_SHIFT_REG = rnode_344to346_bb4__26_i533_0_reg_346_NO_SHIFT_REG;
assign rnode_344to346_bb4__26_i533_0_stall_in_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_344to346_bb4__26_i533_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_378_379_0_inputs_ready;
 reg SFC_3_VALID_378_379_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_378_379_0_stall_in;
wire SFC_3_VALID_378_379_0_output_regs_ready;
 reg SFC_3_VALID_378_379_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_378_379_0_causedstall;

assign SFC_3_VALID_378_379_0_inputs_ready = 1'b1;
assign SFC_3_VALID_378_379_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_377_378_0_stall_in = 1'b0;
assign SFC_3_VALID_378_379_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_378_379_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_378_379_0_output_regs_ready)
		begin
			SFC_3_VALID_378_379_0_NO_SHIFT_REG <= SFC_3_VALID_377_378_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or112_i403_stall_local;
wire [31:0] local_bb4_or112_i403;

assign local_bb4_or112_i403 = (local_bb4_and108_i401 | (local_bb4_cond111_i402 & 32'h7F800000));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_345to346_bb4_var__u42_0_valid_out_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u42_0_stall_in_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u42_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u42_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u42_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u42_0_valid_out_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u42_0_stall_in_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u42_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_345to346_bb4_var__u42_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to346_bb4_var__u42_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to346_bb4_var__u42_0_stall_in_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_345to346_bb4_var__u42_0_valid_out_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_345to346_bb4_var__u42_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in(rnode_344to345_bb4_var__u42_0_NO_SHIFT_REG),
	.data_out(rnode_345to346_bb4_var__u42_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_345to346_bb4_var__u42_0_reg_346_fifo.DEPTH = 1;
defparam rnode_345to346_bb4_var__u42_0_reg_346_fifo.DATA_WIDTH = 1;
defparam rnode_345to346_bb4_var__u42_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to346_bb4_var__u42_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_345to346_bb4_var__u42_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_344to345_bb4_var__u42_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_var__u42_0_NO_SHIFT_REG = rnode_345to346_bb4_var__u42_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4_var__u42_0_stall_in_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_var__u42_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and194_i_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and194_i_1_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and194_i_2_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and194_i_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_valid_out_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_stall_in_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and194_i_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4_and194_i_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4_and194_i_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4_and194_i_0_stall_in_0_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4_and194_i_0_valid_out_0_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4_and194_i_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((local_bb4_and194_i & 32'hFFFFFFF)),
	.data_out(rnode_344to345_bb4_and194_i_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4_and194_i_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4_and194_i_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_344to345_bb4_and194_i_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4_and194_i_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4_and194_i_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and194_i_stall_in = 1'b0;
assign rnode_344to345_bb4_and194_i_0_stall_in_0_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_344to345_bb4_and194_i_0_NO_SHIFT_REG = rnode_344to345_bb4_and194_i_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_344to345_bb4_and194_i_1_NO_SHIFT_REG = rnode_344to345_bb4_and194_i_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_344to345_bb4_and194_i_2_NO_SHIFT_REG = rnode_344to345_bb4_and194_i_0_reg_345_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4_and196_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and196_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and196_i_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and196_i_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and196_i_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and196_i_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and196_i_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and196_i_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4_and196_i_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4_and196_i_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4_and196_i_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4_and196_i_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4_and196_i_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((local_bb4_and196_i & 32'h1F)),
	.data_out(rnode_344to345_bb4_and196_i_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4_and196_i_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4_and196_i_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_344to345_bb4_and196_i_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4_and196_i_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4_and196_i_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and196_i_stall_in = 1'b0;
assign rnode_344to345_bb4_and196_i_0_NO_SHIFT_REG = rnode_344to345_bb4_and196_i_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4_and196_i_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and196_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4_and199_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and199_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and199_i_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and199_i_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4_and199_i_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and199_i_0_valid_out_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and199_i_0_stall_in_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4_and199_i_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4_and199_i_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4_and199_i_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4_and199_i_0_stall_in_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4_and199_i_0_valid_out_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4_and199_i_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((local_bb4_and199_i & 32'h1)),
	.data_out(rnode_344to345_bb4_and199_i_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4_and199_i_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4_and199_i_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_344to345_bb4_and199_i_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4_and199_i_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4_and199_i_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and199_i_stall_in = 1'b0;
assign rnode_344to345_bb4_and199_i_0_NO_SHIFT_REG = rnode_344to345_bb4_and199_i_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4_and199_i_0_stall_in_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and199_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i559_stall_local;
wire [31:0] local_bb4_shr_i_i559;

assign local_bb4_shr_i_i559 = ((local_bb4_and202_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_346to347_bb4__26_i533_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_2_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_valid_out_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_stall_in_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4__26_i533_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_346to347_bb4__26_i533_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to347_bb4__26_i533_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to347_bb4__26_i533_0_stall_in_0_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_346to347_bb4__26_i533_0_valid_out_0_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_346to347_bb4__26_i533_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in(rnode_344to346_bb4__26_i533_0_NO_SHIFT_REG),
	.data_out(rnode_346to347_bb4__26_i533_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_346to347_bb4__26_i533_0_reg_347_fifo.DEPTH = 1;
defparam rnode_346to347_bb4__26_i533_0_reg_347_fifo.DATA_WIDTH = 1;
defparam rnode_346to347_bb4__26_i533_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to347_bb4__26_i533_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_346to347_bb4__26_i533_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_344to346_bb4__26_i533_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__26_i533_0_stall_in_0_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__26_i533_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4__26_i533_0_NO_SHIFT_REG = rnode_346to347_bb4__26_i533_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4__26_i533_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4__26_i533_1_NO_SHIFT_REG = rnode_346to347_bb4__26_i533_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4__26_i533_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4__26_i533_2_NO_SHIFT_REG = rnode_346to347_bb4__26_i533_0_reg_347_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_379_380_0_inputs_ready;
 reg SFC_3_VALID_379_380_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_379_380_0_stall_in;
wire SFC_3_VALID_379_380_0_output_regs_ready;
 reg SFC_3_VALID_379_380_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_379_380_0_causedstall;

assign SFC_3_VALID_379_380_0_inputs_ready = 1'b1;
assign SFC_3_VALID_379_380_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_378_379_0_stall_in = 1'b0;
assign SFC_3_VALID_379_380_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_379_380_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_379_380_0_output_regs_ready)
		begin
			SFC_3_VALID_379_380_0_NO_SHIFT_REG <= SFC_3_VALID_378_379_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u50_valid_out;
wire local_bb4_var__u50_stall_in;
wire local_bb4_var__u50_inputs_ready;
wire local_bb4_var__u50_stall_local;
wire [31:0] local_bb4_var__u50;

assign local_bb4_var__u50_inputs_ready = (rnode_344to345_bb4_xor_i316_0_valid_out_NO_SHIFT_REG & rnode_344to345_bb4__29_i345_0_valid_out_NO_SHIFT_REG & rnode_343to345_bb4_or581_i374_0_valid_out_1_NO_SHIFT_REG & rnode_343to345_bb4_or581_i374_0_valid_out_0_NO_SHIFT_REG & rnode_344to345_bb4_reduction_0_i375_0_valid_out_NO_SHIFT_REG & rnode_343to345_bb4_cmp68_i377_0_valid_out_NO_SHIFT_REG & rnode_343to345_bb4_cmp71_not_i394_0_valid_out_NO_SHIFT_REG & rnode_343to345_bb4_shl_i381_0_valid_out_NO_SHIFT_REG & rnode_343to345_bb4_and75_i378_0_valid_out_NO_SHIFT_REG & rnode_344to345_bb4__40_i387_0_valid_out_NO_SHIFT_REG);
assign local_bb4_var__u50 = (rnode_344to345_bb4__29_i345_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb4_or112_i403);
assign local_bb4_var__u50_valid_out = 1'b1;
assign rnode_344to345_bb4_xor_i316_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__29_i345_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_or581_i374_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_or581_i374_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_reduction_0_i375_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp68_i377_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp71_not_i394_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_shl_i381_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_and75_i378_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__40_i387_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr217_i_stall_local;
wire [31:0] local_bb4_shr217_i;

assign local_bb4_shr217_i = ((rnode_344to345_bb4_and194_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i573_stall_local;
wire [31:0] local_bb4__pre_i573;

assign local_bb4__pre_i573 = ((rnode_344to345_bb4_and196_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i560_stall_local;
wire [31:0] local_bb4_or_i_i560;

assign local_bb4_or_i_i560 = ((local_bb4_shr_i_i559 & 32'h3FFFFFF) | (local_bb4_and202_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond293_i_stall_local;
wire [31:0] local_bb4_cond293_i;

assign local_bb4_cond293_i = (rnode_346to347_bb4__26_i533_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u51_stall_local;
wire [31:0] local_bb4_var__u51;

assign local_bb4_var__u51[31:1] = 31'h0;
assign local_bb4_var__u51[0] = rnode_346to347_bb4__26_i533_2_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_380_381_0_inputs_ready;
 reg SFC_3_VALID_380_381_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_380_381_0_stall_in;
wire SFC_3_VALID_380_381_0_output_regs_ready;
 reg SFC_3_VALID_380_381_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_380_381_0_causedstall;

assign SFC_3_VALID_380_381_0_inputs_ready = 1'b1;
assign SFC_3_VALID_380_381_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_379_380_0_stall_in = 1'b0;
assign SFC_3_VALID_380_381_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_380_381_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_380_381_0_output_regs_ready)
		begin
			SFC_3_VALID_380_381_0_NO_SHIFT_REG <= SFC_3_VALID_379_380_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_345to346_bb4_var__u50_0_valid_out_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u50_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_var__u50_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u50_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_var__u50_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u50_0_valid_out_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u50_0_stall_in_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_var__u50_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_345to346_bb4_var__u50_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to346_bb4_var__u50_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to346_bb4_var__u50_0_stall_in_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_345to346_bb4_var__u50_0_valid_out_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_345to346_bb4_var__u50_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in(local_bb4_var__u50),
	.data_out(rnode_345to346_bb4_var__u50_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_345to346_bb4_var__u50_0_reg_346_fifo.DEPTH = 1;
defparam rnode_345to346_bb4_var__u50_0_reg_346_fifo.DATA_WIDTH = 32;
defparam rnode_345to346_bb4_var__u50_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to346_bb4_var__u50_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_345to346_bb4_var__u50_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u50_stall_in = 1'b0;
assign rnode_345to346_bb4_var__u50_0_NO_SHIFT_REG = rnode_345to346_bb4_var__u50_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4_var__u50_0_stall_in_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_var__u50_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or220_i_stall_local;
wire [31:0] local_bb4_or220_i;

assign local_bb4_or220_i = ((local_bb4_shr217_i & 32'h7FFFFFF) | (rnode_344to345_bb4_and199_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool214_i_stall_local;
wire local_bb4_tobool214_i;

assign local_bb4_tobool214_i = ((local_bb4__pre_i573 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i561_stall_local;
wire [31:0] local_bb4_shr1_i_i561;

assign local_bb4_shr1_i_i561 = ((local_bb4_or_i_i560 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i590_stall_local;
wire [31:0] local_bb4_lnot_ext_i590;

assign local_bb4_lnot_ext_i590 = ((local_bb4_var__u51 & 32'h1) ^ 32'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_381_382_0_inputs_ready;
 reg SFC_3_VALID_381_382_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_381_382_0_stall_in;
wire SFC_3_VALID_381_382_0_output_regs_ready;
 reg SFC_3_VALID_381_382_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_381_382_0_causedstall;

assign SFC_3_VALID_381_382_0_inputs_ready = 1'b1;
assign SFC_3_VALID_381_382_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_380_381_0_stall_in = 1'b0;
assign SFC_3_VALID_381_382_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_381_382_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_381_382_0_output_regs_ready)
		begin
			SFC_3_VALID_381_382_0_NO_SHIFT_REG <= SFC_3_VALID_380_381_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 36
//  * capacity = 36
 logic rnode_346to382_bb4_var__u50_0_valid_out_NO_SHIFT_REG;
 logic rnode_346to382_bb4_var__u50_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_346to382_bb4_var__u50_0_NO_SHIFT_REG;
 logic rnode_346to382_bb4_var__u50_0_reg_382_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_346to382_bb4_var__u50_0_reg_382_NO_SHIFT_REG;
 logic rnode_346to382_bb4_var__u50_0_valid_out_reg_382_NO_SHIFT_REG;
 logic rnode_346to382_bb4_var__u50_0_stall_in_reg_382_NO_SHIFT_REG;
 logic rnode_346to382_bb4_var__u50_0_stall_out_reg_382_NO_SHIFT_REG;

acl_data_fifo rnode_346to382_bb4_var__u50_0_reg_382_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to382_bb4_var__u50_0_reg_382_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to382_bb4_var__u50_0_stall_in_reg_382_NO_SHIFT_REG),
	.valid_out(rnode_346to382_bb4_var__u50_0_valid_out_reg_382_NO_SHIFT_REG),
	.stall_out(rnode_346to382_bb4_var__u50_0_stall_out_reg_382_NO_SHIFT_REG),
	.data_in(rnode_345to346_bb4_var__u50_0_NO_SHIFT_REG),
	.data_out(rnode_346to382_bb4_var__u50_0_reg_382_NO_SHIFT_REG)
);

defparam rnode_346to382_bb4_var__u50_0_reg_382_fifo.DEPTH = 36;
defparam rnode_346to382_bb4_var__u50_0_reg_382_fifo.DATA_WIDTH = 32;
defparam rnode_346to382_bb4_var__u50_0_reg_382_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to382_bb4_var__u50_0_reg_382_fifo.IMPL = "shift_reg";

assign rnode_346to382_bb4_var__u50_0_reg_382_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_345to346_bb4_var__u50_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_346to382_bb4_var__u50_0_NO_SHIFT_REG = rnode_346to382_bb4_var__u50_0_reg_382_NO_SHIFT_REG;
assign rnode_346to382_bb4_var__u50_0_stall_in_reg_382_NO_SHIFT_REG = 1'b0;
assign rnode_346to382_bb4_var__u50_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i574_stall_local;
wire local_bb4__40_demorgan_i574;

assign local_bb4__40_demorgan_i574 = (rnode_343to345_bb4_cmp38_i_0_NO_SHIFT_REG | local_bb4_tobool214_i);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i575_stall_local;
wire local_bb4__42_i575;

assign local_bb4__42_i575 = (local_bb4_tobool214_i & local_bb4_not_cmp38_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i562_stall_local;
wire [31:0] local_bb4_or2_i_i562;

assign local_bb4_or2_i_i562 = ((local_bb4_shr1_i_i561 & 32'h1FFFFFF) | (local_bb4_or_i_i560 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_382_383_0_inputs_ready;
 reg SFC_3_VALID_382_383_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_382_383_0_stall_in;
wire SFC_3_VALID_382_383_0_output_regs_ready;
 reg SFC_3_VALID_382_383_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_382_383_0_causedstall;

assign SFC_3_VALID_382_383_0_inputs_ready = 1'b1;
assign SFC_3_VALID_382_383_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_381_382_0_stall_in = 1'b0;
assign SFC_3_VALID_382_383_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_382_383_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_382_383_0_output_regs_ready)
		begin
			SFC_3_VALID_382_383_0_NO_SHIFT_REG <= SFC_3_VALID_381_382_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_382to383_bb4_var__u50_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb4_var__u50_0_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb4_var__u50_1_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb4_var__u50_2_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_reg_383_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_382to383_bb4_var__u50_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_valid_out_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_stall_in_0_reg_383_NO_SHIFT_REG;
 logic rnode_382to383_bb4_var__u50_0_stall_out_reg_383_NO_SHIFT_REG;

acl_data_fifo rnode_382to383_bb4_var__u50_0_reg_383_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_382to383_bb4_var__u50_0_reg_383_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_382to383_bb4_var__u50_0_stall_in_0_reg_383_NO_SHIFT_REG),
	.valid_out(rnode_382to383_bb4_var__u50_0_valid_out_0_reg_383_NO_SHIFT_REG),
	.stall_out(rnode_382to383_bb4_var__u50_0_stall_out_reg_383_NO_SHIFT_REG),
	.data_in(rnode_346to382_bb4_var__u50_0_NO_SHIFT_REG),
	.data_out(rnode_382to383_bb4_var__u50_0_reg_383_NO_SHIFT_REG)
);

defparam rnode_382to383_bb4_var__u50_0_reg_383_fifo.DEPTH = 1;
defparam rnode_382to383_bb4_var__u50_0_reg_383_fifo.DATA_WIDTH = 32;
defparam rnode_382to383_bb4_var__u50_0_reg_383_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_382to383_bb4_var__u50_0_reg_383_fifo.IMPL = "shift_reg";

assign rnode_382to383_bb4_var__u50_0_reg_383_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_346to382_bb4_var__u50_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb4_var__u50_0_stall_in_0_reg_383_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb4_var__u50_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb4_var__u50_0_NO_SHIFT_REG = rnode_382to383_bb4_var__u50_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb4_var__u50_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb4_var__u50_1_NO_SHIFT_REG = rnode_382to383_bb4_var__u50_0_reg_383_NO_SHIFT_REG;
assign rnode_382to383_bb4_var__u50_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_382to383_bb4_var__u50_2_NO_SHIFT_REG = rnode_382to383_bb4_var__u50_0_reg_383_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__43_i576_stall_local;
wire [31:0] local_bb4__43_i576;

assign local_bb4__43_i576 = (local_bb4__42_i575 ? 32'h0 : (local_bb4__pre_i573 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i563_stall_local;
wire [31:0] local_bb4_shr3_i_i563;

assign local_bb4_shr3_i_i563 = ((local_bb4_or2_i_i562 & 32'h7FFFFFF) >> 32'h4);

// This section implements a registered operation.
// 
wire SFC_3_VALID_383_384_0_inputs_ready;
 reg SFC_3_VALID_383_384_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_383_384_0_stall_in;
wire SFC_3_VALID_383_384_0_output_regs_ready;
 reg SFC_3_VALID_383_384_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_383_384_0_causedstall;

assign SFC_3_VALID_383_384_0_inputs_ready = 1'b1;
assign SFC_3_VALID_383_384_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_382_383_0_stall_in = 1'b0;
assign SFC_3_VALID_383_384_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_383_384_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_383_384_0_output_regs_ready)
		begin
			SFC_3_VALID_383_384_0_NO_SHIFT_REG <= SFC_3_VALID_382_383_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr_i220_stall_local;
wire [31:0] local_bb4_shr_i220;

assign local_bb4_shr_i220 = (rnode_382to383_bb4_var__u50_0_NO_SHIFT_REG >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and5_i226_stall_local;
wire [31:0] local_bb4_and5_i226;

assign local_bb4_and5_i226 = (rnode_382to383_bb4_var__u50_2_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i564_stall_local;
wire [31:0] local_bb4_or4_i_i564;

assign local_bb4_or4_i_i564 = ((local_bb4_shr3_i_i563 & 32'h7FFFFF) | (local_bb4_or2_i_i562 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_384_385_0_inputs_ready;
 reg SFC_3_VALID_384_385_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_384_385_0_stall_in;
wire SFC_3_VALID_384_385_0_output_regs_ready;
 reg SFC_3_VALID_384_385_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_384_385_0_causedstall;

assign SFC_3_VALID_384_385_0_inputs_ready = 1'b1;
assign SFC_3_VALID_384_385_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_383_384_0_stall_in = 1'b0;
assign SFC_3_VALID_384_385_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_384_385_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_384_385_0_output_regs_ready)
		begin
			SFC_3_VALID_384_385_0_NO_SHIFT_REG <= SFC_3_VALID_383_384_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and_i221_stall_local;
wire [31:0] local_bb4_and_i221;

assign local_bb4_and_i221 = ((local_bb4_shr_i220 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i232_stall_local;
wire local_bb4_lnot14_i232;

assign local_bb4_lnot14_i232 = ((local_bb4_and5_i226 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i254_stall_local;
wire [31:0] local_bb4_or_i254;

assign local_bb4_or_i254 = ((local_bb4_and5_i226 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i565_stall_local;
wire [31:0] local_bb4_shr5_i_i565;

assign local_bb4_shr5_i_i565 = ((local_bb4_or4_i_i564 & 32'h7FFFFFF) >> 32'h8);

// This section implements a registered operation.
// 
wire SFC_3_VALID_385_386_0_inputs_ready;
 reg SFC_3_VALID_385_386_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_385_386_0_stall_in;
wire SFC_3_VALID_385_386_0_output_regs_ready;
 reg SFC_3_VALID_385_386_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_385_386_0_causedstall;

assign SFC_3_VALID_385_386_0_inputs_ready = 1'b1;
assign SFC_3_VALID_385_386_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_384_385_0_stall_in = 1'b0;
assign SFC_3_VALID_385_386_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_385_386_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_385_386_0_output_regs_ready)
		begin
			SFC_3_VALID_385_386_0_NO_SHIFT_REG <= SFC_3_VALID_384_385_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i228_stall_local;
wire local_bb4_lnot_i228;

assign local_bb4_lnot_i228 = ((local_bb4_and_i221 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i230_stall_local;
wire local_bb4_cmp_i230;

assign local_bb4_cmp_i230 = ((local_bb4_and_i221 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i232_valid_out;
wire local_bb4_lnot14_i232_stall_in;
wire local_bb4_conv_i_i256_valid_out;
wire local_bb4_conv_i_i256_stall_in;
wire local_bb4_conv_i_i256_inputs_ready;
wire local_bb4_conv_i_i256_stall_local;
wire [63:0] local_bb4_conv_i_i256;

assign local_bb4_conv_i_i256_inputs_ready = rnode_382to383_bb4_var__u50_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_conv_i_i256[63:32] = 32'h0;
assign local_bb4_conv_i_i256[31:0] = ((local_bb4_or_i254 & 32'hFFFFFF) | 32'h800000);
assign local_bb4_lnot14_i232_valid_out = 1'b1;
assign local_bb4_conv_i_i256_valid_out = 1'b1;
assign rnode_382to383_bb4_var__u50_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i566_stall_local;
wire [31:0] local_bb4_or6_i_i566;

assign local_bb4_or6_i_i566 = ((local_bb4_shr5_i_i565 & 32'h7FFFF) | (local_bb4_or4_i_i564 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_386_387_0_inputs_ready;
 reg SFC_3_VALID_386_387_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_386_387_0_stall_in;
wire SFC_3_VALID_386_387_0_output_regs_ready;
 reg SFC_3_VALID_386_387_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_386_387_0_causedstall;

assign SFC_3_VALID_386_387_0_inputs_ready = 1'b1;
assign SFC_3_VALID_386_387_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_385_386_0_stall_in = 1'b0;
assign SFC_3_VALID_386_387_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_386_387_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_386_387_0_output_regs_ready)
		begin
			SFC_3_VALID_386_387_0_NO_SHIFT_REG <= SFC_3_VALID_385_386_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_lnot14_i232_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot14_i232_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_lnot14_i232_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_lnot14_i232_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_lnot14_i232_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_lnot14_i232_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_lnot14_i232_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_lnot14_i232),
	.data_out(rnode_383to384_bb4_lnot14_i232_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_lnot14_i232_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_lnot14_i232_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_lnot14_i232_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_lnot14_i232_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_lnot14_i232_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot14_i232_stall_in = 1'b0;
assign rnode_383to384_bb4_lnot14_i232_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot14_i232_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_lnot14_i232_0_NO_SHIFT_REG = rnode_383to384_bb4_lnot14_i232_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_lnot14_i232_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_lnot14_i232_1_NO_SHIFT_REG = rnode_383to384_bb4_lnot14_i232_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_lnot14_i232_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_lnot14_i232_2_NO_SHIFT_REG = rnode_383to384_bb4_lnot14_i232_0_reg_384_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i567_stall_local;
wire [31:0] local_bb4_shr7_i_i567;

assign local_bb4_shr7_i_i567 = ((local_bb4_or6_i_i566 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i568_stall_local;
wire [31:0] local_bb4_or6_masked_i_i568;

assign local_bb4_or6_masked_i_i568 = ((local_bb4_or6_i_i566 & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_387_388_0_inputs_ready;
 reg SFC_3_VALID_387_388_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_387_388_0_stall_in_0;
 reg SFC_3_VALID_387_388_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_387_388_0_stall_in_1;
wire SFC_3_VALID_387_388_0_output_regs_ready;
 reg SFC_3_VALID_387_388_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_387_388_0_causedstall;

assign SFC_3_VALID_387_388_0_inputs_ready = 1'b1;
assign SFC_3_VALID_387_388_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_386_387_0_stall_in = 1'b0;
assign SFC_3_VALID_387_388_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_387_388_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_387_388_0_output_regs_ready)
		begin
			SFC_3_VALID_387_388_0_NO_SHIFT_REG <= SFC_3_VALID_386_387_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_not_i251_stall_local;
wire local_bb4_lnot14_not_i251;

assign local_bb4_lnot14_not_i251 = (rnode_383to384_bb4_lnot14_i232_2_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i569_stall_local;
wire [31:0] local_bb4_neg_i_i569;

assign local_bb4_neg_i_i569 = ((local_bb4_or6_masked_i_i568 & 32'h7FFFFFF) | (local_bb4_shr7_i_i567 & 32'h7FF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_388_389_0_inputs_ready;
 reg SFC_3_VALID_388_389_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_388_389_0_stall_in;
wire SFC_3_VALID_388_389_0_output_regs_ready;
 reg SFC_3_VALID_388_389_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_388_389_0_causedstall;

assign SFC_3_VALID_388_389_0_inputs_ready = 1'b1;
assign SFC_3_VALID_388_389_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_387_388_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_388_389_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_388_389_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_388_389_0_output_regs_ready)
		begin
			SFC_3_VALID_388_389_0_NO_SHIFT_REG <= SFC_3_VALID_387_388_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_sum_312_pop9_c1_ene6_valid_out;
wire local_bb4_sum_312_pop9_c1_ene6_stall_in;
wire local_bb4_sum_312_pop9_c1_ene6_inputs_ready;
wire local_bb4_sum_312_pop9_c1_ene6_stall_local;
wire [31:0] local_bb4_sum_312_pop9_c1_ene6;
wire local_bb4_sum_312_pop9_c1_ene6_fu_valid_out;
wire local_bb4_sum_312_pop9_c1_ene6_fu_stall_out;

acl_pop local_bb4_sum_312_pop9_c1_ene6_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_387to388_bb4_c1_ene5_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_387to388_bb4_c1_ene6_0_NO_SHIFT_REG),
	.stall_out(local_bb4_sum_312_pop9_c1_ene6_fu_stall_out),
	.valid_in(SFC_3_VALID_387_388_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sum_312_pop9_c1_ene6_fu_valid_out),
	.stall_in(local_bb4_sum_312_pop9_c1_ene6_stall_local),
	.data_out(local_bb4_sum_312_pop9_c1_ene6),
	.feedback_in(feedback_data_in_9),
	.feedback_valid_in(feedback_valid_in_9),
	.feedback_stall_out(feedback_stall_out_9)
);

defparam local_bb4_sum_312_pop9_c1_ene6_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_sum_312_pop9_c1_ene6_feedback.DATA_WIDTH = 32;
defparam local_bb4_sum_312_pop9_c1_ene6_feedback.STYLE = "REGULAR";

assign local_bb4_sum_312_pop9_c1_ene6_inputs_ready = (SFC_3_VALID_387_388_0_valid_out_1_NO_SHIFT_REG & rnode_387to388_bb4_c1_ene5_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG);
assign local_bb4_sum_312_pop9_c1_ene6_stall_local = 1'b0;
assign local_bb4_sum_312_pop9_c1_ene6_valid_out = 1'b1;
assign SFC_3_VALID_387_388_0_stall_in_1 = 1'b0;
assign rnode_387to388_bb4_c1_ene5_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i570_stall_local;
wire [31:0] local_bb4_and_i_i570;

assign local_bb4_and_i_i570 = ((local_bb4_neg_i_i569 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_389_390_0_inputs_ready;
 reg SFC_3_VALID_389_390_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_389_390_0_stall_in;
wire SFC_3_VALID_389_390_0_output_regs_ready;
 reg SFC_3_VALID_389_390_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_389_390_0_causedstall;

assign SFC_3_VALID_389_390_0_inputs_ready = 1'b1;
assign SFC_3_VALID_389_390_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_388_389_0_stall_in = 1'b0;
assign SFC_3_VALID_389_390_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_389_390_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_389_390_0_output_regs_ready)
		begin
			SFC_3_VALID_389_390_0_NO_SHIFT_REG <= SFC_3_VALID_388_389_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_sum_312_pop9_c1_ene6_1_NO_SHIFT_REG;
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_valid_out_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_in_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_in_0_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_valid_out_0_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb4_sum_312_pop9_c1_ene6),
	.data_out(rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_sum_312_pop9_c1_ene6_stall_in = 1'b0;
assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_in_0_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG = rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_1_NO_SHIFT_REG = rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_reg_389_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i570_valid_out;
wire local_bb4__and_i_i570_stall_in;
wire local_bb4__and_i_i570_inputs_ready;
wire local_bb4__and_i_i570_stall_local;
wire [31:0] local_bb4__and_i_i570;

thirtysix_six_comp local_bb4__and_i_i570_popcnt_instance (
	.data((local_bb4_and_i_i570 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i570)
);


assign local_bb4__and_i_i570_inputs_ready = rnode_343to344_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i570_valid_out = 1'b1;
assign rnode_343to344_bb4_add193_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_390_391_0_inputs_ready;
 reg SFC_3_VALID_390_391_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_390_391_0_stall_in;
wire SFC_3_VALID_390_391_0_output_regs_ready;
 reg SFC_3_VALID_390_391_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_390_391_0_causedstall;

assign SFC_3_VALID_390_391_0_inputs_ready = 1'b1;
assign SFC_3_VALID_390_391_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_389_390_0_stall_in = 1'b0;
assign SFC_3_VALID_390_391_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_390_391_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_390_391_0_output_regs_ready)
		begin
			SFC_3_VALID_390_391_0_NO_SHIFT_REG <= SFC_3_VALID_389_390_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u52_stall_local;
wire [31:0] local_bb4_var__u52;

assign local_bb4_var__u52 = rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_valid_out_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_valid_out_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(rnode_388to389_bb4_sum_312_pop9_c1_ene6_1_NO_SHIFT_REG),
	.data_out(rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_fifo.DATA_WIDTH = 32;
defparam rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG = rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_344to345_bb4__and_i_i570_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4__and_i_i570_0_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4__and_i_i570_1_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4__and_i_i570_2_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_reg_345_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_344to345_bb4__and_i_i570_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_valid_out_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_stall_in_0_reg_345_NO_SHIFT_REG;
 logic rnode_344to345_bb4__and_i_i570_0_stall_out_reg_345_NO_SHIFT_REG;

acl_data_fifo rnode_344to345_bb4__and_i_i570_0_reg_345_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_344to345_bb4__and_i_i570_0_reg_345_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_344to345_bb4__and_i_i570_0_stall_in_0_reg_345_NO_SHIFT_REG),
	.valid_out(rnode_344to345_bb4__and_i_i570_0_valid_out_0_reg_345_NO_SHIFT_REG),
	.stall_out(rnode_344to345_bb4__and_i_i570_0_stall_out_reg_345_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i570 & 32'h3F)),
	.data_out(rnode_344to345_bb4__and_i_i570_0_reg_345_NO_SHIFT_REG)
);

defparam rnode_344to345_bb4__and_i_i570_0_reg_345_fifo.DEPTH = 1;
defparam rnode_344to345_bb4__and_i_i570_0_reg_345_fifo.DATA_WIDTH = 32;
defparam rnode_344to345_bb4__and_i_i570_0_reg_345_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_344to345_bb4__and_i_i570_0_reg_345_fifo.IMPL = "shift_reg";

assign rnode_344to345_bb4__and_i_i570_0_reg_345_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i570_stall_in = 1'b0;
assign rnode_344to345_bb4__and_i_i570_0_stall_in_0_reg_345_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__and_i_i570_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_344to345_bb4__and_i_i570_0_NO_SHIFT_REG = rnode_344to345_bb4__and_i_i570_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4__and_i_i570_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_344to345_bb4__and_i_i570_1_NO_SHIFT_REG = rnode_344to345_bb4__and_i_i570_0_reg_345_NO_SHIFT_REG;
assign rnode_344to345_bb4__and_i_i570_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_344to345_bb4__and_i_i570_2_NO_SHIFT_REG = rnode_344to345_bb4__and_i_i570_0_reg_345_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_391_392_0_inputs_ready;
 reg SFC_3_VALID_391_392_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_391_392_0_stall_in;
wire SFC_3_VALID_391_392_0_output_regs_ready;
 reg SFC_3_VALID_391_392_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_391_392_0_causedstall;

assign SFC_3_VALID_391_392_0_inputs_ready = 1'b1;
assign SFC_3_VALID_391_392_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_390_391_0_stall_in = 1'b0;
assign SFC_3_VALID_391_392_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_391_392_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_391_392_0_output_regs_ready)
		begin
			SFC_3_VALID_391_392_0_NO_SHIFT_REG <= SFC_3_VALID_390_391_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and2_i2_stall_local;
wire [31:0] local_bb4_and2_i2;

assign local_bb4_and2_i2 = (local_bb4_var__u52 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i_stall_local;
wire [31:0] local_bb4_and12_i;

assign local_bb4_and12_i = (local_bb4_var__u52 & 32'hFFFF);

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_NO_SHIFT_REG;
 logic rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_fifo.DEPTH = 5;
defparam rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4_sum_312_pop9_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG = rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_reg_395_NO_SHIFT_REG;
assign rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i571_stall_local;
wire [31:0] local_bb4_and9_i_i571;

assign local_bb4_and9_i_i571 = ((rnode_344to345_bb4__and_i_i570_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and204_i_stall_local;
wire [31:0] local_bb4_and204_i;

assign local_bb4_and204_i = ((rnode_344to345_bb4__and_i_i570_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and207_i_stall_local;
wire [31:0] local_bb4_and207_i;

assign local_bb4_and207_i = ((rnode_344to345_bb4__and_i_i570_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements a registered operation.
// 
wire SFC_3_VALID_392_393_0_inputs_ready;
 reg SFC_3_VALID_392_393_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_392_393_0_stall_in_0;
 reg SFC_3_VALID_392_393_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_392_393_0_stall_in_1;
wire SFC_3_VALID_392_393_0_output_regs_ready;
 reg SFC_3_VALID_392_393_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_392_393_0_causedstall;

assign SFC_3_VALID_392_393_0_inputs_ready = 1'b1;
assign SFC_3_VALID_392_393_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_391_392_0_stall_in = 1'b0;
assign SFC_3_VALID_392_393_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_392_393_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_392_393_0_output_regs_ready)
		begin
			SFC_3_VALID_392_393_0_NO_SHIFT_REG <= SFC_3_VALID_391_392_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_stall_local;
wire [31:0] local_bb4_shr3_i;

assign local_bb4_shr3_i = ((local_bb4_and2_i2 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_fifo.DATA_WIDTH = 32;
defparam rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_390to395_bb4_sum_312_pop9_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG = rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_sub240_i_stall_local;
wire [31:0] local_bb4_sub240_i;

assign local_bb4_sub240_i = (32'h0 - (local_bb4_and9_i_i571 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl205_i_stall_local;
wire [31:0] local_bb4_shl205_i;

assign local_bb4_shl205_i = ((rnode_344to345_bb4_and194_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and204_i & 32'h18));

// This section implements a registered operation.
// 
wire SFC_3_VALID_393_394_0_inputs_ready;
 reg SFC_3_VALID_393_394_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_393_394_0_stall_in;
wire SFC_3_VALID_393_394_0_output_regs_ready;
 reg SFC_3_VALID_393_394_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_393_394_0_causedstall;

assign SFC_3_VALID_393_394_0_inputs_ready = 1'b1;
assign SFC_3_VALID_393_394_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_392_393_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_393_394_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_393_394_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_393_394_0_output_regs_ready)
		begin
			SFC_3_VALID_393_394_0_NO_SHIFT_REG <= SFC_3_VALID_392_393_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_t_313_pop8_c1_ene4_valid_out;
wire local_bb4_t_313_pop8_c1_ene4_stall_in;
wire local_bb4_t_313_pop8_c1_ene4_inputs_ready;
wire local_bb4_t_313_pop8_c1_ene4_stall_local;
wire [31:0] local_bb4_t_313_pop8_c1_ene4;
wire local_bb4_t_313_pop8_c1_ene4_fu_valid_out;
wire local_bb4_t_313_pop8_c1_ene4_fu_stall_out;

acl_pop local_bb4_t_313_pop8_c1_ene4_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_392to393_bb4_c1_ene5_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_392to393_bb4_c1_ene4_0_NO_SHIFT_REG),
	.stall_out(local_bb4_t_313_pop8_c1_ene4_fu_stall_out),
	.valid_in(SFC_3_VALID_392_393_0_NO_SHIFT_REG),
	.valid_out(local_bb4_t_313_pop8_c1_ene4_fu_valid_out),
	.stall_in(local_bb4_t_313_pop8_c1_ene4_stall_local),
	.data_out(local_bb4_t_313_pop8_c1_ene4),
	.feedback_in(feedback_data_in_8),
	.feedback_valid_in(feedback_valid_in_8),
	.feedback_stall_out(feedback_stall_out_8)
);

defparam local_bb4_t_313_pop8_c1_ene4_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_t_313_pop8_c1_ene4_feedback.DATA_WIDTH = 32;
defparam local_bb4_t_313_pop8_c1_ene4_feedback.STYLE = "REGULAR";

assign local_bb4_t_313_pop8_c1_ene4_inputs_ready = (SFC_3_VALID_392_393_0_valid_out_1_NO_SHIFT_REG & rnode_392to393_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG);
assign local_bb4_t_313_pop8_c1_ene4_stall_local = 1'b0;
assign local_bb4_t_313_pop8_c1_ene4_valid_out = 1'b1;
assign SFC_3_VALID_392_393_0_stall_in_1 = 1'b0;
assign rnode_392to393_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cond245_i_stall_local;
wire [31:0] local_bb4_cond245_i;

assign local_bb4_cond245_i = (rnode_343to345_bb4_cmp38_i_2_NO_SHIFT_REG ? local_bb4_sub240_i : (local_bb4__43_i576 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i572_stall_local;
wire [31:0] local_bb4_and206_i572;

assign local_bb4_and206_i572 = (local_bb4_shl205_i & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_394_395_0_inputs_ready;
 reg SFC_3_VALID_394_395_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_394_395_0_stall_in;
wire SFC_3_VALID_394_395_0_output_regs_ready;
 reg SFC_3_VALID_394_395_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_394_395_0_causedstall;

assign SFC_3_VALID_394_395_0_inputs_ready = 1'b1;
assign SFC_3_VALID_394_395_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_393_394_0_stall_in = 1'b0;
assign SFC_3_VALID_394_395_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_394_395_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_394_395_0_output_regs_ready)
		begin
			SFC_3_VALID_394_395_0_NO_SHIFT_REG <= SFC_3_VALID_393_394_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_t_313_pop8_c1_ene4_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_valid_out_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_in_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_in_0_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb4_t_313_pop8_c1_ene4_0_valid_out_0_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in(local_bb4_t_313_pop8_c1_ene4),
	.data_out(rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_t_313_pop8_c1_ene4_stall_in = 1'b0;
assign rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_in_0_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_t_313_pop8_c1_ene4_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG = rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_t_313_pop8_c1_ene4_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_t_313_pop8_c1_ene4_1_NO_SHIFT_REG = rnode_393to394_bb4_t_313_pop8_c1_ene4_0_reg_394_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add246_i_stall_local;
wire [31:0] local_bb4_add246_i;

assign local_bb4_add246_i = (local_bb4_cond245_i + (rnode_343to345_bb4_and17_i511_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i581_stall_local;
wire [31:0] local_bb4_fold_i581;

assign local_bb4_fold_i581 = (local_bb4_cond245_i + (rnode_343to345_bb4_shr16_i510_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl208_i_stall_local;
wire [31:0] local_bb4_shl208_i;

assign local_bb4_shl208_i = ((local_bb4_and206_i572 & 32'h7FFFFFF) << (local_bb4_and207_i & 32'h7));

// This section implements a registered operation.
// 
wire SFC_3_VALID_395_396_0_inputs_ready;
 reg SFC_3_VALID_395_396_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_395_396_0_stall_in;
wire SFC_3_VALID_395_396_0_output_regs_ready;
 reg SFC_3_VALID_395_396_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_395_396_0_causedstall;

assign SFC_3_VALID_395_396_0_inputs_ready = 1'b1;
assign SFC_3_VALID_395_396_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_394_395_0_stall_in = 1'b0;
assign SFC_3_VALID_395_396_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_395_396_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_395_396_0_output_regs_ready)
		begin
			SFC_3_VALID_395_396_0_NO_SHIFT_REG <= SFC_3_VALID_394_395_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u53_stall_local;
wire [31:0] local_bb4_var__u53;

assign local_bb4_var__u53 = rnode_393to394_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_t_313_pop8_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_394to395_bb4_t_313_pop8_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_t_313_pop8_c1_ene4_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_t_313_pop8_c1_ene4_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(rnode_393to394_bb4_t_313_pop8_c1_ene4_1_NO_SHIFT_REG),
	.data_out(rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG = rnode_394to395_bb4_t_313_pop8_c1_ene4_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_t_313_pop8_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and251_i_stall_local;
wire [31:0] local_bb4_and251_i;

assign local_bb4_and251_i = (local_bb4_fold_i581 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i586_stall_local;
wire [31:0] local_bb4_and270_i586;

assign local_bb4_and270_i586 = (local_bb4_fold_i581 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and209_i_stall_local;
wire [31:0] local_bb4_and209_i;

assign local_bb4_and209_i = (local_bb4_shl208_i & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_396_397_0_inputs_ready;
 reg SFC_3_VALID_396_397_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_396_397_0_stall_in_0;
 reg SFC_3_VALID_396_397_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_396_397_0_stall_in_1;
wire SFC_3_VALID_396_397_0_output_regs_ready;
 reg SFC_3_VALID_396_397_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_396_397_0_causedstall;

assign SFC_3_VALID_396_397_0_inputs_ready = 1'b1;
assign SFC_3_VALID_396_397_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_395_396_0_stall_in = 1'b0;
assign SFC_3_VALID_396_397_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_396_397_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_396_397_0_output_regs_ready)
		begin
			SFC_3_VALID_396_397_0_NO_SHIFT_REG <= SFC_3_VALID_395_396_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and2_i13_stall_local;
wire [31:0] local_bb4_and2_i13;

assign local_bb4_and2_i13 = (local_bb4_var__u53 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i18_stall_local;
wire [31:0] local_bb4_and12_i18;

assign local_bb4_and12_i18 = (local_bb4_var__u53 & 32'hFFFF);

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_395to400_bb4_t_313_pop8_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_395to400_bb4_t_313_pop8_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_395to400_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_NO_SHIFT_REG;
 logic rnode_395to400_bb4_t_313_pop8_c1_ene4_0_valid_out_reg_400_NO_SHIFT_REG;
 logic rnode_395to400_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_400_NO_SHIFT_REG;
 logic rnode_395to400_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to400_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_395to400_bb4_t_313_pop8_c1_ene4_0_valid_out_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_395to400_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in(rnode_394to395_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_fifo.DEPTH = 5;
defparam rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_fifo.DATA_WIDTH = 32;
defparam rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4_t_313_pop8_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to400_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG = rnode_395to400_bb4_t_313_pop8_c1_ene4_0_reg_400_NO_SHIFT_REG;
assign rnode_395to400_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_395to400_bb4_t_313_pop8_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__44_i577_stall_local;
wire [31:0] local_bb4__44_i577;

assign local_bb4__44_i577 = (local_bb4__40_demorgan_i574 ? (local_bb4_and209_i & 32'h7FFFFFF) : (local_bb4_or220_i & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_397_398_0_inputs_ready;
 reg SFC_3_VALID_397_398_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_397_398_0_stall_in;
wire SFC_3_VALID_397_398_0_output_regs_ready;
 reg SFC_3_VALID_397_398_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_397_398_0_causedstall;

assign SFC_3_VALID_397_398_0_inputs_ready = 1'b1;
assign SFC_3_VALID_397_398_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_396_397_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_397_398_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_397_398_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_397_398_0_output_regs_ready)
		begin
			SFC_3_VALID_397_398_0_NO_SHIFT_REG <= SFC_3_VALID_396_397_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i14_stall_local;
wire [31:0] local_bb4_shr3_i14;

assign local_bb4_shr3_i14 = ((local_bb4_and2_i13 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4_t_313_pop8_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_400to401_bb4_t_313_pop8_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_400to401_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_t_313_pop8_c1_ene4_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4_t_313_pop8_c1_ene4_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4_t_313_pop8_c1_ene4_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(rnode_395to400_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_fifo.DATA_WIDTH = 32;
defparam rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_395to400_bb4_t_313_pop8_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG = rnode_400to401_bb4_t_313_pop8_c1_ene4_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_t_313_pop8_c1_ene4_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_t_313_pop8_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and251_i_valid_out;
wire local_bb4_and251_i_stall_in;
wire local_bb4_and270_i586_valid_out;
wire local_bb4_and270_i586_stall_in;
wire local_bb4_add246_i_valid_out;
wire local_bb4_add246_i_stall_in;
wire local_bb4__45_i578_valid_out;
wire local_bb4__45_i578_stall_in;
wire local_bb4_not_cmp38_i_valid_out_1;
wire local_bb4_not_cmp38_i_stall_in_1;
wire local_bb4__45_i578_inputs_ready;
wire local_bb4__45_i578_stall_local;
wire [31:0] local_bb4__45_i578;

assign local_bb4__45_i578_inputs_ready = (rnode_343to345_bb4_shr16_i510_0_valid_out_NO_SHIFT_REG & rnode_343to345_bb4_and17_i511_0_valid_out_NO_SHIFT_REG & rnode_343to345_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG & rnode_343to345_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG & rnode_344to345_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG & rnode_343to345_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG & rnode_344to345_bb4_and196_i_0_valid_out_NO_SHIFT_REG & rnode_344to345_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG & rnode_344to345_bb4_and199_i_0_valid_out_NO_SHIFT_REG & rnode_344to345_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG & rnode_344to345_bb4__and_i_i570_0_valid_out_1_NO_SHIFT_REG & rnode_344to345_bb4__and_i_i570_0_valid_out_2_NO_SHIFT_REG & rnode_344to345_bb4__and_i_i570_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i578 = (local_bb4__42_i575 ? (rnode_344to345_bb4_and194_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i577 & 32'h7FFFFFF));
assign local_bb4_and251_i_valid_out = 1'b1;
assign local_bb4_and270_i586_valid_out = 1'b1;
assign local_bb4_add246_i_valid_out = 1'b1;
assign local_bb4__45_i578_valid_out = 1'b1;
assign local_bb4_not_cmp38_i_valid_out_1 = 1'b1;
assign rnode_343to345_bb4_shr16_i510_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_and17_i511_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp38_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and194_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_343to345_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and196_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and194_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and199_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4_and194_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__and_i_i570_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__and_i_i570_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_344to345_bb4__and_i_i570_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_398_399_0_inputs_ready;
 reg SFC_3_VALID_398_399_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_398_399_0_stall_in;
wire SFC_3_VALID_398_399_0_output_regs_ready;
 reg SFC_3_VALID_398_399_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_398_399_0_causedstall;

assign SFC_3_VALID_398_399_0_inputs_ready = 1'b1;
assign SFC_3_VALID_398_399_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_397_398_0_stall_in = 1'b0;
assign SFC_3_VALID_398_399_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_398_399_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_398_399_0_output_regs_ready)
		begin
			SFC_3_VALID_398_399_0_NO_SHIFT_REG <= SFC_3_VALID_397_398_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_345to346_bb4_and251_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and251_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_and251_i_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and251_i_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_and251_i_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and251_i_0_valid_out_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and251_i_0_stall_in_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_and251_i_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_345to346_bb4_and251_i_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to346_bb4_and251_i_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to346_bb4_and251_i_0_stall_in_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_345to346_bb4_and251_i_0_valid_out_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_345to346_bb4_and251_i_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in((local_bb4_and251_i & 32'hFF)),
	.data_out(rnode_345to346_bb4_and251_i_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_345to346_bb4_and251_i_0_reg_346_fifo.DEPTH = 1;
defparam rnode_345to346_bb4_and251_i_0_reg_346_fifo.DATA_WIDTH = 32;
defparam rnode_345to346_bb4_and251_i_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to346_bb4_and251_i_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_345to346_bb4_and251_i_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and251_i_stall_in = 1'b0;
assign rnode_345to346_bb4_and251_i_0_NO_SHIFT_REG = rnode_345to346_bb4_and251_i_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4_and251_i_0_stall_in_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_and251_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_345to347_bb4_and270_i586_0_valid_out_NO_SHIFT_REG;
 logic rnode_345to347_bb4_and270_i586_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_345to347_bb4_and270_i586_0_NO_SHIFT_REG;
 logic rnode_345to347_bb4_and270_i586_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_345to347_bb4_and270_i586_0_reg_347_NO_SHIFT_REG;
 logic rnode_345to347_bb4_and270_i586_0_valid_out_reg_347_NO_SHIFT_REG;
 logic rnode_345to347_bb4_and270_i586_0_stall_in_reg_347_NO_SHIFT_REG;
 logic rnode_345to347_bb4_and270_i586_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_345to347_bb4_and270_i586_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to347_bb4_and270_i586_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to347_bb4_and270_i586_0_stall_in_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_345to347_bb4_and270_i586_0_valid_out_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_345to347_bb4_and270_i586_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in((local_bb4_and270_i586 & 32'hFF800000)),
	.data_out(rnode_345to347_bb4_and270_i586_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_345to347_bb4_and270_i586_0_reg_347_fifo.DEPTH = 2;
defparam rnode_345to347_bb4_and270_i586_0_reg_347_fifo.DATA_WIDTH = 32;
defparam rnode_345to347_bb4_and270_i586_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to347_bb4_and270_i586_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_345to347_bb4_and270_i586_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and270_i586_stall_in = 1'b0;
assign rnode_345to347_bb4_and270_i586_0_NO_SHIFT_REG = rnode_345to347_bb4_and270_i586_0_reg_347_NO_SHIFT_REG;
assign rnode_345to347_bb4_and270_i586_0_stall_in_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_345to347_bb4_and270_i586_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_345to346_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4_add246_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_add246_i_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_345to346_bb4_add246_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_add246_i_1_NO_SHIFT_REG;
 logic rnode_345to346_bb4_add246_i_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4_add246_i_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_add246_i_0_valid_out_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_add246_i_0_stall_in_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_add246_i_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_345to346_bb4_add246_i_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to346_bb4_add246_i_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to346_bb4_add246_i_0_stall_in_0_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_345to346_bb4_add246_i_0_valid_out_0_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_345to346_bb4_add246_i_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in(local_bb4_add246_i),
	.data_out(rnode_345to346_bb4_add246_i_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_345to346_bb4_add246_i_0_reg_346_fifo.DEPTH = 1;
defparam rnode_345to346_bb4_add246_i_0_reg_346_fifo.DATA_WIDTH = 32;
defparam rnode_345to346_bb4_add246_i_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to346_bb4_add246_i_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_345to346_bb4_add246_i_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add246_i_stall_in = 1'b0;
assign rnode_345to346_bb4_add246_i_0_stall_in_0_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_345to346_bb4_add246_i_0_NO_SHIFT_REG = rnode_345to346_bb4_add246_i_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_345to346_bb4_add246_i_1_NO_SHIFT_REG = rnode_345to346_bb4_add246_i_0_reg_346_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_345to346_bb4__45_i578_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4__45_i578_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4__45_i578_1_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4__45_i578_2_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_345to346_bb4__45_i578_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_valid_out_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_stall_in_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4__45_i578_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_345to346_bb4__45_i578_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to346_bb4__45_i578_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to346_bb4__45_i578_0_stall_in_0_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_345to346_bb4__45_i578_0_valid_out_0_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_345to346_bb4__45_i578_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in((local_bb4__45_i578 & 32'hFFFFFFF)),
	.data_out(rnode_345to346_bb4__45_i578_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_345to346_bb4__45_i578_0_reg_346_fifo.DEPTH = 1;
defparam rnode_345to346_bb4__45_i578_0_reg_346_fifo.DATA_WIDTH = 32;
defparam rnode_345to346_bb4__45_i578_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to346_bb4__45_i578_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_345to346_bb4__45_i578_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i578_stall_in = 1'b0;
assign rnode_345to346_bb4__45_i578_0_stall_in_0_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4__45_i578_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_345to346_bb4__45_i578_0_NO_SHIFT_REG = rnode_345to346_bb4__45_i578_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4__45_i578_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_345to346_bb4__45_i578_1_NO_SHIFT_REG = rnode_345to346_bb4__45_i578_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4__45_i578_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_345to346_bb4__45_i578_2_NO_SHIFT_REG = rnode_345to346_bb4__45_i578_0_reg_346_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_345to346_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_345to346_bb4_not_cmp38_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_345to346_bb4_not_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_345to346_bb4_not_cmp38_i_0_reg_346_inputs_ready_NO_SHIFT_REG;
 logic rnode_345to346_bb4_not_cmp38_i_0_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_not_cmp38_i_0_valid_out_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_not_cmp38_i_0_stall_in_reg_346_NO_SHIFT_REG;
 logic rnode_345to346_bb4_not_cmp38_i_0_stall_out_reg_346_NO_SHIFT_REG;

acl_data_fifo rnode_345to346_bb4_not_cmp38_i_0_reg_346_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_345to346_bb4_not_cmp38_i_0_reg_346_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_345to346_bb4_not_cmp38_i_0_stall_in_reg_346_NO_SHIFT_REG),
	.valid_out(rnode_345to346_bb4_not_cmp38_i_0_valid_out_reg_346_NO_SHIFT_REG),
	.stall_out(rnode_345to346_bb4_not_cmp38_i_0_stall_out_reg_346_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp38_i),
	.data_out(rnode_345to346_bb4_not_cmp38_i_0_reg_346_NO_SHIFT_REG)
);

defparam rnode_345to346_bb4_not_cmp38_i_0_reg_346_fifo.DEPTH = 1;
defparam rnode_345to346_bb4_not_cmp38_i_0_reg_346_fifo.DATA_WIDTH = 1;
defparam rnode_345to346_bb4_not_cmp38_i_0_reg_346_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_345to346_bb4_not_cmp38_i_0_reg_346_fifo.IMPL = "shift_reg";

assign rnode_345to346_bb4_not_cmp38_i_0_reg_346_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp38_i_stall_in_1 = 1'b0;
assign rnode_345to346_bb4_not_cmp38_i_0_NO_SHIFT_REG = rnode_345to346_bb4_not_cmp38_i_0_reg_346_NO_SHIFT_REG;
assign rnode_345to346_bb4_not_cmp38_i_0_stall_in_reg_346_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_399_400_0_inputs_ready;
 reg SFC_3_VALID_399_400_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_399_400_0_stall_in;
wire SFC_3_VALID_399_400_0_output_regs_ready;
 reg SFC_3_VALID_399_400_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_399_400_0_causedstall;

assign SFC_3_VALID_399_400_0_inputs_ready = 1'b1;
assign SFC_3_VALID_399_400_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_398_399_0_stall_in = 1'b0;
assign SFC_3_VALID_399_400_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_399_400_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_399_400_0_output_regs_ready)
		begin
			SFC_3_VALID_399_400_0_NO_SHIFT_REG <= SFC_3_VALID_398_399_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i583_stall_local;
wire local_bb4_notrhs_i583;

assign local_bb4_notrhs_i583 = ((rnode_345to346_bb4_and251_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl274_i_stall_local;
wire [31:0] local_bb4_shl274_i;

assign local_bb4_shl274_i = ((rnode_345to347_bb4_and270_i586_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and248_i_stall_local;
wire [31:0] local_bb4_and248_i;

assign local_bb4_and248_i = (rnode_345to346_bb4_add246_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp259_i_stall_local;
wire local_bb4_cmp259_i;

assign local_bb4_cmp259_i = ($signed(rnode_345to346_bb4_add246_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and226_i_stall_local;
wire [31:0] local_bb4_and226_i;

assign local_bb4_and226_i = ((rnode_345to346_bb4__45_i578_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and271_i_stall_local;
wire [31:0] local_bb4_and271_i;

assign local_bb4_and271_i = ((rnode_345to346_bb4__45_i578_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr272_i_valid_out;
wire local_bb4_shr272_i_stall_in;
wire local_bb4_shr272_i_inputs_ready;
wire local_bb4_shr272_i_stall_local;
wire [31:0] local_bb4_shr272_i;

assign local_bb4_shr272_i_inputs_ready = rnode_345to346_bb4__45_i578_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr272_i = ((rnode_345to346_bb4__45_i578_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr272_i_valid_out = 1'b1;
assign rnode_345to346_bb4__45_i578_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_400_401_0_inputs_ready;
 reg SFC_3_VALID_400_401_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_400_401_0_stall_in;
wire SFC_3_VALID_400_401_0_output_regs_ready;
 reg SFC_3_VALID_400_401_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_400_401_0_causedstall;

assign SFC_3_VALID_400_401_0_inputs_ready = 1'b1;
assign SFC_3_VALID_400_401_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_399_400_0_stall_in = 1'b0;
assign SFC_3_VALID_400_401_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_400_401_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_400_401_0_output_regs_ready)
		begin
			SFC_3_VALID_400_401_0_NO_SHIFT_REG <= SFC_3_VALID_399_400_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i582_stall_local;
wire local_bb4_notlhs_i582;

assign local_bb4_notlhs_i582 = ((local_bb4_and248_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp227_i_stall_local;
wire local_bb4_cmp227_i;

assign local_bb4_cmp227_i = ((local_bb4_and226_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp297_i_stall_local;
wire local_bb4_cmp297_i;

assign local_bb4_cmp297_i = ((local_bb4_and271_i & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp297_i_valid_out;
wire local_bb4_cmp297_i_stall_in;
wire local_bb4_cmp300_i_valid_out;
wire local_bb4_cmp300_i_stall_in;
wire local_bb4_cmp300_i_inputs_ready;
wire local_bb4_cmp300_i_stall_local;
wire local_bb4_cmp300_i;

assign local_bb4_cmp300_i_inputs_ready = rnode_345to346_bb4__45_i578_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp300_i = ((local_bb4_and271_i & 32'h7) == 32'h4);
assign local_bb4_cmp297_i_valid_out = 1'b1;
assign local_bb4_cmp300_i_valid_out = 1'b1;
assign rnode_345to346_bb4__45_i578_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_346to347_bb4_shr272_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_346to347_bb4_shr272_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_346to347_bb4_shr272_i_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4_shr272_i_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_346to347_bb4_shr272_i_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_shr272_i_0_valid_out_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_shr272_i_0_stall_in_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_shr272_i_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_346to347_bb4_shr272_i_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to347_bb4_shr272_i_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to347_bb4_shr272_i_0_stall_in_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_346to347_bb4_shr272_i_0_valid_out_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_346to347_bb4_shr272_i_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in((local_bb4_shr272_i & 32'h1FFFFFF)),
	.data_out(rnode_346to347_bb4_shr272_i_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_346to347_bb4_shr272_i_0_reg_347_fifo.DEPTH = 1;
defparam rnode_346to347_bb4_shr272_i_0_reg_347_fifo.DATA_WIDTH = 32;
defparam rnode_346to347_bb4_shr272_i_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to347_bb4_shr272_i_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_346to347_bb4_shr272_i_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr272_i_stall_in = 1'b0;
assign rnode_346to347_bb4_shr272_i_0_NO_SHIFT_REG = rnode_346to347_bb4_shr272_i_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4_shr272_i_0_stall_in_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_shr272_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_401_402_0_inputs_ready;
 reg SFC_3_VALID_401_402_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_401_402_0_stall_in_0;
 reg SFC_3_VALID_401_402_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_401_402_0_stall_in_1;
wire SFC_3_VALID_401_402_0_output_regs_ready;
 reg SFC_3_VALID_401_402_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_401_402_0_causedstall;

assign SFC_3_VALID_401_402_0_inputs_ready = 1'b1;
assign SFC_3_VALID_401_402_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_400_401_0_stall_in = 1'b0;
assign SFC_3_VALID_401_402_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_401_402_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_401_402_0_output_regs_ready)
		begin
			SFC_3_VALID_401_402_0_NO_SHIFT_REG <= SFC_3_VALID_400_401_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i584_stall_local;
wire local_bb4_not__46_i584;

assign local_bb4_not__46_i584 = (local_bb4_notrhs_i583 | local_bb4_notlhs_i582);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp227_not_i_stall_local;
wire local_bb4_cmp227_not_i;

assign local_bb4_cmp227_not_i = (local_bb4_cmp227_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_346to347_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp297_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp297_i_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp297_i_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp297_i_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp297_i_0_valid_out_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp297_i_0_stall_in_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp297_i_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_346to347_bb4_cmp297_i_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to347_bb4_cmp297_i_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to347_bb4_cmp297_i_0_stall_in_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_346to347_bb4_cmp297_i_0_valid_out_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_346to347_bb4_cmp297_i_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in(local_bb4_cmp297_i),
	.data_out(rnode_346to347_bb4_cmp297_i_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_346to347_bb4_cmp297_i_0_reg_347_fifo.DEPTH = 1;
defparam rnode_346to347_bb4_cmp297_i_0_reg_347_fifo.DATA_WIDTH = 1;
defparam rnode_346to347_bb4_cmp297_i_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to347_bb4_cmp297_i_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_346to347_bb4_cmp297_i_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp297_i_stall_in = 1'b0;
assign rnode_346to347_bb4_cmp297_i_0_NO_SHIFT_REG = rnode_346to347_bb4_cmp297_i_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4_cmp297_i_0_stall_in_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_346to347_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp300_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp300_i_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp300_i_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp300_i_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp300_i_0_valid_out_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp300_i_0_stall_in_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_cmp300_i_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_346to347_bb4_cmp300_i_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to347_bb4_cmp300_i_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to347_bb4_cmp300_i_0_stall_in_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_346to347_bb4_cmp300_i_0_valid_out_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_346to347_bb4_cmp300_i_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in(local_bb4_cmp300_i),
	.data_out(rnode_346to347_bb4_cmp300_i_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_346to347_bb4_cmp300_i_0_reg_347_fifo.DEPTH = 1;
defparam rnode_346to347_bb4_cmp300_i_0_reg_347_fifo.DATA_WIDTH = 1;
defparam rnode_346to347_bb4_cmp300_i_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to347_bb4_cmp300_i_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_346to347_bb4_cmp300_i_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp300_i_stall_in = 1'b0;
assign rnode_346to347_bb4_cmp300_i_0_NO_SHIFT_REG = rnode_346to347_bb4_cmp300_i_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4_cmp300_i_0_stall_in_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and273_i_stall_local;
wire [31:0] local_bb4_and273_i;

assign local_bb4_and273_i = ((rnode_346to347_bb4_shr272_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_402_403_0_inputs_ready;
 reg SFC_3_VALID_402_403_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_402_403_0_stall_in_0;
 reg SFC_3_VALID_402_403_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_402_403_0_stall_in_1;
 reg SFC_3_VALID_402_403_0_valid_out_2_NO_SHIFT_REG;
wire SFC_3_VALID_402_403_0_stall_in_2;
wire SFC_3_VALID_402_403_0_output_regs_ready;
 reg SFC_3_VALID_402_403_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_402_403_0_causedstall;

assign SFC_3_VALID_402_403_0_inputs_ready = 1'b1;
assign SFC_3_VALID_402_403_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_401_402_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_402_403_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_402_403_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_402_403_0_output_regs_ready)
		begin
			SFC_3_VALID_402_403_0_NO_SHIFT_REG <= SFC_3_VALID_401_402_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__47_i585_stall_local;
wire local_bb4__47_i585;

assign local_bb4__47_i585 = (local_bb4_cmp227_i | local_bb4_not__46_i584);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i579_stall_local;
wire local_bb4_brmerge12_i579;

assign local_bb4_brmerge12_i579 = (local_bb4_cmp227_not_i | rnode_345to346_bb4_not_cmp38_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot263__i_stall_local;
wire local_bb4_lnot263__i;

assign local_bb4_lnot263__i = (local_bb4_cmp259_i & local_bb4_cmp227_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29749_i_stall_local;
wire [31:0] local_bb4_cmp29749_i;

assign local_bb4_cmp29749_i[31:1] = 31'h0;
assign local_bb4_cmp29749_i[0] = rnode_346to347_bb4_cmp297_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv301_i_stall_local;
wire [31:0] local_bb4_conv301_i;

assign local_bb4_conv301_i[31:1] = 31'h0;
assign local_bb4_conv301_i[0] = rnode_346to347_bb4_cmp300_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i587_stall_local;
wire [31:0] local_bb4_or275_i587;

assign local_bb4_or275_i587 = ((local_bb4_and273_i & 32'h7FFFFF) | (local_bb4_shl274_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i580_stall_local;
wire [31:0] local_bb4_resultSign_0_i580;

assign local_bb4_resultSign_0_i580 = (local_bb4_brmerge12_i579 ? (rnode_345to346_bb4_and35_i520_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i580_valid_out;
wire local_bb4_resultSign_0_i580_stall_in;
wire local_bb4__47_i585_valid_out;
wire local_bb4__47_i585_stall_in;
wire local_bb4_or2672_i_valid_out;
wire local_bb4_or2672_i_stall_in;
wire local_bb4_or2672_i_inputs_ready;
wire local_bb4_or2672_i_stall_local;
wire local_bb4_or2672_i;

assign local_bb4_or2672_i_inputs_ready = (rnode_345to346_bb4_and35_i520_0_valid_out_NO_SHIFT_REG & rnode_345to346_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG & rnode_345to346_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG & rnode_345to346_bb4_and251_i_0_valid_out_NO_SHIFT_REG & rnode_345to346_bb4__45_i578_0_valid_out_0_NO_SHIFT_REG & rnode_345to346_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG & rnode_345to346_bb4_var__u42_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2672_i = (rnode_345to346_bb4_var__u42_0_NO_SHIFT_REG | local_bb4_lnot263__i);
assign local_bb4_resultSign_0_i580_valid_out = 1'b1;
assign local_bb4__47_i585_valid_out = 1'b1;
assign local_bb4_or2672_i_valid_out = 1'b1;
assign rnode_345to346_bb4_and35_i520_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_not_cmp38_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_add246_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_and251_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4__45_i578_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_add246_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_345to346_bb4_var__u42_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_346to347_bb4_resultSign_0_i580_0_valid_out_NO_SHIFT_REG;
 logic rnode_346to347_bb4_resultSign_0_i580_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_346to347_bb4_resultSign_0_i580_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4_resultSign_0_i580_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_346to347_bb4_resultSign_0_i580_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_resultSign_0_i580_0_valid_out_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_resultSign_0_i580_0_stall_in_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_resultSign_0_i580_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_346to347_bb4_resultSign_0_i580_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to347_bb4_resultSign_0_i580_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to347_bb4_resultSign_0_i580_0_stall_in_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_346to347_bb4_resultSign_0_i580_0_valid_out_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_346to347_bb4_resultSign_0_i580_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i580 & 32'h80000000)),
	.data_out(rnode_346to347_bb4_resultSign_0_i580_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_346to347_bb4_resultSign_0_i580_0_reg_347_fifo.DEPTH = 1;
defparam rnode_346to347_bb4_resultSign_0_i580_0_reg_347_fifo.DATA_WIDTH = 32;
defparam rnode_346to347_bb4_resultSign_0_i580_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to347_bb4_resultSign_0_i580_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_346to347_bb4_resultSign_0_i580_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i580_stall_in = 1'b0;
assign rnode_346to347_bb4_resultSign_0_i580_0_NO_SHIFT_REG = rnode_346to347_bb4_resultSign_0_i580_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4_resultSign_0_i580_0_stall_in_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_resultSign_0_i580_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_346to347_bb4__47_i585_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_valid_out_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_stall_in_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4__47_i585_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_346to347_bb4__47_i585_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to347_bb4__47_i585_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to347_bb4__47_i585_0_stall_in_0_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_346to347_bb4__47_i585_0_valid_out_0_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_346to347_bb4__47_i585_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in(local_bb4__47_i585),
	.data_out(rnode_346to347_bb4__47_i585_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_346to347_bb4__47_i585_0_reg_347_fifo.DEPTH = 1;
defparam rnode_346to347_bb4__47_i585_0_reg_347_fifo.DATA_WIDTH = 1;
defparam rnode_346to347_bb4__47_i585_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to347_bb4__47_i585_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_346to347_bb4__47_i585_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i585_stall_in = 1'b0;
assign rnode_346to347_bb4__47_i585_0_stall_in_0_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__47_i585_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4__47_i585_0_NO_SHIFT_REG = rnode_346to347_bb4__47_i585_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4__47_i585_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4__47_i585_1_NO_SHIFT_REG = rnode_346to347_bb4__47_i585_0_reg_347_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_346to347_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_1_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_2_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_reg_347_inputs_ready_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_valid_out_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_stall_in_0_reg_347_NO_SHIFT_REG;
 logic rnode_346to347_bb4_or2672_i_0_stall_out_reg_347_NO_SHIFT_REG;

acl_data_fifo rnode_346to347_bb4_or2672_i_0_reg_347_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_346to347_bb4_or2672_i_0_reg_347_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_346to347_bb4_or2672_i_0_stall_in_0_reg_347_NO_SHIFT_REG),
	.valid_out(rnode_346to347_bb4_or2672_i_0_valid_out_0_reg_347_NO_SHIFT_REG),
	.stall_out(rnode_346to347_bb4_or2672_i_0_stall_out_reg_347_NO_SHIFT_REG),
	.data_in(local_bb4_or2672_i),
	.data_out(rnode_346to347_bb4_or2672_i_0_reg_347_NO_SHIFT_REG)
);

defparam rnode_346to347_bb4_or2672_i_0_reg_347_fifo.DEPTH = 1;
defparam rnode_346to347_bb4_or2672_i_0_reg_347_fifo.DATA_WIDTH = 1;
defparam rnode_346to347_bb4_or2672_i_0_reg_347_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_346to347_bb4_or2672_i_0_reg_347_fifo.IMPL = "shift_reg";

assign rnode_346to347_bb4_or2672_i_0_reg_347_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2672_i_stall_in = 1'b0;
assign rnode_346to347_bb4_or2672_i_0_stall_in_0_reg_347_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4_or2672_i_0_NO_SHIFT_REG = rnode_346to347_bb4_or2672_i_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4_or2672_i_1_NO_SHIFT_REG = rnode_346to347_bb4_or2672_i_0_reg_347_NO_SHIFT_REG;
assign rnode_346to347_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_346to347_bb4_or2672_i_2_NO_SHIFT_REG = rnode_346to347_bb4_or2672_i_0_reg_347_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or276_i_stall_local;
wire [31:0] local_bb4_or276_i;

assign local_bb4_or276_i = ((local_bb4_or275_i587 & 32'h7FFFFFFF) | (rnode_346to347_bb4_resultSign_0_i580_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u54_stall_local;
wire [31:0] local_bb4_var__u54;

assign local_bb4_var__u54[31:1] = 31'h0;
assign local_bb4_var__u54[0] = rnode_346to347_bb4__47_i585_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2814_i_stall_local;
wire local_bb4_or2814_i;

assign local_bb4_or2814_i = (rnode_346to347_bb4__47_i585_0_NO_SHIFT_REG | rnode_346to347_bb4_or2672_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2885_i_stall_local;
wire local_bb4_or2885_i;

assign local_bb4_or2885_i = (rnode_346to347_bb4_or2672_i_1_NO_SHIFT_REG | rnode_346to347_bb4__26_i533_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u55_stall_local;
wire [31:0] local_bb4_var__u55;

assign local_bb4_var__u55[31:1] = 31'h0;
assign local_bb4_var__u55[0] = rnode_346to347_bb4_or2672_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext315_i_stall_local;
wire [31:0] local_bb4_lnot_ext315_i;

assign local_bb4_lnot_ext315_i = ((local_bb4_var__u54 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond283_i_stall_local;
wire [31:0] local_bb4_cond283_i;

assign local_bb4_cond283_i = (local_bb4_or2814_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond290_i_stall_local;
wire [31:0] local_bb4_cond290_i;

assign local_bb4_cond290_i = (local_bb4_or2885_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext311_i_stall_local;
wire [31:0] local_bb4_lnot_ext311_i;

assign local_bb4_lnot_ext311_i = ((local_bb4_var__u55 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and294_i_stall_local;
wire [31:0] local_bb4_and294_i;

assign local_bb4_and294_i = ((local_bb4_cond283_i | 32'h80000000) & local_bb4_or276_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i588_stall_local;
wire [31:0] local_bb4_or295_i588;

assign local_bb4_or295_i588 = ((local_bb4_cond290_i & 32'h7F800000) | (local_bb4_cond293_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i591_stall_local;
wire [31:0] local_bb4_reduction_0_i591;

assign local_bb4_reduction_0_i591 = ((local_bb4_lnot_ext311_i & 32'h1) & (local_bb4_lnot_ext_i590 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and303_i_stall_local;
wire [31:0] local_bb4_and303_i;

assign local_bb4_and303_i = ((local_bb4_conv301_i & 32'h1) & local_bb4_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or296_i_stall_local;
wire [31:0] local_bb4_or296_i;

assign local_bb4_or296_i = ((local_bb4_or295_i588 & 32'h7FC00000) | local_bb4_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i589_stall_local;
wire [31:0] local_bb4_lor_ext_i589;

assign local_bb4_lor_ext_i589 = ((local_bb4_cmp29749_i & 32'h1) | (local_bb4_and303_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i592_stall_local;
wire [31:0] local_bb4_reduction_1_i592;

assign local_bb4_reduction_1_i592 = ((local_bb4_lnot_ext315_i & 32'h1) & (local_bb4_lor_ext_i589 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i593_stall_local;
wire [31:0] local_bb4_reduction_2_i593;

assign local_bb4_reduction_2_i593 = ((local_bb4_reduction_0_i591 & 32'h1) & (local_bb4_reduction_1_i592 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_add321_i_stall_local;
wire [31:0] local_bb4_add321_i;

assign local_bb4_add321_i = ((local_bb4_reduction_2_i593 & 32'h1) + local_bb4_or296_i);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i404_stall_local;
wire [31:0] local_bb4_shr_i404;

assign local_bb4_shr_i404 = (local_bb4_add321_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i406_stall_local;
wire [31:0] local_bb4_shr2_i406;

assign local_bb4_shr2_i406 = (local_bb4_add321_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and5_i410_stall_local;
wire [31:0] local_bb4_and5_i410;

assign local_bb4_and5_i410 = (local_bb4_add321_i & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and6_i411_stall_local;
wire [31:0] local_bb4_and6_i411;

assign local_bb4_and6_i411 = (local_bb4_add321_i & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i438_stall_local;
wire [31:0] local_bb4_or_i438;

assign local_bb4_or_i438 = ((local_bb4_and5_i410 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_or47_i439_stall_local;
wire [31:0] local_bb4_or47_i439;

assign local_bb4_or47_i439 = ((local_bb4_and6_i411 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_conv_i_i440_stall_local;
wire [63:0] local_bb4_conv_i_i440;

assign local_bb4_conv_i_i440[63:32] = 32'h0;
assign local_bb4_conv_i_i440[31:0] = ((local_bb4_or_i438 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i404_valid_out;
wire local_bb4_shr_i404_stall_in;
wire local_bb4_shr2_i406_valid_out;
wire local_bb4_shr2_i406_stall_in;
wire local_bb4_and5_i410_valid_out_1;
wire local_bb4_and5_i410_stall_in_1;
wire local_bb4_and6_i411_valid_out_1;
wire local_bb4_and6_i411_stall_in_1;
wire local_bb4_conv_i_i440_valid_out;
wire local_bb4_conv_i_i440_stall_in;
wire local_bb4_conv1_i_i441_valid_out;
wire local_bb4_conv1_i_i441_stall_in;
wire local_bb4_conv1_i_i441_inputs_ready;
wire local_bb4_conv1_i_i441_stall_local;
wire [63:0] local_bb4_conv1_i_i441;

assign local_bb4_conv1_i_i441_inputs_ready = (rnode_345to347_bb4_and270_i586_0_valid_out_NO_SHIFT_REG & rnode_346to347_bb4_resultSign_0_i580_0_valid_out_NO_SHIFT_REG & rnode_346to347_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG & rnode_346to347_bb4__26_i533_0_valid_out_0_NO_SHIFT_REG & rnode_346to347_bb4__26_i533_0_valid_out_1_NO_SHIFT_REG & rnode_346to347_bb4__47_i585_0_valid_out_0_NO_SHIFT_REG & rnode_346to347_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG & rnode_346to347_bb4__26_i533_0_valid_out_2_NO_SHIFT_REG & rnode_346to347_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG & rnode_346to347_bb4_shr272_i_0_valid_out_NO_SHIFT_REG & rnode_346to347_bb4__47_i585_0_valid_out_1_NO_SHIFT_REG & rnode_346to347_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG & rnode_346to347_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_conv1_i_i441[63:32] = 32'h0;
assign local_bb4_conv1_i_i441[31:0] = ((local_bb4_or47_i439 & 32'hFFFFFF) | 32'h800000);
assign local_bb4_shr_i404_valid_out = 1'b1;
assign local_bb4_shr2_i406_valid_out = 1'b1;
assign local_bb4_and5_i410_valid_out_1 = 1'b1;
assign local_bb4_and6_i411_valid_out_1 = 1'b1;
assign local_bb4_conv_i_i440_valid_out = 1'b1;
assign local_bb4_conv1_i_i441_valid_out = 1'b1;
assign rnode_345to347_bb4_and270_i586_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_resultSign_0_i580_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_or2672_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__26_i533_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__26_i533_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__47_i585_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_or2672_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__26_i533_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_or2672_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_shr272_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4__47_i585_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_cmp297_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_346to347_bb4_cmp300_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_347to348_bb4_shr_i404_0_valid_out_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr_i404_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_shr_i404_0_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr_i404_0_reg_348_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_shr_i404_0_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr_i404_0_valid_out_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr_i404_0_stall_in_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr_i404_0_stall_out_reg_348_NO_SHIFT_REG;

acl_data_fifo rnode_347to348_bb4_shr_i404_0_reg_348_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_347to348_bb4_shr_i404_0_reg_348_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_347to348_bb4_shr_i404_0_stall_in_reg_348_NO_SHIFT_REG),
	.valid_out(rnode_347to348_bb4_shr_i404_0_valid_out_reg_348_NO_SHIFT_REG),
	.stall_out(rnode_347to348_bb4_shr_i404_0_stall_out_reg_348_NO_SHIFT_REG),
	.data_in((local_bb4_shr_i404 & 32'h1FF)),
	.data_out(rnode_347to348_bb4_shr_i404_0_reg_348_NO_SHIFT_REG)
);

defparam rnode_347to348_bb4_shr_i404_0_reg_348_fifo.DEPTH = 1;
defparam rnode_347to348_bb4_shr_i404_0_reg_348_fifo.DATA_WIDTH = 32;
defparam rnode_347to348_bb4_shr_i404_0_reg_348_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_347to348_bb4_shr_i404_0_reg_348_fifo.IMPL = "shift_reg";

assign rnode_347to348_bb4_shr_i404_0_reg_348_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr_i404_stall_in = 1'b0;
assign rnode_347to348_bb4_shr_i404_0_NO_SHIFT_REG = rnode_347to348_bb4_shr_i404_0_reg_348_NO_SHIFT_REG;
assign rnode_347to348_bb4_shr_i404_0_stall_in_reg_348_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_shr_i404_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_347to348_bb4_shr2_i406_0_valid_out_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr2_i406_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_shr2_i406_0_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr2_i406_0_reg_348_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_shr2_i406_0_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr2_i406_0_valid_out_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr2_i406_0_stall_in_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_shr2_i406_0_stall_out_reg_348_NO_SHIFT_REG;

acl_data_fifo rnode_347to348_bb4_shr2_i406_0_reg_348_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_347to348_bb4_shr2_i406_0_reg_348_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_347to348_bb4_shr2_i406_0_stall_in_reg_348_NO_SHIFT_REG),
	.valid_out(rnode_347to348_bb4_shr2_i406_0_valid_out_reg_348_NO_SHIFT_REG),
	.stall_out(rnode_347to348_bb4_shr2_i406_0_stall_out_reg_348_NO_SHIFT_REG),
	.data_in((local_bb4_shr2_i406 & 32'h1FF)),
	.data_out(rnode_347to348_bb4_shr2_i406_0_reg_348_NO_SHIFT_REG)
);

defparam rnode_347to348_bb4_shr2_i406_0_reg_348_fifo.DEPTH = 1;
defparam rnode_347to348_bb4_shr2_i406_0_reg_348_fifo.DATA_WIDTH = 32;
defparam rnode_347to348_bb4_shr2_i406_0_reg_348_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_347to348_bb4_shr2_i406_0_reg_348_fifo.IMPL = "shift_reg";

assign rnode_347to348_bb4_shr2_i406_0_reg_348_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr2_i406_stall_in = 1'b0;
assign rnode_347to348_bb4_shr2_i406_0_NO_SHIFT_REG = rnode_347to348_bb4_shr2_i406_0_reg_348_NO_SHIFT_REG;
assign rnode_347to348_bb4_shr2_i406_0_stall_in_reg_348_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_shr2_i406_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_347to348_bb4_and5_i410_0_valid_out_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and5_i410_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_and5_i410_0_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and5_i410_0_reg_348_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_and5_i410_0_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and5_i410_0_valid_out_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and5_i410_0_stall_in_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and5_i410_0_stall_out_reg_348_NO_SHIFT_REG;

acl_data_fifo rnode_347to348_bb4_and5_i410_0_reg_348_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_347to348_bb4_and5_i410_0_reg_348_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_347to348_bb4_and5_i410_0_stall_in_reg_348_NO_SHIFT_REG),
	.valid_out(rnode_347to348_bb4_and5_i410_0_valid_out_reg_348_NO_SHIFT_REG),
	.stall_out(rnode_347to348_bb4_and5_i410_0_stall_out_reg_348_NO_SHIFT_REG),
	.data_in((local_bb4_and5_i410 & 32'h7FFFFF)),
	.data_out(rnode_347to348_bb4_and5_i410_0_reg_348_NO_SHIFT_REG)
);

defparam rnode_347to348_bb4_and5_i410_0_reg_348_fifo.DEPTH = 1;
defparam rnode_347to348_bb4_and5_i410_0_reg_348_fifo.DATA_WIDTH = 32;
defparam rnode_347to348_bb4_and5_i410_0_reg_348_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_347to348_bb4_and5_i410_0_reg_348_fifo.IMPL = "shift_reg";

assign rnode_347to348_bb4_and5_i410_0_reg_348_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and5_i410_stall_in_1 = 1'b0;
assign rnode_347to348_bb4_and5_i410_0_NO_SHIFT_REG = rnode_347to348_bb4_and5_i410_0_reg_348_NO_SHIFT_REG;
assign rnode_347to348_bb4_and5_i410_0_stall_in_reg_348_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_and5_i410_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_347to348_bb4_and6_i411_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_and6_i411_0_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_and6_i411_1_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_and6_i411_2_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_reg_348_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_347to348_bb4_and6_i411_0_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_valid_out_0_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_stall_in_0_reg_348_NO_SHIFT_REG;
 logic rnode_347to348_bb4_and6_i411_0_stall_out_reg_348_NO_SHIFT_REG;

acl_data_fifo rnode_347to348_bb4_and6_i411_0_reg_348_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_347to348_bb4_and6_i411_0_reg_348_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_347to348_bb4_and6_i411_0_stall_in_0_reg_348_NO_SHIFT_REG),
	.valid_out(rnode_347to348_bb4_and6_i411_0_valid_out_0_reg_348_NO_SHIFT_REG),
	.stall_out(rnode_347to348_bb4_and6_i411_0_stall_out_reg_348_NO_SHIFT_REG),
	.data_in((local_bb4_and6_i411 & 32'h7FFFFF)),
	.data_out(rnode_347to348_bb4_and6_i411_0_reg_348_NO_SHIFT_REG)
);

defparam rnode_347to348_bb4_and6_i411_0_reg_348_fifo.DEPTH = 1;
defparam rnode_347to348_bb4_and6_i411_0_reg_348_fifo.DATA_WIDTH = 32;
defparam rnode_347to348_bb4_and6_i411_0_reg_348_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_347to348_bb4_and6_i411_0_reg_348_fifo.IMPL = "shift_reg";

assign rnode_347to348_bb4_and6_i411_0_reg_348_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and6_i411_stall_in_1 = 1'b0;
assign rnode_347to348_bb4_and6_i411_0_stall_in_0_reg_348_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_and6_i411_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_347to348_bb4_and6_i411_0_NO_SHIFT_REG = rnode_347to348_bb4_and6_i411_0_reg_348_NO_SHIFT_REG;
assign rnode_347to348_bb4_and6_i411_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_347to348_bb4_and6_i411_1_NO_SHIFT_REG = rnode_347to348_bb4_and6_i411_0_reg_348_NO_SHIFT_REG;
assign rnode_347to348_bb4_and6_i411_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_347to348_bb4_and6_i411_2_NO_SHIFT_REG = rnode_347to348_bb4_and6_i411_0_reg_348_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_mul_i_i442_inputs_ready;
 reg local_bb4_mul_i_i442_valid_out_0_NO_SHIFT_REG;
wire local_bb4_mul_i_i442_stall_in_0;
 reg local_bb4_mul_i_i442_valid_out_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i442_stall_in_1;
wire local_bb4_mul_i_i442_output_regs_ready;
wire [63:0] local_bb4_mul_i_i442;
 reg local_bb4_mul_i_i442_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul_i_i442_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i442_causedstall;

acl_int_mult int_module_local_bb4_mul_i_i442 (
	.clock(clock),
	.dataa(((local_bb4_conv1_i_i441 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb4_conv_i_i440 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb4_mul_i_i442_output_regs_ready),
	.result(local_bb4_mul_i_i442)
);

defparam int_module_local_bb4_mul_i_i442.INPUT1_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i442.INPUT2_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i442.OUTPUT_WIDTH = 64;
defparam int_module_local_bb4_mul_i_i442.LATENCY = 3;
defparam int_module_local_bb4_mul_i_i442.SIGNED = 0;

assign local_bb4_mul_i_i442_inputs_ready = 1'b1;
assign local_bb4_mul_i_i442_output_regs_ready = 1'b1;
assign local_bb4_conv1_i_i441_stall_in = 1'b0;
assign local_bb4_conv_i_i440_stall_in = 1'b0;
assign local_bb4_mul_i_i442_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i442_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i442_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i442_output_regs_ready)
		begin
			local_bb4_mul_i_i442_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i442_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul_i_i442_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i442_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i442_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i442_output_regs_ready)
		begin
			local_bb4_mul_i_i442_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i442_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul_i_i442_stall_in_0))
			begin
				local_bb4_mul_i_i442_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_mul_i_i442_stall_in_1))
			begin
				local_bb4_mul_i_i442_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and_i405_stall_local;
wire [31:0] local_bb4_and_i405;

assign local_bb4_and_i405 = ((rnode_347to348_bb4_shr_i404_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and3_i407_stall_local;
wire [31:0] local_bb4_and3_i407;

assign local_bb4_and3_i407 = ((rnode_347to348_bb4_shr2_i406_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i416_stall_local;
wire local_bb4_lnot14_i416;

assign local_bb4_lnot14_i416 = ((rnode_347to348_bb4_and5_i410_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_i417_stall_local;
wire local_bb4_lnot17_i417;

assign local_bb4_lnot17_i417 = ((rnode_347to348_bb4_and6_i411_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_conv3_i_i443_stall_local;
wire [31:0] local_bb4_conv3_i_i443;
wire [63:0] local_bb4_conv3_i_i443$ps;

assign local_bb4_conv3_i_i443$ps = (local_bb4_mul_i_i442 & 64'hFFFFFFFFFFFF);
assign local_bb4_conv3_i_i443 = local_bb4_conv3_i_i443$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u56_stall_local;
wire [63:0] local_bb4_var__u56;

assign local_bb4_var__u56 = ((local_bb4_mul_i_i442 & 64'hFFFFFFFFFFFF) >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i412_stall_local;
wire local_bb4_lnot_i412;

assign local_bb4_lnot_i412 = ((local_bb4_and_i405 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i414_stall_local;
wire local_bb4_cmp_i414;

assign local_bb4_cmp_i414 = ((local_bb4_and_i405 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u57_stall_local;
wire [31:0] local_bb4_var__u57;

assign local_bb4_var__u57 = ((rnode_347to348_bb4_and6_i411_2_NO_SHIFT_REG & 32'h7FFFFF) | (local_bb4_and_i405 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot8_i413_stall_local;
wire local_bb4_lnot8_i413;

assign local_bb4_lnot8_i413 = ((local_bb4_and3_i407 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_i415_stall_local;
wire local_bb4_cmp11_i415;

assign local_bb4_cmp11_i415 = ((local_bb4_and3_i407 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u58_stall_local;
wire [31:0] local_bb4_var__u58;

assign local_bb4_var__u58 = ((local_bb4_and3_i407 & 32'hFF) | (rnode_347to348_bb4_and6_i411_1_NO_SHIFT_REG & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i449_stall_local;
wire [31:0] local_bb4_add_i449;

assign local_bb4_add_i449 = ((local_bb4_and3_i407 & 32'hFF) + (local_bb4_and_i405 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_not_i435_stall_local;
wire local_bb4_lnot14_not_i435;

assign local_bb4_lnot14_not_i435 = (local_bb4_lnot14_i416 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_not_i421_stall_local;
wire local_bb4_lnot17_not_i421;

assign local_bb4_lnot17_not_i421 = (local_bb4_lnot17_i417 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i16_i446_stall_local;
wire [31:0] local_bb4_shr_i16_i446;

assign local_bb4_shr_i16_i446 = (local_bb4_conv3_i_i443 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i18_i448_stall_local;
wire [31:0] local_bb4_shl1_i18_i448;

assign local_bb4_shl1_i18_i448 = (local_bb4_conv3_i_i443 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u59_stall_local;
wire [31:0] local_bb4_var__u59;

assign local_bb4_var__u59 = (local_bb4_conv3_i_i443 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i_i456_stall_local;
wire [31:0] local_bb4_shl1_i_i456;

assign local_bb4_shl1_i_i456 = (local_bb4_conv3_i_i443 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb4__tr_i444_stall_local;
wire [31:0] local_bb4__tr_i444;
wire [63:0] local_bb4__tr_i444$ps;

assign local_bb4__tr_i444$ps = (local_bb4_var__u56 & 64'hFFFFFF);
assign local_bb4__tr_i444 = local_bb4__tr_i444$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u60_stall_local;
wire local_bb4_var__u60;

assign local_bb4_var__u60 = ((local_bb4_var__u57 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i467_stall_local;
wire local_bb4_reduction_0_i467;

assign local_bb4_reduction_0_i467 = (local_bb4_lnot_i412 | local_bb4_lnot8_i413);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge8_demorgan_i418_stall_local;
wire local_bb4_brmerge8_demorgan_i418;

assign local_bb4_brmerge8_demorgan_i418 = (local_bb4_cmp11_i415 & local_bb4_lnot17_i417);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_not_i422_stall_local;
wire local_bb4_cmp11_not_i422;

assign local_bb4_cmp11_not_i422 = (local_bb4_cmp11_i415 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u61_stall_local;
wire local_bb4_var__u61;

assign local_bb4_var__u61 = (local_bb4_cmp_i414 | local_bb4_cmp11_i415);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u62_stall_local;
wire local_bb4_var__u62;

assign local_bb4_var__u62 = ((local_bb4_var__u58 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i436_stall_local;
wire local_bb4__28_i436;

assign local_bb4__28_i436 = (local_bb4_cmp_i414 & local_bb4_lnot14_not_i435);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i454_stall_local;
wire [31:0] local_bb4_shr_i_i454;

assign local_bb4_shr_i_i454 = ((local_bb4_var__u59 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i15_i445_stall_local;
wire [31:0] local_bb4_shl_i15_i445;

assign local_bb4_shl_i15_i445 = ((local_bb4__tr_i444 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb4_and48_i450_stall_local;
wire [31:0] local_bb4_and48_i450;

assign local_bb4_and48_i450 = ((local_bb4__tr_i444 & 32'hFFFFFF) & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge10_demorgan_i419_stall_local;
wire local_bb4_brmerge10_demorgan_i419;

assign local_bb4_brmerge10_demorgan_i419 = (local_bb4_brmerge8_demorgan_i418 & local_bb4_lnot_i412);

// This section implements an unregistered operation.
// 
wire local_bb4__mux9_mux_i420_stall_local;
wire local_bb4__mux9_mux_i420;

assign local_bb4__mux9_mux_i420 = (local_bb4_brmerge8_demorgan_i418 ^ local_bb4_cmp11_i415);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge3_i423_stall_local;
wire local_bb4_brmerge3_i423;

assign local_bb4_brmerge3_i423 = (local_bb4_var__u62 | local_bb4_cmp11_not_i422);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_i425_stall_local;
wire local_bb4__mux_mux_i425;

assign local_bb4__mux_mux_i425 = (local_bb4_var__u62 | local_bb4_cmp11_i415);

// This section implements an unregistered operation.
// 
wire local_bb4__not_i427_stall_local;
wire local_bb4__not_i427;

assign local_bb4__not_i427 = (local_bb4_var__u62 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i17_i447_stall_local;
wire [31:0] local_bb4_or_i17_i447;

assign local_bb4_or_i17_i447 = ((local_bb4_shl_i15_i445 & 32'hFFFF00) | (local_bb4_shr_i16_i446 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool49_i451_stall_local;
wire local_bb4_tobool49_i451;

assign local_bb4_tobool49_i451 = ((local_bb4_and48_i450 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__26_demorgan_i433_stall_local;
wire local_bb4__26_demorgan_i433;

assign local_bb4__26_demorgan_i433 = (local_bb4_cmp_i414 | local_bb4_brmerge10_demorgan_i419);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge5_i424_stall_local;
wire local_bb4_brmerge5_i424;

assign local_bb4_brmerge5_i424 = (local_bb4_brmerge3_i423 | local_bb4_lnot17_not_i421);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i428_stall_local;
wire local_bb4_reduction_3_i428;

assign local_bb4_reduction_3_i428 = (local_bb4_cmp11_i415 & local_bb4__not_i427);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_i453_stall_local;
wire [31:0] local_bb4_shl_i_i453;

assign local_bb4_shl_i_i453 = ((local_bb4_or_i17_i447 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_mux_i426_stall_local;
wire local_bb4__mux_mux_mux_i426;

assign local_bb4__mux_mux_mux_i426 = (local_bb4_brmerge5_i424 & local_bb4__mux_mux_i425);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i429_stall_local;
wire local_bb4_reduction_5_i429;

assign local_bb4_reduction_5_i429 = (local_bb4_lnot14_i416 & local_bb4_reduction_3_i428);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i455_stall_local;
wire [31:0] local_bb4_or_i_i455;

assign local_bb4_or_i_i455 = ((local_bb4_shl_i_i453 & 32'h1FFFFFE) | (local_bb4_shr_i_i454 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i430_stall_local;
wire local_bb4_reduction_6_i430;

assign local_bb4_reduction_6_i430 = (local_bb4_var__u60 & local_bb4_reduction_5_i429);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i431_stall_local;
wire local_bb4__24_i431;

assign local_bb4__24_i431 = (local_bb4_cmp_i414 ? local_bb4_reduction_6_i430 : local_bb4_brmerge10_demorgan_i419);

// This section implements an unregistered operation.
// 
wire local_bb4__25_i432_stall_local;
wire local_bb4__25_i432;

assign local_bb4__25_i432 = (local_bb4__24_i431 ? local_bb4_lnot14_i416 : local_bb4__mux_mux_mux_i426);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i434_stall_local;
wire local_bb4__27_i434;

assign local_bb4__27_i434 = (local_bb4__26_demorgan_i433 ? local_bb4__25_i432 : local_bb4__mux9_mux_i420);

// This section implements an unregistered operation.
// 
wire local_bb4_add_i449_valid_out;
wire local_bb4_add_i449_stall_in;
wire local_bb4_reduction_0_i467_valid_out;
wire local_bb4_reduction_0_i467_stall_in;
wire local_bb4_var__u61_valid_out;
wire local_bb4_var__u61_stall_in;
wire local_bb4__29_i437_valid_out;
wire local_bb4__29_i437_stall_in;
wire local_bb4__29_i437_inputs_ready;
wire local_bb4__29_i437_stall_local;
wire local_bb4__29_i437;

assign local_bb4__29_i437_inputs_ready = (rnode_347to348_bb4_shr_i404_0_valid_out_NO_SHIFT_REG & rnode_347to348_bb4_and6_i411_0_valid_out_2_NO_SHIFT_REG & rnode_347to348_bb4_shr2_i406_0_valid_out_NO_SHIFT_REG & rnode_347to348_bb4_and6_i411_0_valid_out_1_NO_SHIFT_REG & rnode_347to348_bb4_and6_i411_0_valid_out_0_NO_SHIFT_REG & rnode_347to348_bb4_and5_i410_0_valid_out_NO_SHIFT_REG);
assign local_bb4__29_i437 = (local_bb4__28_i436 | local_bb4__27_i434);
assign local_bb4_add_i449_valid_out = 1'b1;
assign local_bb4_reduction_0_i467_valid_out = 1'b1;
assign local_bb4_var__u61_valid_out = 1'b1;
assign local_bb4__29_i437_valid_out = 1'b1;
assign rnode_347to348_bb4_shr_i404_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_and6_i411_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_shr2_i406_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_and6_i411_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_and6_i411_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_347to348_bb4_and5_i410_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_348to350_bb4_add_i449_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_348to350_bb4_add_i449_0_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_348to350_bb4_add_i449_1_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_348to350_bb4_add_i449_2_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_reg_350_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_348to350_bb4_add_i449_0_reg_350_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_valid_out_0_reg_350_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_stall_in_0_reg_350_NO_SHIFT_REG;
 logic rnode_348to350_bb4_add_i449_0_stall_out_reg_350_NO_SHIFT_REG;

acl_data_fifo rnode_348to350_bb4_add_i449_0_reg_350_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_348to350_bb4_add_i449_0_reg_350_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_348to350_bb4_add_i449_0_stall_in_0_reg_350_NO_SHIFT_REG),
	.valid_out(rnode_348to350_bb4_add_i449_0_valid_out_0_reg_350_NO_SHIFT_REG),
	.stall_out(rnode_348to350_bb4_add_i449_0_stall_out_reg_350_NO_SHIFT_REG),
	.data_in((local_bb4_add_i449 & 32'h1FF)),
	.data_out(rnode_348to350_bb4_add_i449_0_reg_350_NO_SHIFT_REG)
);

defparam rnode_348to350_bb4_add_i449_0_reg_350_fifo.DEPTH = 2;
defparam rnode_348to350_bb4_add_i449_0_reg_350_fifo.DATA_WIDTH = 32;
defparam rnode_348to350_bb4_add_i449_0_reg_350_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_348to350_bb4_add_i449_0_reg_350_fifo.IMPL = "shift_reg";

assign rnode_348to350_bb4_add_i449_0_reg_350_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add_i449_stall_in = 1'b0;
assign rnode_348to350_bb4_add_i449_0_stall_in_0_reg_350_NO_SHIFT_REG = 1'b0;
assign rnode_348to350_bb4_add_i449_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_348to350_bb4_add_i449_0_NO_SHIFT_REG = rnode_348to350_bb4_add_i449_0_reg_350_NO_SHIFT_REG;
assign rnode_348to350_bb4_add_i449_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_348to350_bb4_add_i449_1_NO_SHIFT_REG = rnode_348to350_bb4_add_i449_0_reg_350_NO_SHIFT_REG;
assign rnode_348to350_bb4_add_i449_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_348to350_bb4_add_i449_2_NO_SHIFT_REG = rnode_348to350_bb4_add_i449_0_reg_350_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_348to349_bb4_reduction_0_i467_0_valid_out_NO_SHIFT_REG;
 logic rnode_348to349_bb4_reduction_0_i467_0_stall_in_NO_SHIFT_REG;
 logic rnode_348to349_bb4_reduction_0_i467_0_NO_SHIFT_REG;
 logic rnode_348to349_bb4_reduction_0_i467_0_reg_349_inputs_ready_NO_SHIFT_REG;
 logic rnode_348to349_bb4_reduction_0_i467_0_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4_reduction_0_i467_0_valid_out_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4_reduction_0_i467_0_stall_in_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4_reduction_0_i467_0_stall_out_reg_349_NO_SHIFT_REG;

acl_data_fifo rnode_348to349_bb4_reduction_0_i467_0_reg_349_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_348to349_bb4_reduction_0_i467_0_reg_349_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_348to349_bb4_reduction_0_i467_0_stall_in_reg_349_NO_SHIFT_REG),
	.valid_out(rnode_348to349_bb4_reduction_0_i467_0_valid_out_reg_349_NO_SHIFT_REG),
	.stall_out(rnode_348to349_bb4_reduction_0_i467_0_stall_out_reg_349_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_0_i467),
	.data_out(rnode_348to349_bb4_reduction_0_i467_0_reg_349_NO_SHIFT_REG)
);

defparam rnode_348to349_bb4_reduction_0_i467_0_reg_349_fifo.DEPTH = 1;
defparam rnode_348to349_bb4_reduction_0_i467_0_reg_349_fifo.DATA_WIDTH = 1;
defparam rnode_348to349_bb4_reduction_0_i467_0_reg_349_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_348to349_bb4_reduction_0_i467_0_reg_349_fifo.IMPL = "shift_reg";

assign rnode_348to349_bb4_reduction_0_i467_0_reg_349_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_0_i467_stall_in = 1'b0;
assign rnode_348to349_bb4_reduction_0_i467_0_NO_SHIFT_REG = rnode_348to349_bb4_reduction_0_i467_0_reg_349_NO_SHIFT_REG;
assign rnode_348to349_bb4_reduction_0_i467_0_stall_in_reg_349_NO_SHIFT_REG = 1'b0;
assign rnode_348to349_bb4_reduction_0_i467_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_348to349_bb4_var__u61_0_valid_out_NO_SHIFT_REG;
 logic rnode_348to349_bb4_var__u61_0_stall_in_NO_SHIFT_REG;
 logic rnode_348to349_bb4_var__u61_0_NO_SHIFT_REG;
 logic rnode_348to349_bb4_var__u61_0_reg_349_inputs_ready_NO_SHIFT_REG;
 logic rnode_348to349_bb4_var__u61_0_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4_var__u61_0_valid_out_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4_var__u61_0_stall_in_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4_var__u61_0_stall_out_reg_349_NO_SHIFT_REG;

acl_data_fifo rnode_348to349_bb4_var__u61_0_reg_349_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_348to349_bb4_var__u61_0_reg_349_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_348to349_bb4_var__u61_0_stall_in_reg_349_NO_SHIFT_REG),
	.valid_out(rnode_348to349_bb4_var__u61_0_valid_out_reg_349_NO_SHIFT_REG),
	.stall_out(rnode_348to349_bb4_var__u61_0_stall_out_reg_349_NO_SHIFT_REG),
	.data_in(local_bb4_var__u61),
	.data_out(rnode_348to349_bb4_var__u61_0_reg_349_NO_SHIFT_REG)
);

defparam rnode_348to349_bb4_var__u61_0_reg_349_fifo.DEPTH = 1;
defparam rnode_348to349_bb4_var__u61_0_reg_349_fifo.DATA_WIDTH = 1;
defparam rnode_348to349_bb4_var__u61_0_reg_349_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_348to349_bb4_var__u61_0_reg_349_fifo.IMPL = "shift_reg";

assign rnode_348to349_bb4_var__u61_0_reg_349_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u61_stall_in = 1'b0;
assign rnode_348to349_bb4_var__u61_0_NO_SHIFT_REG = rnode_348to349_bb4_var__u61_0_reg_349_NO_SHIFT_REG;
assign rnode_348to349_bb4_var__u61_0_stall_in_reg_349_NO_SHIFT_REG = 1'b0;
assign rnode_348to349_bb4_var__u61_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_348to349_bb4__29_i437_0_valid_out_NO_SHIFT_REG;
 logic rnode_348to349_bb4__29_i437_0_stall_in_NO_SHIFT_REG;
 logic rnode_348to349_bb4__29_i437_0_NO_SHIFT_REG;
 logic rnode_348to349_bb4__29_i437_0_reg_349_inputs_ready_NO_SHIFT_REG;
 logic rnode_348to349_bb4__29_i437_0_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4__29_i437_0_valid_out_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4__29_i437_0_stall_in_reg_349_NO_SHIFT_REG;
 logic rnode_348to349_bb4__29_i437_0_stall_out_reg_349_NO_SHIFT_REG;

acl_data_fifo rnode_348to349_bb4__29_i437_0_reg_349_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_348to349_bb4__29_i437_0_reg_349_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_348to349_bb4__29_i437_0_stall_in_reg_349_NO_SHIFT_REG),
	.valid_out(rnode_348to349_bb4__29_i437_0_valid_out_reg_349_NO_SHIFT_REG),
	.stall_out(rnode_348to349_bb4__29_i437_0_stall_out_reg_349_NO_SHIFT_REG),
	.data_in(local_bb4__29_i437),
	.data_out(rnode_348to349_bb4__29_i437_0_reg_349_NO_SHIFT_REG)
);

defparam rnode_348to349_bb4__29_i437_0_reg_349_fifo.DEPTH = 1;
defparam rnode_348to349_bb4__29_i437_0_reg_349_fifo.DATA_WIDTH = 1;
defparam rnode_348to349_bb4__29_i437_0_reg_349_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_348to349_bb4__29_i437_0_reg_349_fifo.IMPL = "shift_reg";

assign rnode_348to349_bb4__29_i437_0_reg_349_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__29_i437_stall_in = 1'b0;
assign rnode_348to349_bb4__29_i437_0_NO_SHIFT_REG = rnode_348to349_bb4__29_i437_0_reg_349_NO_SHIFT_REG;
assign rnode_348to349_bb4__29_i437_0_stall_in_reg_349_NO_SHIFT_REG = 1'b0;
assign rnode_348to349_bb4__29_i437_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_inc_i452_stall_local;
wire [31:0] local_bb4_inc_i452;

assign local_bb4_inc_i452 = ((rnode_348to350_bb4_add_i449_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp50_not_i457_stall_local;
wire local_bb4_cmp50_not_i457;

assign local_bb4_cmp50_not_i457 = ((rnode_348to350_bb4_add_i449_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_349to351_bb4_reduction_0_i467_0_valid_out_NO_SHIFT_REG;
 logic rnode_349to351_bb4_reduction_0_i467_0_stall_in_NO_SHIFT_REG;
 logic rnode_349to351_bb4_reduction_0_i467_0_NO_SHIFT_REG;
 logic rnode_349to351_bb4_reduction_0_i467_0_reg_351_inputs_ready_NO_SHIFT_REG;
 logic rnode_349to351_bb4_reduction_0_i467_0_reg_351_NO_SHIFT_REG;
 logic rnode_349to351_bb4_reduction_0_i467_0_valid_out_reg_351_NO_SHIFT_REG;
 logic rnode_349to351_bb4_reduction_0_i467_0_stall_in_reg_351_NO_SHIFT_REG;
 logic rnode_349to351_bb4_reduction_0_i467_0_stall_out_reg_351_NO_SHIFT_REG;

acl_data_fifo rnode_349to351_bb4_reduction_0_i467_0_reg_351_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_349to351_bb4_reduction_0_i467_0_reg_351_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_349to351_bb4_reduction_0_i467_0_stall_in_reg_351_NO_SHIFT_REG),
	.valid_out(rnode_349to351_bb4_reduction_0_i467_0_valid_out_reg_351_NO_SHIFT_REG),
	.stall_out(rnode_349to351_bb4_reduction_0_i467_0_stall_out_reg_351_NO_SHIFT_REG),
	.data_in(rnode_348to349_bb4_reduction_0_i467_0_NO_SHIFT_REG),
	.data_out(rnode_349to351_bb4_reduction_0_i467_0_reg_351_NO_SHIFT_REG)
);

defparam rnode_349to351_bb4_reduction_0_i467_0_reg_351_fifo.DEPTH = 2;
defparam rnode_349to351_bb4_reduction_0_i467_0_reg_351_fifo.DATA_WIDTH = 1;
defparam rnode_349to351_bb4_reduction_0_i467_0_reg_351_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_349to351_bb4_reduction_0_i467_0_reg_351_fifo.IMPL = "shift_reg";

assign rnode_349to351_bb4_reduction_0_i467_0_reg_351_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_348to349_bb4_reduction_0_i467_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_349to351_bb4_reduction_0_i467_0_NO_SHIFT_REG = rnode_349to351_bb4_reduction_0_i467_0_reg_351_NO_SHIFT_REG;
assign rnode_349to351_bb4_reduction_0_i467_0_stall_in_reg_351_NO_SHIFT_REG = 1'b0;
assign rnode_349to351_bb4_reduction_0_i467_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_349to350_bb4_var__u61_0_valid_out_NO_SHIFT_REG;
 logic rnode_349to350_bb4_var__u61_0_stall_in_NO_SHIFT_REG;
 logic rnode_349to350_bb4_var__u61_0_NO_SHIFT_REG;
 logic rnode_349to350_bb4_var__u61_0_reg_350_inputs_ready_NO_SHIFT_REG;
 logic rnode_349to350_bb4_var__u61_0_reg_350_NO_SHIFT_REG;
 logic rnode_349to350_bb4_var__u61_0_valid_out_reg_350_NO_SHIFT_REG;
 logic rnode_349to350_bb4_var__u61_0_stall_in_reg_350_NO_SHIFT_REG;
 logic rnode_349to350_bb4_var__u61_0_stall_out_reg_350_NO_SHIFT_REG;

acl_data_fifo rnode_349to350_bb4_var__u61_0_reg_350_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_349to350_bb4_var__u61_0_reg_350_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_349to350_bb4_var__u61_0_stall_in_reg_350_NO_SHIFT_REG),
	.valid_out(rnode_349to350_bb4_var__u61_0_valid_out_reg_350_NO_SHIFT_REG),
	.stall_out(rnode_349to350_bb4_var__u61_0_stall_out_reg_350_NO_SHIFT_REG),
	.data_in(rnode_348to349_bb4_var__u61_0_NO_SHIFT_REG),
	.data_out(rnode_349to350_bb4_var__u61_0_reg_350_NO_SHIFT_REG)
);

defparam rnode_349to350_bb4_var__u61_0_reg_350_fifo.DEPTH = 1;
defparam rnode_349to350_bb4_var__u61_0_reg_350_fifo.DATA_WIDTH = 1;
defparam rnode_349to350_bb4_var__u61_0_reg_350_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_349to350_bb4_var__u61_0_reg_350_fifo.IMPL = "shift_reg";

assign rnode_349to350_bb4_var__u61_0_reg_350_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_348to349_bb4_var__u61_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_349to350_bb4_var__u61_0_NO_SHIFT_REG = rnode_349to350_bb4_var__u61_0_reg_350_NO_SHIFT_REG;
assign rnode_349to350_bb4_var__u61_0_stall_in_reg_350_NO_SHIFT_REG = 1'b0;
assign rnode_349to350_bb4_var__u61_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_349to352_bb4__29_i437_0_valid_out_NO_SHIFT_REG;
 logic rnode_349to352_bb4__29_i437_0_stall_in_NO_SHIFT_REG;
 logic rnode_349to352_bb4__29_i437_0_NO_SHIFT_REG;
 logic rnode_349to352_bb4__29_i437_0_reg_352_inputs_ready_NO_SHIFT_REG;
 logic rnode_349to352_bb4__29_i437_0_reg_352_NO_SHIFT_REG;
 logic rnode_349to352_bb4__29_i437_0_valid_out_reg_352_NO_SHIFT_REG;
 logic rnode_349to352_bb4__29_i437_0_stall_in_reg_352_NO_SHIFT_REG;
 logic rnode_349to352_bb4__29_i437_0_stall_out_reg_352_NO_SHIFT_REG;

acl_data_fifo rnode_349to352_bb4__29_i437_0_reg_352_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_349to352_bb4__29_i437_0_reg_352_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_349to352_bb4__29_i437_0_stall_in_reg_352_NO_SHIFT_REG),
	.valid_out(rnode_349to352_bb4__29_i437_0_valid_out_reg_352_NO_SHIFT_REG),
	.stall_out(rnode_349to352_bb4__29_i437_0_stall_out_reg_352_NO_SHIFT_REG),
	.data_in(rnode_348to349_bb4__29_i437_0_NO_SHIFT_REG),
	.data_out(rnode_349to352_bb4__29_i437_0_reg_352_NO_SHIFT_REG)
);

defparam rnode_349to352_bb4__29_i437_0_reg_352_fifo.DEPTH = 3;
defparam rnode_349to352_bb4__29_i437_0_reg_352_fifo.DATA_WIDTH = 1;
defparam rnode_349to352_bb4__29_i437_0_reg_352_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_349to352_bb4__29_i437_0_reg_352_fifo.IMPL = "shift_reg";

assign rnode_349to352_bb4__29_i437_0_reg_352_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_348to349_bb4__29_i437_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_349to352_bb4__29_i437_0_NO_SHIFT_REG = rnode_349to352_bb4__29_i437_0_reg_352_NO_SHIFT_REG;
assign rnode_349to352_bb4__29_i437_0_stall_in_reg_352_NO_SHIFT_REG = 1'b0;
assign rnode_349to352_bb4__29_i437_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__31_i458_stall_local;
wire local_bb4__31_i458;

assign local_bb4__31_i458 = (local_bb4_tobool49_i451 & local_bb4_cmp50_not_i457);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_351to352_bb4_reduction_0_i467_0_valid_out_NO_SHIFT_REG;
 logic rnode_351to352_bb4_reduction_0_i467_0_stall_in_NO_SHIFT_REG;
 logic rnode_351to352_bb4_reduction_0_i467_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4_reduction_0_i467_0_reg_352_inputs_ready_NO_SHIFT_REG;
 logic rnode_351to352_bb4_reduction_0_i467_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_reduction_0_i467_0_valid_out_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_reduction_0_i467_0_stall_in_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_reduction_0_i467_0_stall_out_reg_352_NO_SHIFT_REG;

acl_data_fifo rnode_351to352_bb4_reduction_0_i467_0_reg_352_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_351to352_bb4_reduction_0_i467_0_reg_352_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_351to352_bb4_reduction_0_i467_0_stall_in_reg_352_NO_SHIFT_REG),
	.valid_out(rnode_351to352_bb4_reduction_0_i467_0_valid_out_reg_352_NO_SHIFT_REG),
	.stall_out(rnode_351to352_bb4_reduction_0_i467_0_stall_out_reg_352_NO_SHIFT_REG),
	.data_in(rnode_349to351_bb4_reduction_0_i467_0_NO_SHIFT_REG),
	.data_out(rnode_351to352_bb4_reduction_0_i467_0_reg_352_NO_SHIFT_REG)
);

defparam rnode_351to352_bb4_reduction_0_i467_0_reg_352_fifo.DEPTH = 1;
defparam rnode_351to352_bb4_reduction_0_i467_0_reg_352_fifo.DATA_WIDTH = 1;
defparam rnode_351to352_bb4_reduction_0_i467_0_reg_352_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_351to352_bb4_reduction_0_i467_0_reg_352_fifo.IMPL = "shift_reg";

assign rnode_351to352_bb4_reduction_0_i467_0_reg_352_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_349to351_bb4_reduction_0_i467_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_reduction_0_i467_0_NO_SHIFT_REG = rnode_351to352_bb4_reduction_0_i467_0_reg_352_NO_SHIFT_REG;
assign rnode_351to352_bb4_reduction_0_i467_0_stall_in_reg_352_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_reduction_0_i467_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_350to351_bb4_var__u61_0_valid_out_NO_SHIFT_REG;
 logic rnode_350to351_bb4_var__u61_0_stall_in_NO_SHIFT_REG;
 logic rnode_350to351_bb4_var__u61_0_NO_SHIFT_REG;
 logic rnode_350to351_bb4_var__u61_0_reg_351_inputs_ready_NO_SHIFT_REG;
 logic rnode_350to351_bb4_var__u61_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_var__u61_0_valid_out_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_var__u61_0_stall_in_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_var__u61_0_stall_out_reg_351_NO_SHIFT_REG;

acl_data_fifo rnode_350to351_bb4_var__u61_0_reg_351_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_350to351_bb4_var__u61_0_reg_351_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_350to351_bb4_var__u61_0_stall_in_reg_351_NO_SHIFT_REG),
	.valid_out(rnode_350to351_bb4_var__u61_0_valid_out_reg_351_NO_SHIFT_REG),
	.stall_out(rnode_350to351_bb4_var__u61_0_stall_out_reg_351_NO_SHIFT_REG),
	.data_in(rnode_349to350_bb4_var__u61_0_NO_SHIFT_REG),
	.data_out(rnode_350to351_bb4_var__u61_0_reg_351_NO_SHIFT_REG)
);

defparam rnode_350to351_bb4_var__u61_0_reg_351_fifo.DEPTH = 1;
defparam rnode_350to351_bb4_var__u61_0_reg_351_fifo.DATA_WIDTH = 1;
defparam rnode_350to351_bb4_var__u61_0_reg_351_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_350to351_bb4_var__u61_0_reg_351_fifo.IMPL = "shift_reg";

assign rnode_350to351_bb4_var__u61_0_reg_351_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_349to350_bb4_var__u61_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4_var__u61_0_NO_SHIFT_REG = rnode_350to351_bb4_var__u61_0_reg_351_NO_SHIFT_REG;
assign rnode_350to351_bb4_var__u61_0_stall_in_reg_351_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4_var__u61_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_352to353_bb4__29_i437_0_valid_out_NO_SHIFT_REG;
 logic rnode_352to353_bb4__29_i437_0_stall_in_NO_SHIFT_REG;
 logic rnode_352to353_bb4__29_i437_0_NO_SHIFT_REG;
 logic rnode_352to353_bb4__29_i437_0_reg_353_inputs_ready_NO_SHIFT_REG;
 logic rnode_352to353_bb4__29_i437_0_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4__29_i437_0_valid_out_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4__29_i437_0_stall_in_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4__29_i437_0_stall_out_reg_353_NO_SHIFT_REG;

acl_data_fifo rnode_352to353_bb4__29_i437_0_reg_353_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_352to353_bb4__29_i437_0_reg_353_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_352to353_bb4__29_i437_0_stall_in_reg_353_NO_SHIFT_REG),
	.valid_out(rnode_352to353_bb4__29_i437_0_valid_out_reg_353_NO_SHIFT_REG),
	.stall_out(rnode_352to353_bb4__29_i437_0_stall_out_reg_353_NO_SHIFT_REG),
	.data_in(rnode_349to352_bb4__29_i437_0_NO_SHIFT_REG),
	.data_out(rnode_352to353_bb4__29_i437_0_reg_353_NO_SHIFT_REG)
);

defparam rnode_352to353_bb4__29_i437_0_reg_353_fifo.DEPTH = 1;
defparam rnode_352to353_bb4__29_i437_0_reg_353_fifo.DATA_WIDTH = 1;
defparam rnode_352to353_bb4__29_i437_0_reg_353_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_352to353_bb4__29_i437_0_reg_353_fifo.IMPL = "shift_reg";

assign rnode_352to353_bb4__29_i437_0_reg_353_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_349to352_bb4__29_i437_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_352to353_bb4__29_i437_0_NO_SHIFT_REG = rnode_352to353_bb4__29_i437_0_reg_353_NO_SHIFT_REG;
assign rnode_352to353_bb4__29_i437_0_stall_in_reg_353_NO_SHIFT_REG = 1'b0;
assign rnode_352to353_bb4__29_i437_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__32_i459_stall_local;
wire [31:0] local_bb4__32_i459;

assign local_bb4__32_i459 = (local_bb4__31_i458 ? (local_bb4_shl1_i_i456 & 32'hFFFFFE00) : (local_bb4_shl1_i18_i448 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__34_i461_stall_local;
wire [31:0] local_bb4__34_i461;

assign local_bb4__34_i461 = (local_bb4__31_i458 ? (local_bb4_or_i_i455 & 32'h1FFFFFF) : (local_bb4_or_i17_i447 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__36_i463_stall_local;
wire [31:0] local_bb4__36_i463;

assign local_bb4__36_i463 = (local_bb4__31_i458 ? (rnode_348to350_bb4_add_i449_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i460_stall_local;
wire [31:0] local_bb4__33_i460;

assign local_bb4__33_i460 = (local_bb4_tobool49_i451 ? (local_bb4__32_i459 & 32'hFFFFFF00) : (local_bb4_shl1_i18_i448 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__35_i462_stall_local;
wire [31:0] local_bb4__35_i462;

assign local_bb4__35_i462 = (local_bb4_tobool49_i451 ? (local_bb4__34_i461 & 32'h1FFFFFF) : (local_bb4_or_i17_i447 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__37_i464_stall_local;
wire [31:0] local_bb4__37_i464;

assign local_bb4__37_i464 = (local_bb4_tobool49_i451 ? (local_bb4__36_i463 & 32'h1FF) : (local_bb4_inc_i452 & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i470_stall_local;
wire [31:0] local_bb4_and75_i470;

assign local_bb4_and75_i470 = ((local_bb4__35_i462 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i460_valid_out;
wire local_bb4__33_i460_stall_in;
wire local_bb4__37_i464_valid_out;
wire local_bb4__37_i464_stall_in;
wire local_bb4_and75_i470_valid_out;
wire local_bb4_and75_i470_stall_in;
wire local_bb4_and83_i476_valid_out;
wire local_bb4_and83_i476_stall_in;
wire local_bb4_and83_i476_inputs_ready;
wire local_bb4_and83_i476_stall_local;
wire [31:0] local_bb4_and83_i476;

assign local_bb4_and83_i476_inputs_ready = (local_bb4_mul_i_i442_valid_out_0_NO_SHIFT_REG & rnode_348to350_bb4_add_i449_0_valid_out_1_NO_SHIFT_REG & rnode_348to350_bb4_add_i449_0_valid_out_0_NO_SHIFT_REG & rnode_348to350_bb4_add_i449_0_valid_out_2_NO_SHIFT_REG & local_bb4_mul_i_i442_valid_out_1_NO_SHIFT_REG);
assign local_bb4_and83_i476 = ((local_bb4__35_i462 & 32'h1FFFFFF) & 32'h1);
assign local_bb4__33_i460_valid_out = 1'b1;
assign local_bb4__37_i464_valid_out = 1'b1;
assign local_bb4_and75_i470_valid_out = 1'b1;
assign local_bb4_and83_i476_valid_out = 1'b1;
assign local_bb4_mul_i_i442_stall_in_0 = 1'b0;
assign rnode_348to350_bb4_add_i449_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_348to350_bb4_add_i449_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_348to350_bb4_add_i449_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign local_bb4_mul_i_i442_stall_in_1 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_350to351_bb4__33_i460_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_350to351_bb4__33_i460_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__33_i460_0_NO_SHIFT_REG;
 logic rnode_350to351_bb4__33_i460_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_350to351_bb4__33_i460_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__33_i460_1_NO_SHIFT_REG;
 logic rnode_350to351_bb4__33_i460_0_reg_351_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__33_i460_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4__33_i460_0_valid_out_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4__33_i460_0_stall_in_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4__33_i460_0_stall_out_reg_351_NO_SHIFT_REG;

acl_data_fifo rnode_350to351_bb4__33_i460_0_reg_351_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_350to351_bb4__33_i460_0_reg_351_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_350to351_bb4__33_i460_0_stall_in_0_reg_351_NO_SHIFT_REG),
	.valid_out(rnode_350to351_bb4__33_i460_0_valid_out_0_reg_351_NO_SHIFT_REG),
	.stall_out(rnode_350to351_bb4__33_i460_0_stall_out_reg_351_NO_SHIFT_REG),
	.data_in((local_bb4__33_i460 & 32'hFFFFFF00)),
	.data_out(rnode_350to351_bb4__33_i460_0_reg_351_NO_SHIFT_REG)
);

defparam rnode_350to351_bb4__33_i460_0_reg_351_fifo.DEPTH = 1;
defparam rnode_350to351_bb4__33_i460_0_reg_351_fifo.DATA_WIDTH = 32;
defparam rnode_350to351_bb4__33_i460_0_reg_351_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_350to351_bb4__33_i460_0_reg_351_fifo.IMPL = "shift_reg";

assign rnode_350to351_bb4__33_i460_0_reg_351_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__33_i460_stall_in = 1'b0;
assign rnode_350to351_bb4__33_i460_0_stall_in_0_reg_351_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4__33_i460_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_350to351_bb4__33_i460_0_NO_SHIFT_REG = rnode_350to351_bb4__33_i460_0_reg_351_NO_SHIFT_REG;
assign rnode_350to351_bb4__33_i460_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_350to351_bb4__33_i460_1_NO_SHIFT_REG = rnode_350to351_bb4__33_i460_0_reg_351_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_350to351_bb4__37_i464_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__37_i464_0_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__37_i464_1_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__37_i464_2_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__37_i464_3_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_reg_351_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4__37_i464_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_valid_out_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_stall_in_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4__37_i464_0_stall_out_reg_351_NO_SHIFT_REG;

acl_data_fifo rnode_350to351_bb4__37_i464_0_reg_351_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_350to351_bb4__37_i464_0_reg_351_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_350to351_bb4__37_i464_0_stall_in_0_reg_351_NO_SHIFT_REG),
	.valid_out(rnode_350to351_bb4__37_i464_0_valid_out_0_reg_351_NO_SHIFT_REG),
	.stall_out(rnode_350to351_bb4__37_i464_0_stall_out_reg_351_NO_SHIFT_REG),
	.data_in((local_bb4__37_i464 & 32'h3FF)),
	.data_out(rnode_350to351_bb4__37_i464_0_reg_351_NO_SHIFT_REG)
);

defparam rnode_350to351_bb4__37_i464_0_reg_351_fifo.DEPTH = 1;
defparam rnode_350to351_bb4__37_i464_0_reg_351_fifo.DATA_WIDTH = 32;
defparam rnode_350to351_bb4__37_i464_0_reg_351_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_350to351_bb4__37_i464_0_reg_351_fifo.IMPL = "shift_reg";

assign rnode_350to351_bb4__37_i464_0_reg_351_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__37_i464_stall_in = 1'b0;
assign rnode_350to351_bb4__37_i464_0_stall_in_0_reg_351_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4__37_i464_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_350to351_bb4__37_i464_0_NO_SHIFT_REG = rnode_350to351_bb4__37_i464_0_reg_351_NO_SHIFT_REG;
assign rnode_350to351_bb4__37_i464_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_350to351_bb4__37_i464_1_NO_SHIFT_REG = rnode_350to351_bb4__37_i464_0_reg_351_NO_SHIFT_REG;
assign rnode_350to351_bb4__37_i464_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_350to351_bb4__37_i464_2_NO_SHIFT_REG = rnode_350to351_bb4__37_i464_0_reg_351_NO_SHIFT_REG;
assign rnode_350to351_bb4__37_i464_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_350to351_bb4__37_i464_3_NO_SHIFT_REG = rnode_350to351_bb4__37_i464_0_reg_351_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_350to351_bb4_and75_i470_0_valid_out_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and75_i470_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4_and75_i470_0_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and75_i470_0_reg_351_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4_and75_i470_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and75_i470_0_valid_out_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and75_i470_0_stall_in_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and75_i470_0_stall_out_reg_351_NO_SHIFT_REG;

acl_data_fifo rnode_350to351_bb4_and75_i470_0_reg_351_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_350to351_bb4_and75_i470_0_reg_351_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_350to351_bb4_and75_i470_0_stall_in_reg_351_NO_SHIFT_REG),
	.valid_out(rnode_350to351_bb4_and75_i470_0_valid_out_reg_351_NO_SHIFT_REG),
	.stall_out(rnode_350to351_bb4_and75_i470_0_stall_out_reg_351_NO_SHIFT_REG),
	.data_in((local_bb4_and75_i470 & 32'h7FFFFF)),
	.data_out(rnode_350to351_bb4_and75_i470_0_reg_351_NO_SHIFT_REG)
);

defparam rnode_350to351_bb4_and75_i470_0_reg_351_fifo.DEPTH = 1;
defparam rnode_350to351_bb4_and75_i470_0_reg_351_fifo.DATA_WIDTH = 32;
defparam rnode_350to351_bb4_and75_i470_0_reg_351_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_350to351_bb4_and75_i470_0_reg_351_fifo.IMPL = "shift_reg";

assign rnode_350to351_bb4_and75_i470_0_reg_351_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and75_i470_stall_in = 1'b0;
assign rnode_350to351_bb4_and75_i470_0_NO_SHIFT_REG = rnode_350to351_bb4_and75_i470_0_reg_351_NO_SHIFT_REG;
assign rnode_350to351_bb4_and75_i470_0_stall_in_reg_351_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4_and75_i470_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_350to351_bb4_and83_i476_0_valid_out_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and83_i476_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4_and83_i476_0_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and83_i476_0_reg_351_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_350to351_bb4_and83_i476_0_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and83_i476_0_valid_out_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and83_i476_0_stall_in_reg_351_NO_SHIFT_REG;
 logic rnode_350to351_bb4_and83_i476_0_stall_out_reg_351_NO_SHIFT_REG;

acl_data_fifo rnode_350to351_bb4_and83_i476_0_reg_351_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_350to351_bb4_and83_i476_0_reg_351_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_350to351_bb4_and83_i476_0_stall_in_reg_351_NO_SHIFT_REG),
	.valid_out(rnode_350to351_bb4_and83_i476_0_valid_out_reg_351_NO_SHIFT_REG),
	.stall_out(rnode_350to351_bb4_and83_i476_0_stall_out_reg_351_NO_SHIFT_REG),
	.data_in((local_bb4_and83_i476 & 32'h1)),
	.data_out(rnode_350to351_bb4_and83_i476_0_reg_351_NO_SHIFT_REG)
);

defparam rnode_350to351_bb4_and83_i476_0_reg_351_fifo.DEPTH = 1;
defparam rnode_350to351_bb4_and83_i476_0_reg_351_fifo.DATA_WIDTH = 32;
defparam rnode_350to351_bb4_and83_i476_0_reg_351_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_350to351_bb4_and83_i476_0_reg_351_fifo.IMPL = "shift_reg";

assign rnode_350to351_bb4_and83_i476_0_reg_351_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and83_i476_stall_in = 1'b0;
assign rnode_350to351_bb4_and83_i476_0_NO_SHIFT_REG = rnode_350to351_bb4_and83_i476_0_reg_351_NO_SHIFT_REG;
assign rnode_350to351_bb4_and83_i476_0_stall_in_reg_351_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4_and83_i476_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i475_stall_local;
wire local_bb4_cmp77_i475;

assign local_bb4_cmp77_i475 = ((rnode_350to351_bb4__33_i460_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u63_stall_local;
wire local_bb4_var__u63;

assign local_bb4_var__u63 = ($signed((rnode_350to351_bb4__33_i460_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp53_i465_stall_local;
wire local_bb4_cmp53_i465;

assign local_bb4_cmp53_i465 = ((rnode_350to351_bb4__37_i464_0_NO_SHIFT_REG & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp68_i469_valid_out;
wire local_bb4_cmp68_i469_stall_in;
wire local_bb4_cmp68_i469_inputs_ready;
wire local_bb4_cmp68_i469_stall_local;
wire local_bb4_cmp68_i469;

assign local_bb4_cmp68_i469_inputs_ready = rnode_350to351_bb4__37_i464_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp68_i469 = ((rnode_350to351_bb4__37_i464_1_NO_SHIFT_REG & 32'h3FF) < 32'h80);
assign local_bb4_cmp68_i469_valid_out = 1'b1;
assign rnode_350to351_bb4__37_i464_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i471_stall_local;
wire [31:0] local_bb4_sub_i471;

assign local_bb4_sub_i471 = ((rnode_350to351_bb4__37_i464_2_NO_SHIFT_REG & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp71_not_i486_valid_out;
wire local_bb4_cmp71_not_i486_stall_in;
wire local_bb4_cmp71_not_i486_inputs_ready;
wire local_bb4_cmp71_not_i486_stall_local;
wire local_bb4_cmp71_not_i486;

assign local_bb4_cmp71_not_i486_inputs_ready = rnode_350to351_bb4__37_i464_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4_cmp71_not_i486 = ((rnode_350to351_bb4__37_i464_3_NO_SHIFT_REG & 32'h3FF) != 32'h7F);
assign local_bb4_cmp71_not_i486_valid_out = 1'b1;
assign rnode_350to351_bb4__37_i464_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool84_i477_stall_local;
wire local_bb4_tobool84_i477;

assign local_bb4_tobool84_i477 = ((rnode_350to351_bb4_and83_i476_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or581_i466_valid_out;
wire local_bb4_or581_i466_stall_in;
wire local_bb4_or581_i466_inputs_ready;
wire local_bb4_or581_i466_stall_local;
wire local_bb4_or581_i466;

assign local_bb4_or581_i466_inputs_ready = (rnode_350to351_bb4_var__u61_0_valid_out_NO_SHIFT_REG & rnode_350to351_bb4__37_i464_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_or581_i466 = (rnode_350to351_bb4_var__u61_0_NO_SHIFT_REG | local_bb4_cmp53_i465);
assign local_bb4_or581_i466_valid_out = 1'b1;
assign rnode_350to351_bb4_var__u61_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4__37_i464_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_351to352_bb4_cmp68_i469_0_valid_out_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp68_i469_0_stall_in_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp68_i469_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp68_i469_0_reg_352_inputs_ready_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp68_i469_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp68_i469_0_valid_out_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp68_i469_0_stall_in_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp68_i469_0_stall_out_reg_352_NO_SHIFT_REG;

acl_data_fifo rnode_351to352_bb4_cmp68_i469_0_reg_352_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_351to352_bb4_cmp68_i469_0_reg_352_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_351to352_bb4_cmp68_i469_0_stall_in_reg_352_NO_SHIFT_REG),
	.valid_out(rnode_351to352_bb4_cmp68_i469_0_valid_out_reg_352_NO_SHIFT_REG),
	.stall_out(rnode_351to352_bb4_cmp68_i469_0_stall_out_reg_352_NO_SHIFT_REG),
	.data_in(local_bb4_cmp68_i469),
	.data_out(rnode_351to352_bb4_cmp68_i469_0_reg_352_NO_SHIFT_REG)
);

defparam rnode_351to352_bb4_cmp68_i469_0_reg_352_fifo.DEPTH = 1;
defparam rnode_351to352_bb4_cmp68_i469_0_reg_352_fifo.DATA_WIDTH = 1;
defparam rnode_351to352_bb4_cmp68_i469_0_reg_352_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_351to352_bb4_cmp68_i469_0_reg_352_fifo.IMPL = "shift_reg";

assign rnode_351to352_bb4_cmp68_i469_0_reg_352_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp68_i469_stall_in = 1'b0;
assign rnode_351to352_bb4_cmp68_i469_0_NO_SHIFT_REG = rnode_351to352_bb4_cmp68_i469_0_reg_352_NO_SHIFT_REG;
assign rnode_351to352_bb4_cmp68_i469_0_stall_in_reg_352_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_cmp68_i469_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and74_i472_stall_local;
wire [31:0] local_bb4_and74_i472;

assign local_bb4_and74_i472 = ((local_bb4_sub_i471 & 32'hFF800000) + 32'h40800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_351to352_bb4_cmp71_not_i486_0_valid_out_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp71_not_i486_0_stall_in_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp71_not_i486_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp71_not_i486_0_reg_352_inputs_ready_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp71_not_i486_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp71_not_i486_0_valid_out_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp71_not_i486_0_stall_in_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_cmp71_not_i486_0_stall_out_reg_352_NO_SHIFT_REG;

acl_data_fifo rnode_351to352_bb4_cmp71_not_i486_0_reg_352_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_351to352_bb4_cmp71_not_i486_0_reg_352_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_351to352_bb4_cmp71_not_i486_0_stall_in_reg_352_NO_SHIFT_REG),
	.valid_out(rnode_351to352_bb4_cmp71_not_i486_0_valid_out_reg_352_NO_SHIFT_REG),
	.stall_out(rnode_351to352_bb4_cmp71_not_i486_0_stall_out_reg_352_NO_SHIFT_REG),
	.data_in(local_bb4_cmp71_not_i486),
	.data_out(rnode_351to352_bb4_cmp71_not_i486_0_reg_352_NO_SHIFT_REG)
);

defparam rnode_351to352_bb4_cmp71_not_i486_0_reg_352_fifo.DEPTH = 1;
defparam rnode_351to352_bb4_cmp71_not_i486_0_reg_352_fifo.DATA_WIDTH = 1;
defparam rnode_351to352_bb4_cmp71_not_i486_0_reg_352_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_351to352_bb4_cmp71_not_i486_0_reg_352_fifo.IMPL = "shift_reg";

assign rnode_351to352_bb4_cmp71_not_i486_0_reg_352_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp71_not_i486_stall_in = 1'b0;
assign rnode_351to352_bb4_cmp71_not_i486_0_NO_SHIFT_REG = rnode_351to352_bb4_cmp71_not_i486_0_reg_352_NO_SHIFT_REG;
assign rnode_351to352_bb4_cmp71_not_i486_0_stall_in_reg_352_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_cmp71_not_i486_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__39_i478_stall_local;
wire local_bb4__39_i478;

assign local_bb4__39_i478 = (local_bb4_tobool84_i477 & local_bb4_var__u63);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_351to352_bb4_or581_i466_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_1_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_reg_352_inputs_ready_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_valid_out_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_stall_in_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or581_i466_0_stall_out_reg_352_NO_SHIFT_REG;

acl_data_fifo rnode_351to352_bb4_or581_i466_0_reg_352_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_351to352_bb4_or581_i466_0_reg_352_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_351to352_bb4_or581_i466_0_stall_in_0_reg_352_NO_SHIFT_REG),
	.valid_out(rnode_351to352_bb4_or581_i466_0_valid_out_0_reg_352_NO_SHIFT_REG),
	.stall_out(rnode_351to352_bb4_or581_i466_0_stall_out_reg_352_NO_SHIFT_REG),
	.data_in(local_bb4_or581_i466),
	.data_out(rnode_351to352_bb4_or581_i466_0_reg_352_NO_SHIFT_REG)
);

defparam rnode_351to352_bb4_or581_i466_0_reg_352_fifo.DEPTH = 1;
defparam rnode_351to352_bb4_or581_i466_0_reg_352_fifo.DATA_WIDTH = 1;
defparam rnode_351to352_bb4_or581_i466_0_reg_352_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_351to352_bb4_or581_i466_0_reg_352_fifo.IMPL = "shift_reg";

assign rnode_351to352_bb4_or581_i466_0_reg_352_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or581_i466_stall_in = 1'b0;
assign rnode_351to352_bb4_or581_i466_0_stall_in_0_reg_352_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_or581_i466_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_351to352_bb4_or581_i466_0_NO_SHIFT_REG = rnode_351to352_bb4_or581_i466_0_reg_352_NO_SHIFT_REG;
assign rnode_351to352_bb4_or581_i466_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_351to352_bb4_or581_i466_1_NO_SHIFT_REG = rnode_351to352_bb4_or581_i466_0_reg_352_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u64_stall_local;
wire [31:0] local_bb4_var__u64;

assign local_bb4_var__u64[31:1] = 31'h0;
assign local_bb4_var__u64[0] = rnode_351to352_bb4_cmp68_i469_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i473_stall_local;
wire [31:0] local_bb4_shl_i473;

assign local_bb4_shl_i473 = ((local_bb4_and74_i472 & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4__40_i479_valid_out;
wire local_bb4__40_i479_stall_in;
wire local_bb4__40_i479_inputs_ready;
wire local_bb4__40_i479_stall_local;
wire local_bb4__40_i479;

assign local_bb4__40_i479_inputs_ready = (rnode_350to351_bb4__33_i460_0_valid_out_0_NO_SHIFT_REG & rnode_350to351_bb4__33_i460_0_valid_out_1_NO_SHIFT_REG & rnode_350to351_bb4_and83_i476_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40_i479 = (local_bb4_cmp77_i475 | local_bb4__39_i478);
assign local_bb4__40_i479_valid_out = 1'b1;
assign rnode_350to351_bb4__33_i460_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4__33_i460_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4_and83_i476_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i468_stall_local;
wire local_bb4_reduction_2_i468;

assign local_bb4_reduction_2_i468 = (rnode_351to352_bb4_reduction_0_i467_0_NO_SHIFT_REG | rnode_351to352_bb4_or581_i466_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_352to353_bb4_or581_i466_0_valid_out_NO_SHIFT_REG;
 logic rnode_352to353_bb4_or581_i466_0_stall_in_NO_SHIFT_REG;
 logic rnode_352to353_bb4_or581_i466_0_NO_SHIFT_REG;
 logic rnode_352to353_bb4_or581_i466_0_reg_353_inputs_ready_NO_SHIFT_REG;
 logic rnode_352to353_bb4_or581_i466_0_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4_or581_i466_0_valid_out_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4_or581_i466_0_stall_in_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4_or581_i466_0_stall_out_reg_353_NO_SHIFT_REG;

acl_data_fifo rnode_352to353_bb4_or581_i466_0_reg_353_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_352to353_bb4_or581_i466_0_reg_353_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_352to353_bb4_or581_i466_0_stall_in_reg_353_NO_SHIFT_REG),
	.valid_out(rnode_352to353_bb4_or581_i466_0_valid_out_reg_353_NO_SHIFT_REG),
	.stall_out(rnode_352to353_bb4_or581_i466_0_stall_out_reg_353_NO_SHIFT_REG),
	.data_in(rnode_351to352_bb4_or581_i466_1_NO_SHIFT_REG),
	.data_out(rnode_352to353_bb4_or581_i466_0_reg_353_NO_SHIFT_REG)
);

defparam rnode_352to353_bb4_or581_i466_0_reg_353_fifo.DEPTH = 1;
defparam rnode_352to353_bb4_or581_i466_0_reg_353_fifo.DATA_WIDTH = 1;
defparam rnode_352to353_bb4_or581_i466_0_reg_353_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_352to353_bb4_or581_i466_0_reg_353_fifo.IMPL = "shift_reg";

assign rnode_352to353_bb4_or581_i466_0_reg_353_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_351to352_bb4_or581_i466_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_352to353_bb4_or581_i466_0_NO_SHIFT_REG = rnode_352to353_bb4_or581_i466_0_reg_353_NO_SHIFT_REG;
assign rnode_352to353_bb4_or581_i466_0_stall_in_reg_353_NO_SHIFT_REG = 1'b0;
assign rnode_352to353_bb4_or581_i466_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or76_i474_valid_out;
wire local_bb4_or76_i474_stall_in;
wire local_bb4_or76_i474_inputs_ready;
wire local_bb4_or76_i474_stall_local;
wire [31:0] local_bb4_or76_i474;

assign local_bb4_or76_i474_inputs_ready = (rnode_350to351_bb4__37_i464_0_valid_out_2_NO_SHIFT_REG & rnode_350to351_bb4_and75_i470_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or76_i474 = ((local_bb4_shl_i473 & 32'h7F800000) | (rnode_350to351_bb4_and75_i470_0_NO_SHIFT_REG & 32'h7FFFFF));
assign local_bb4_or76_i474_valid_out = 1'b1;
assign rnode_350to351_bb4__37_i464_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_350to351_bb4_and75_i470_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_351to352_bb4__40_i479_0_valid_out_NO_SHIFT_REG;
 logic rnode_351to352_bb4__40_i479_0_stall_in_NO_SHIFT_REG;
 logic rnode_351to352_bb4__40_i479_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4__40_i479_0_reg_352_inputs_ready_NO_SHIFT_REG;
 logic rnode_351to352_bb4__40_i479_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4__40_i479_0_valid_out_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4__40_i479_0_stall_in_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4__40_i479_0_stall_out_reg_352_NO_SHIFT_REG;

acl_data_fifo rnode_351to352_bb4__40_i479_0_reg_352_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_351to352_bb4__40_i479_0_reg_352_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_351to352_bb4__40_i479_0_stall_in_reg_352_NO_SHIFT_REG),
	.valid_out(rnode_351to352_bb4__40_i479_0_valid_out_reg_352_NO_SHIFT_REG),
	.stall_out(rnode_351to352_bb4__40_i479_0_stall_out_reg_352_NO_SHIFT_REG),
	.data_in(local_bb4__40_i479),
	.data_out(rnode_351to352_bb4__40_i479_0_reg_352_NO_SHIFT_REG)
);

defparam rnode_351to352_bb4__40_i479_0_reg_352_fifo.DEPTH = 1;
defparam rnode_351to352_bb4__40_i479_0_reg_352_fifo.DATA_WIDTH = 1;
defparam rnode_351to352_bb4__40_i479_0_reg_352_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_351to352_bb4__40_i479_0_reg_352_fifo.IMPL = "shift_reg";

assign rnode_351to352_bb4__40_i479_0_reg_352_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_i479_stall_in = 1'b0;
assign rnode_351to352_bb4__40_i479_0_NO_SHIFT_REG = rnode_351to352_bb4__40_i479_0_reg_352_NO_SHIFT_REG;
assign rnode_351to352_bb4__40_i479_0_stall_in_reg_352_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4__40_i479_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_conv101_i489_stall_local;
wire [31:0] local_bb4_conv101_i489;

assign local_bb4_conv101_i489[31:1] = 31'h0;
assign local_bb4_conv101_i489[0] = local_bb4_reduction_2_i468;

// This section implements an unregistered operation.
// 
wire local_bb4_cond111_i494_stall_local;
wire [31:0] local_bb4_cond111_i494;

assign local_bb4_cond111_i494 = (rnode_352to353_bb4_or581_i466_0_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_351to352_bb4_or76_i474_0_valid_out_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or76_i474_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_351to352_bb4_or76_i474_0_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or76_i474_0_reg_352_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_351to352_bb4_or76_i474_0_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or76_i474_0_valid_out_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or76_i474_0_stall_in_reg_352_NO_SHIFT_REG;
 logic rnode_351to352_bb4_or76_i474_0_stall_out_reg_352_NO_SHIFT_REG;

acl_data_fifo rnode_351to352_bb4_or76_i474_0_reg_352_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_351to352_bb4_or76_i474_0_reg_352_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_351to352_bb4_or76_i474_0_stall_in_reg_352_NO_SHIFT_REG),
	.valid_out(rnode_351to352_bb4_or76_i474_0_valid_out_reg_352_NO_SHIFT_REG),
	.stall_out(rnode_351to352_bb4_or76_i474_0_stall_out_reg_352_NO_SHIFT_REG),
	.data_in((local_bb4_or76_i474 & 32'h7FFFFFFF)),
	.data_out(rnode_351to352_bb4_or76_i474_0_reg_352_NO_SHIFT_REG)
);

defparam rnode_351to352_bb4_or76_i474_0_reg_352_fifo.DEPTH = 1;
defparam rnode_351to352_bb4_or76_i474_0_reg_352_fifo.DATA_WIDTH = 32;
defparam rnode_351to352_bb4_or76_i474_0_reg_352_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_351to352_bb4_or76_i474_0_reg_352_fifo.IMPL = "shift_reg";

assign rnode_351to352_bb4_or76_i474_0_reg_352_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or76_i474_stall_in = 1'b0;
assign rnode_351to352_bb4_or76_i474_0_NO_SHIFT_REG = rnode_351to352_bb4_or76_i474_0_reg_352_NO_SHIFT_REG;
assign rnode_351to352_bb4_or76_i474_0_stall_in_reg_352_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_or76_i474_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cond_i480_stall_local;
wire [31:0] local_bb4_cond_i480;

assign local_bb4_cond_i480[31:1] = 31'h0;
assign local_bb4_cond_i480[0] = rnode_351to352_bb4__40_i479_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add87_i481_stall_local;
wire [31:0] local_bb4_add87_i481;

assign local_bb4_add87_i481 = ((local_bb4_cond_i480 & 32'h1) + (rnode_351to352_bb4_or76_i474_0_NO_SHIFT_REG & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i484_stall_local;
wire [31:0] local_bb4_and90_i484;

assign local_bb4_and90_i484 = (local_bb4_add87_i481 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i485_stall_local;
wire local_bb4_cmp91_i485;

assign local_bb4_cmp91_i485 = ((local_bb4_and90_i484 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge14_i487_stall_local;
wire local_bb4_brmerge14_i487;

assign local_bb4_brmerge14_i487 = (local_bb4_cmp91_i485 | rnode_351to352_bb4_cmp71_not_i486_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_conv99_i488_stall_local;
wire [31:0] local_bb4_conv99_i488;

assign local_bb4_conv99_i488 = (local_bb4_brmerge14_i487 ? (local_bb4_var__u64 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or102_i490_stall_local;
wire [31:0] local_bb4_or102_i490;

assign local_bb4_or102_i490 = ((local_bb4_conv99_i488 & 32'h1) | (local_bb4_conv101_i489 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_sext_stall_local;
wire [31:0] local_bb4_sext;

assign local_bb4_sext = ((local_bb4_or102_i490 & 32'h1) + 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and108_i493_valid_out;
wire local_bb4_and108_i493_stall_in;
wire local_bb4_and108_i493_inputs_ready;
wire local_bb4_and108_i493_stall_local;
wire [31:0] local_bb4_and108_i493;

assign local_bb4_and108_i493_inputs_ready = (rnode_351to352_bb4_or581_i466_0_valid_out_0_NO_SHIFT_REG & rnode_351to352_bb4_reduction_0_i467_0_valid_out_NO_SHIFT_REG & rnode_351to352_bb4_cmp68_i469_0_valid_out_NO_SHIFT_REG & rnode_351to352_bb4_cmp71_not_i486_0_valid_out_NO_SHIFT_REG & rnode_351to352_bb4__40_i479_0_valid_out_NO_SHIFT_REG & rnode_351to352_bb4_or76_i474_0_valid_out_NO_SHIFT_REG);
assign local_bb4_and108_i493 = (local_bb4_sext & local_bb4_add87_i481);
assign local_bb4_and108_i493_valid_out = 1'b1;
assign rnode_351to352_bb4_or581_i466_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_reduction_0_i467_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_cmp68_i469_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_cmp71_not_i486_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4__40_i479_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_351to352_bb4_or76_i474_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_352to353_bb4_and108_i493_0_valid_out_NO_SHIFT_REG;
 logic rnode_352to353_bb4_and108_i493_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_352to353_bb4_and108_i493_0_NO_SHIFT_REG;
 logic rnode_352to353_bb4_and108_i493_0_reg_353_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_352to353_bb4_and108_i493_0_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4_and108_i493_0_valid_out_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4_and108_i493_0_stall_in_reg_353_NO_SHIFT_REG;
 logic rnode_352to353_bb4_and108_i493_0_stall_out_reg_353_NO_SHIFT_REG;

acl_data_fifo rnode_352to353_bb4_and108_i493_0_reg_353_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_352to353_bb4_and108_i493_0_reg_353_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_352to353_bb4_and108_i493_0_stall_in_reg_353_NO_SHIFT_REG),
	.valid_out(rnode_352to353_bb4_and108_i493_0_valid_out_reg_353_NO_SHIFT_REG),
	.stall_out(rnode_352to353_bb4_and108_i493_0_stall_out_reg_353_NO_SHIFT_REG),
	.data_in(local_bb4_and108_i493),
	.data_out(rnode_352to353_bb4_and108_i493_0_reg_353_NO_SHIFT_REG)
);

defparam rnode_352to353_bb4_and108_i493_0_reg_353_fifo.DEPTH = 1;
defparam rnode_352to353_bb4_and108_i493_0_reg_353_fifo.DATA_WIDTH = 32;
defparam rnode_352to353_bb4_and108_i493_0_reg_353_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_352to353_bb4_and108_i493_0_reg_353_fifo.IMPL = "shift_reg";

assign rnode_352to353_bb4_and108_i493_0_reg_353_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and108_i493_stall_in = 1'b0;
assign rnode_352to353_bb4_and108_i493_0_NO_SHIFT_REG = rnode_352to353_bb4_and108_i493_0_reg_353_NO_SHIFT_REG;
assign rnode_352to353_bb4_and108_i493_0_stall_in_reg_353_NO_SHIFT_REG = 1'b0;
assign rnode_352to353_bb4_and108_i493_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or112_i495_stall_local;
wire [31:0] local_bb4_or112_i495;

assign local_bb4_or112_i495 = (rnode_352to353_bb4_and108_i493_0_NO_SHIFT_REG | (local_bb4_cond111_i494 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_or112_i495_op_stall_local;
wire [31:0] local_bb4_or112_i495_op;

assign local_bb4_or112_i495_op = (local_bb4_or112_i495 | 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u65_stall_local;
wire [31:0] local_bb4_var__u65;

assign local_bb4_var__u65 = (local_bb4_or112_i495_op | 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_cast_after_negation_valid_out;
wire local_bb4_cast_after_negation_stall_in;
wire local_bb4_cast_after_negation_inputs_ready;
wire local_bb4_cast_after_negation_stall_local;
wire [31:0] local_bb4_cast_after_negation;

assign local_bb4_cast_after_negation_inputs_ready = (rnode_352to353_bb4__29_i437_0_valid_out_NO_SHIFT_REG & rnode_352to353_bb4_or581_i466_0_valid_out_NO_SHIFT_REG & rnode_352to353_bb4_and108_i493_0_valid_out_NO_SHIFT_REG);
assign local_bb4_cast_after_negation = (rnode_352to353_bb4__29_i437_0_NO_SHIFT_REG ? 32'hFFC00000 : local_bb4_var__u65);
assign local_bb4_cast_after_negation_valid_out = 1'b1;
assign rnode_352to353_bb4__29_i437_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_352to353_bb4_or581_i466_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_352to353_bb4_and108_i493_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_div_inputs_ready;
 reg local_bb4_div_valid_out_NO_SHIFT_REG;
wire local_bb4_div_stall_in;
wire local_bb4_div_output_regs_ready;
wire [31:0] local_bb4_div;
 reg local_bb4_div_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_12_NO_SHIFT_REG;
wire local_bb4_div_causedstall;

acl_fp_div_s5 fp_module_local_bb4_div (
	.clock(clock),
	.dataa(local_bb4_cast_after_negation),
	.datab(input_wii_mul39),
	.enable(local_bb4_div_output_regs_ready),
	.result(local_bb4_div)
);


assign local_bb4_div_inputs_ready = 1'b1;
assign local_bb4_div_output_regs_ready = 1'b1;
assign local_bb4_cast_after_negation_stall_in = 1'b0;
assign local_bb4_div_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_div_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_div_output_regs_ready)
		begin
			local_bb4_div_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_div_valid_pipe_1_NO_SHIFT_REG <= local_bb4_div_valid_pipe_0_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_2_NO_SHIFT_REG <= local_bb4_div_valid_pipe_1_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_3_NO_SHIFT_REG <= local_bb4_div_valid_pipe_2_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_4_NO_SHIFT_REG <= local_bb4_div_valid_pipe_3_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_5_NO_SHIFT_REG <= local_bb4_div_valid_pipe_4_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_6_NO_SHIFT_REG <= local_bb4_div_valid_pipe_5_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_7_NO_SHIFT_REG <= local_bb4_div_valid_pipe_6_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_8_NO_SHIFT_REG <= local_bb4_div_valid_pipe_7_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_9_NO_SHIFT_REG <= local_bb4_div_valid_pipe_8_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_10_NO_SHIFT_REG <= local_bb4_div_valid_pipe_9_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_11_NO_SHIFT_REG <= local_bb4_div_valid_pipe_10_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_12_NO_SHIFT_REG <= local_bb4_div_valid_pipe_11_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_div_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_div_output_regs_ready)
		begin
			local_bb4_div_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_div_stall_in))
			begin
				local_bb4_div_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_call_i_div_inputs_ready;
 reg local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG;
wire local_bb4_call_i_div_stall_in_0;
 reg local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG;
wire local_bb4_call_i_div_stall_in_1;
wire local_bb4_call_i_div_output_regs_ready;
wire [31:0] local_bb4_call_i_div;
 reg local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_14_NO_SHIFT_REG;
wire local_bb4_call_i_div_causedstall;

acl_fp_exp_s5 fp_module_local_bb4_call_i_div (
	.clock(clock),
	.dataa(local_bb4_div),
	.enable(local_bb4_call_i_div_output_regs_ready),
	.result(local_bb4_call_i_div)
);


assign local_bb4_call_i_div_inputs_ready = 1'b1;
assign local_bb4_call_i_div_output_regs_ready = 1'b1;
assign local_bb4_div_stall_in = 1'b0;
assign local_bb4_call_i_div_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_14_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_call_i_div_output_regs_ready)
		begin
			local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_14_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_call_i_div_output_regs_ready)
		begin
			local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_call_i_div_stall_in_0))
			begin
				local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_call_i_div_stall_in_1))
			begin
				local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_astype_i_i_stall_local;
wire [31:0] local_bb4_astype_i_i;

assign local_bb4_astype_i_i = local_bb4_call_i_div;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u66_stall_local;
wire [31:0] local_bb4_var__u66;

assign local_bb4_var__u66 = local_bb4_call_i_div;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i_stall_local;
wire [31:0] local_bb4_and_i_i;

assign local_bb4_and_i_i = (local_bb4_astype_i_i & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i_i_stall_local;
wire local_bb4_cmp_i_i;

assign local_bb4_cmp_i_i = ((local_bb4_and_i_i & 32'h7F800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u67_stall_local;
wire [31:0] local_bb4_var__u67;

assign local_bb4_var__u67 = (local_bb4_cmp_i_i ? 32'h0 : local_bb4_var__u66);

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i222_stall_local;
wire [31:0] local_bb4_shr2_i222;

assign local_bb4_shr2_i222 = (local_bb4_var__u67 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i224_stall_local;
wire [31:0] local_bb4_xor_i224;

assign local_bb4_xor_i224 = (local_bb4_var__u67 ^ rnode_382to383_bb4_var__u50_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and6_i227_stall_local;
wire [31:0] local_bb4_and6_i227;

assign local_bb4_and6_i227 = (local_bb4_var__u67 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and3_i223_stall_local;
wire [31:0] local_bb4_and3_i223;

assign local_bb4_and3_i223 = ((local_bb4_shr2_i222 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_i233_stall_local;
wire local_bb4_lnot17_i233;

assign local_bb4_lnot17_i233 = ((local_bb4_and6_i227 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u68_stall_local;
wire [31:0] local_bb4_var__u68;

assign local_bb4_var__u68 = ((local_bb4_and6_i227 & 32'h7FFFFF) | (local_bb4_and_i221 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_or47_i255_stall_local;
wire [31:0] local_bb4_or47_i255;

assign local_bb4_or47_i255 = ((local_bb4_and6_i227 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot8_i229_stall_local;
wire local_bb4_lnot8_i229;

assign local_bb4_lnot8_i229 = ((local_bb4_and3_i223 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_i231_stall_local;
wire local_bb4_cmp11_i231;

assign local_bb4_cmp11_i231 = ((local_bb4_and3_i223 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u69_stall_local;
wire [31:0] local_bb4_var__u69;

assign local_bb4_var__u69 = ((local_bb4_and3_i223 & 32'hFF) | (local_bb4_and6_i227 & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i265_stall_local;
wire [31:0] local_bb4_add_i265;

assign local_bb4_add_i265 = ((local_bb4_and3_i223 & 32'hFF) + (local_bb4_and_i221 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u70_stall_local;
wire local_bb4_var__u70;

assign local_bb4_var__u70 = ((local_bb4_var__u68 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_conv1_i_i257_stall_local;
wire [63:0] local_bb4_conv1_i_i257;

assign local_bb4_conv1_i_i257[63:32] = 32'h0;
assign local_bb4_conv1_i_i257[31:0] = ((local_bb4_or47_i255 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i228_valid_out;
wire local_bb4_lnot_i228_stall_in;
wire local_bb4_cmp_i230_valid_out;
wire local_bb4_cmp_i230_stall_in;
wire local_bb4_add_i265_valid_out;
wire local_bb4_add_i265_stall_in;
wire local_bb4_var__u70_valid_out;
wire local_bb4_var__u70_stall_in;
wire local_bb4_xor_i224_valid_out;
wire local_bb4_xor_i224_stall_in;
wire local_bb4_lnot17_i233_valid_out;
wire local_bb4_lnot17_i233_stall_in;
wire local_bb4_lnot8_i229_valid_out;
wire local_bb4_lnot8_i229_stall_in;
wire local_bb4_cmp11_i231_valid_out;
wire local_bb4_cmp11_i231_stall_in;
wire local_bb4_var__u71_valid_out;
wire local_bb4_var__u71_stall_in;
wire local_bb4_conv1_i_i257_valid_out;
wire local_bb4_conv1_i_i257_stall_in;
wire local_bb4_var__u71_inputs_ready;
wire local_bb4_var__u71_stall_local;
wire local_bb4_var__u71;

assign local_bb4_var__u71_inputs_ready = (rnode_382to383_bb4_var__u50_0_valid_out_0_NO_SHIFT_REG & rnode_382to383_bb4_var__u50_0_valid_out_1_NO_SHIFT_REG & local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG & local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG);
assign local_bb4_var__u71 = ((local_bb4_var__u69 & 32'h7FFFFF) == 32'h0);
assign local_bb4_lnot_i228_valid_out = 1'b1;
assign local_bb4_cmp_i230_valid_out = 1'b1;
assign local_bb4_add_i265_valid_out = 1'b1;
assign local_bb4_var__u70_valid_out = 1'b1;
assign local_bb4_xor_i224_valid_out = 1'b1;
assign local_bb4_lnot17_i233_valid_out = 1'b1;
assign local_bb4_lnot8_i229_valid_out = 1'b1;
assign local_bb4_cmp11_i231_valid_out = 1'b1;
assign local_bb4_var__u71_valid_out = 1'b1;
assign local_bb4_conv1_i_i257_valid_out = 1'b1;
assign rnode_382to383_bb4_var__u50_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_382to383_bb4_var__u50_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign local_bb4_call_i_div_stall_in_1 = 1'b0;
assign local_bb4_call_i_div_stall_in_0 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_lnot_i228_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot_i228_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_lnot_i228_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_lnot_i228_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_lnot_i228_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_lnot_i228_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_lnot_i228_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_lnot_i228),
	.data_out(rnode_383to384_bb4_lnot_i228_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_lnot_i228_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_lnot_i228_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_lnot_i228_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_lnot_i228_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_lnot_i228_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot_i228_stall_in = 1'b0;
assign rnode_383to384_bb4_lnot_i228_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot_i228_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_lnot_i228_0_NO_SHIFT_REG = rnode_383to384_bb4_lnot_i228_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_lnot_i228_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_lnot_i228_1_NO_SHIFT_REG = rnode_383to384_bb4_lnot_i228_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_cmp_i230_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_3_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp_i230_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_cmp_i230_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_cmp_i230_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_cmp_i230_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_cmp_i230_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_cmp_i230_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_cmp_i230),
	.data_out(rnode_383to384_bb4_cmp_i230_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_cmp_i230_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_cmp_i230_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_cmp_i230_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_cmp_i230_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_cmp_i230_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp_i230_stall_in = 1'b0;
assign rnode_383to384_bb4_cmp_i230_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp_i230_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp_i230_0_NO_SHIFT_REG = rnode_383to384_bb4_cmp_i230_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp_i230_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp_i230_1_NO_SHIFT_REG = rnode_383to384_bb4_cmp_i230_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp_i230_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp_i230_2_NO_SHIFT_REG = rnode_383to384_bb4_cmp_i230_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp_i230_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp_i230_3_NO_SHIFT_REG = rnode_383to384_bb4_cmp_i230_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_add_i265_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb4_add_i265_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb4_add_i265_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_add_i265_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb4_add_i265_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_add_i265_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_add_i265_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_add_i265_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_add_i265_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_add_i265_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_add_i265_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_add_i265_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_add_i265_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in((local_bb4_add_i265 & 32'h1FF)),
	.data_out(rnode_383to384_bb4_add_i265_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_add_i265_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_add_i265_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb4_add_i265_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_add_i265_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_add_i265_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add_i265_stall_in = 1'b0;
assign rnode_383to384_bb4_add_i265_0_NO_SHIFT_REG = rnode_383to384_bb4_add_i265_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_add_i265_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_add_i265_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_var__u70_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u70_0_stall_in_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u70_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u70_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u70_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u70_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u70_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u70_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_var__u70_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_var__u70_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_var__u70_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_var__u70_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_var__u70_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_var__u70),
	.data_out(rnode_383to384_bb4_var__u70_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_var__u70_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_var__u70_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_var__u70_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_var__u70_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_var__u70_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u70_stall_in = 1'b0;
assign rnode_383to384_bb4_var__u70_0_NO_SHIFT_REG = rnode_383to384_bb4_var__u70_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_var__u70_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_var__u70_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb4_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb4_xor_i224_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_xor_i224_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_383to384_bb4_xor_i224_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_xor_i224_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_xor_i224_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_xor_i224_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_xor_i224_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_xor_i224_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_xor_i224_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_xor_i224_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_xor_i224_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i224),
	.data_out(rnode_383to384_bb4_xor_i224_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_xor_i224_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_xor_i224_0_reg_384_fifo.DATA_WIDTH = 32;
defparam rnode_383to384_bb4_xor_i224_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_xor_i224_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_xor_i224_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i224_stall_in = 1'b0;
assign rnode_383to384_bb4_xor_i224_0_NO_SHIFT_REG = rnode_383to384_bb4_xor_i224_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_xor_i224_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_lnot17_i233_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot17_i233_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_lnot17_i233_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_lnot17_i233_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_lnot17_i233_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_lnot17_i233_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_lnot17_i233_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_lnot17_i233),
	.data_out(rnode_383to384_bb4_lnot17_i233_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_lnot17_i233_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_lnot17_i233_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_lnot17_i233_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_lnot17_i233_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_lnot17_i233_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot17_i233_stall_in = 1'b0;
assign rnode_383to384_bb4_lnot17_i233_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot17_i233_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_lnot17_i233_0_NO_SHIFT_REG = rnode_383to384_bb4_lnot17_i233_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_lnot17_i233_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_lnot17_i233_1_NO_SHIFT_REG = rnode_383to384_bb4_lnot17_i233_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_lnot8_i229_0_valid_out_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot8_i229_0_stall_in_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot8_i229_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot8_i229_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot8_i229_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot8_i229_0_valid_out_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot8_i229_0_stall_in_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_lnot8_i229_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_lnot8_i229_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_lnot8_i229_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_lnot8_i229_0_stall_in_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_lnot8_i229_0_valid_out_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_lnot8_i229_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_lnot8_i229),
	.data_out(rnode_383to384_bb4_lnot8_i229_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_lnot8_i229_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_lnot8_i229_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_lnot8_i229_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_lnot8_i229_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_lnot8_i229_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot8_i229_stall_in = 1'b0;
assign rnode_383to384_bb4_lnot8_i229_0_NO_SHIFT_REG = rnode_383to384_bb4_lnot8_i229_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_lnot8_i229_0_stall_in_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot8_i229_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_cmp11_i231_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_3_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_in_4_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_4_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_valid_out_5_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_in_5_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_5_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_cmp11_i231_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_cmp11_i231_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_cmp11_i231_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_cmp11_i231_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_cmp11_i231_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_cmp11_i231_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_cmp11_i231),
	.data_out(rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_cmp11_i231_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_cmp11_i231_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_cmp11_i231_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_cmp11_i231_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_cmp11_i231_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp11_i231_stall_in = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp11_i231_0_NO_SHIFT_REG = rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp11_i231_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp11_i231_1_NO_SHIFT_REG = rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp11_i231_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp11_i231_2_NO_SHIFT_REG = rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp11_i231_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp11_i231_3_NO_SHIFT_REG = rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp11_i231_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp11_i231_4_NO_SHIFT_REG = rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_cmp11_i231_0_valid_out_5_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_cmp11_i231_5_NO_SHIFT_REG = rnode_383to384_bb4_cmp11_i231_0_reg_384_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_383to384_bb4_var__u71_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_1_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_2_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_reg_384_inputs_ready_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_valid_out_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_stall_in_0_reg_384_NO_SHIFT_REG;
 logic rnode_383to384_bb4_var__u71_0_stall_out_reg_384_NO_SHIFT_REG;

acl_data_fifo rnode_383to384_bb4_var__u71_0_reg_384_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_383to384_bb4_var__u71_0_reg_384_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_383to384_bb4_var__u71_0_stall_in_0_reg_384_NO_SHIFT_REG),
	.valid_out(rnode_383to384_bb4_var__u71_0_valid_out_0_reg_384_NO_SHIFT_REG),
	.stall_out(rnode_383to384_bb4_var__u71_0_stall_out_reg_384_NO_SHIFT_REG),
	.data_in(local_bb4_var__u71),
	.data_out(rnode_383to384_bb4_var__u71_0_reg_384_NO_SHIFT_REG)
);

defparam rnode_383to384_bb4_var__u71_0_reg_384_fifo.DEPTH = 1;
defparam rnode_383to384_bb4_var__u71_0_reg_384_fifo.DATA_WIDTH = 1;
defparam rnode_383to384_bb4_var__u71_0_reg_384_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_383to384_bb4_var__u71_0_reg_384_fifo.IMPL = "shift_reg";

assign rnode_383to384_bb4_var__u71_0_reg_384_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u71_stall_in = 1'b0;
assign rnode_383to384_bb4_var__u71_0_stall_in_0_reg_384_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_var__u71_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_var__u71_0_NO_SHIFT_REG = rnode_383to384_bb4_var__u71_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_var__u71_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_var__u71_1_NO_SHIFT_REG = rnode_383to384_bb4_var__u71_0_reg_384_NO_SHIFT_REG;
assign rnode_383to384_bb4_var__u71_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_var__u71_2_NO_SHIFT_REG = rnode_383to384_bb4_var__u71_0_reg_384_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_mul_i_i258_inputs_ready;
 reg local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG;
wire local_bb4_mul_i_i258_stall_in_0;
 reg local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i258_stall_in_1;
wire local_bb4_mul_i_i258_output_regs_ready;
wire [63:0] local_bb4_mul_i_i258;
 reg local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul_i_i258_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i258_causedstall;

acl_int_mult int_module_local_bb4_mul_i_i258 (
	.clock(clock),
	.dataa(((local_bb4_conv1_i_i257 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb4_conv_i_i256 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb4_mul_i_i258_output_regs_ready),
	.result(local_bb4_mul_i_i258)
);

defparam int_module_local_bb4_mul_i_i258.INPUT1_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i258.INPUT2_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i258.OUTPUT_WIDTH = 64;
defparam int_module_local_bb4_mul_i_i258.LATENCY = 3;
defparam int_module_local_bb4_mul_i_i258.SIGNED = 0;

assign local_bb4_mul_i_i258_inputs_ready = 1'b1;
assign local_bb4_mul_i_i258_output_regs_ready = 1'b1;
assign local_bb4_conv1_i_i257_stall_in = 1'b0;
assign local_bb4_conv_i_i256_stall_in = 1'b0;
assign local_bb4_mul_i_i258_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i258_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i258_output_regs_ready)
		begin
			local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i258_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i258_output_regs_ready)
		begin
			local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul_i_i258_stall_in_0))
			begin
				local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_mul_i_i258_stall_in_1))
			begin
				local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__28_i252_stall_local;
wire local_bb4__28_i252;

assign local_bb4__28_i252 = (rnode_383to384_bb4_cmp_i230_2_NO_SHIFT_REG & local_bb4_lnot14_not_i251);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb4_add_i265_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb4_add_i265_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb4_add_i265_0_NO_SHIFT_REG;
 logic rnode_384to385_bb4_add_i265_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to385_bb4_add_i265_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4_add_i265_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4_add_i265_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4_add_i265_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb4_add_i265_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb4_add_i265_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb4_add_i265_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb4_add_i265_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb4_add_i265_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in((rnode_383to384_bb4_add_i265_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_384to385_bb4_add_i265_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb4_add_i265_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb4_add_i265_0_reg_385_fifo.DATA_WIDTH = 32;
defparam rnode_384to385_bb4_add_i265_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb4_add_i265_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb4_add_i265_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_add_i265_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb4_add_i265_0_NO_SHIFT_REG = rnode_384to385_bb4_add_i265_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb4_add_i265_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb4_add_i265_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_384to387_bb4_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to387_bb4_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_384to387_bb4_xor_i224_0_NO_SHIFT_REG;
 logic rnode_384to387_bb4_xor_i224_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_384to387_bb4_xor_i224_0_reg_387_NO_SHIFT_REG;
 logic rnode_384to387_bb4_xor_i224_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_384to387_bb4_xor_i224_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_384to387_bb4_xor_i224_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_384to387_bb4_xor_i224_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to387_bb4_xor_i224_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to387_bb4_xor_i224_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_384to387_bb4_xor_i224_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_384to387_bb4_xor_i224_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_383to384_bb4_xor_i224_0_NO_SHIFT_REG),
	.data_out(rnode_384to387_bb4_xor_i224_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_384to387_bb4_xor_i224_0_reg_387_fifo.DEPTH = 3;
defparam rnode_384to387_bb4_xor_i224_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_384to387_bb4_xor_i224_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to387_bb4_xor_i224_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_384to387_bb4_xor_i224_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_383to384_bb4_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_384to387_bb4_xor_i224_0_NO_SHIFT_REG = rnode_384to387_bb4_xor_i224_0_reg_387_NO_SHIFT_REG;
assign rnode_384to387_bb4_xor_i224_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_384to387_bb4_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_not_i237_stall_local;
wire local_bb4_lnot17_not_i237;

assign local_bb4_lnot17_not_i237 = (rnode_383to384_bb4_lnot17_i233_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i283_valid_out;
wire local_bb4_reduction_0_i283_stall_in;
wire local_bb4_reduction_0_i283_inputs_ready;
wire local_bb4_reduction_0_i283_stall_local;
wire local_bb4_reduction_0_i283;

assign local_bb4_reduction_0_i283_inputs_ready = (rnode_383to384_bb4_lnot_i228_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb4_lnot8_i229_0_valid_out_NO_SHIFT_REG);
assign local_bb4_reduction_0_i283 = (rnode_383to384_bb4_lnot_i228_1_NO_SHIFT_REG | rnode_383to384_bb4_lnot8_i229_0_NO_SHIFT_REG);
assign local_bb4_reduction_0_i283_valid_out = 1'b1;
assign rnode_383to384_bb4_lnot_i228_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot8_i229_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge8_demorgan_i234_stall_local;
wire local_bb4_brmerge8_demorgan_i234;

assign local_bb4_brmerge8_demorgan_i234 = (rnode_383to384_bb4_cmp11_i231_0_NO_SHIFT_REG & rnode_383to384_bb4_lnot17_i233_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_not_i238_stall_local;
wire local_bb4_cmp11_not_i238;

assign local_bb4_cmp11_not_i238 = (rnode_383to384_bb4_cmp11_i231_2_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u72_valid_out;
wire local_bb4_var__u72_stall_in;
wire local_bb4_var__u72_inputs_ready;
wire local_bb4_var__u72_stall_local;
wire local_bb4_var__u72;

assign local_bb4_var__u72_inputs_ready = (rnode_383to384_bb4_cmp_i230_0_valid_out_3_NO_SHIFT_REG & rnode_383to384_bb4_cmp11_i231_0_valid_out_5_NO_SHIFT_REG);
assign local_bb4_var__u72 = (rnode_383to384_bb4_cmp_i230_3_NO_SHIFT_REG | rnode_383to384_bb4_cmp11_i231_5_NO_SHIFT_REG);
assign local_bb4_var__u72_valid_out = 1'b1;
assign rnode_383to384_bb4_cmp_i230_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_stall_in_5_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_i241_stall_local;
wire local_bb4__mux_mux_i241;

assign local_bb4__mux_mux_i241 = (rnode_383to384_bb4_var__u71_1_NO_SHIFT_REG | rnode_383to384_bb4_cmp11_i231_3_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__not_i243_stall_local;
wire local_bb4__not_i243;

assign local_bb4__not_i243 = (rnode_383to384_bb4_var__u71_2_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_conv3_i_i259_stall_local;
wire [31:0] local_bb4_conv3_i_i259;
wire [63:0] local_bb4_conv3_i_i259$ps;

assign local_bb4_conv3_i_i259$ps = (local_bb4_mul_i_i258 & 64'hFFFFFFFFFFFF);
assign local_bb4_conv3_i_i259 = local_bb4_conv3_i_i259$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u73_stall_local;
wire [63:0] local_bb4_var__u73;

assign local_bb4_var__u73 = ((local_bb4_mul_i_i258 & 64'hFFFFFFFFFFFF) >> 64'h18);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_385to386_bb4_add_i265_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb4_add_i265_0_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb4_add_i265_1_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb4_add_i265_2_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_385to386_bb4_add_i265_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_valid_out_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_stall_in_0_reg_386_NO_SHIFT_REG;
 logic rnode_385to386_bb4_add_i265_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_385to386_bb4_add_i265_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to386_bb4_add_i265_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to386_bb4_add_i265_0_stall_in_0_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_385to386_bb4_add_i265_0_valid_out_0_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_385to386_bb4_add_i265_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in((rnode_384to385_bb4_add_i265_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_385to386_bb4_add_i265_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_385to386_bb4_add_i265_0_reg_386_fifo.DEPTH = 1;
defparam rnode_385to386_bb4_add_i265_0_reg_386_fifo.DATA_WIDTH = 32;
defparam rnode_385to386_bb4_add_i265_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to386_bb4_add_i265_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_385to386_bb4_add_i265_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb4_add_i265_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb4_add_i265_0_stall_in_0_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb4_add_i265_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb4_add_i265_0_NO_SHIFT_REG = rnode_385to386_bb4_add_i265_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb4_add_i265_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb4_add_i265_1_NO_SHIFT_REG = rnode_385to386_bb4_add_i265_0_reg_386_NO_SHIFT_REG;
assign rnode_385to386_bb4_add_i265_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_385to386_bb4_add_i265_2_NO_SHIFT_REG = rnode_385to386_bb4_add_i265_0_reg_386_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_xor_i224_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_xor_i224_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_xor_i224_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_xor_i224_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_xor_i224_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_xor_i224_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_xor_i224_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_xor_i224_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_xor_i224_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_xor_i224_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_xor_i224_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_384to387_bb4_xor_i224_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb4_xor_i224_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_xor_i224_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_xor_i224_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb4_xor_i224_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_xor_i224_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_xor_i224_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_384to387_bb4_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_xor_i224_0_NO_SHIFT_REG = rnode_387to388_bb4_xor_i224_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_xor_i224_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb4_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_384to385_bb4_reduction_0_i283_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb4_reduction_0_i283_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4_reduction_0_i283_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4_reduction_0_i283_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4_reduction_0_i283_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb4_reduction_0_i283_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb4_reduction_0_i283_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb4_reduction_0_i283_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb4_reduction_0_i283_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb4_reduction_0_i283_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_0_i283),
	.data_out(rnode_384to385_bb4_reduction_0_i283_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb4_reduction_0_i283_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb4_reduction_0_i283_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb4_reduction_0_i283_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb4_reduction_0_i283_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb4_reduction_0_i283_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_0_i283_stall_in = 1'b0;
assign rnode_384to385_bb4_reduction_0_i283_0_NO_SHIFT_REG = rnode_384to385_bb4_reduction_0_i283_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb4_reduction_0_i283_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge10_demorgan_i235_stall_local;
wire local_bb4_brmerge10_demorgan_i235;

assign local_bb4_brmerge10_demorgan_i235 = (local_bb4_brmerge8_demorgan_i234 & rnode_383to384_bb4_lnot_i228_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__mux9_mux_i236_stall_local;
wire local_bb4__mux9_mux_i236;

assign local_bb4__mux9_mux_i236 = (local_bb4_brmerge8_demorgan_i234 ^ rnode_383to384_bb4_cmp11_i231_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge3_i239_stall_local;
wire local_bb4_brmerge3_i239;

assign local_bb4_brmerge3_i239 = (rnode_383to384_bb4_var__u71_0_NO_SHIFT_REG | local_bb4_cmp11_not_i238);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_384to386_bb4_var__u72_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to386_bb4_var__u72_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to386_bb4_var__u72_0_NO_SHIFT_REG;
 logic rnode_384to386_bb4_var__u72_0_reg_386_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to386_bb4_var__u72_0_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb4_var__u72_0_valid_out_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb4_var__u72_0_stall_in_reg_386_NO_SHIFT_REG;
 logic rnode_384to386_bb4_var__u72_0_stall_out_reg_386_NO_SHIFT_REG;

acl_data_fifo rnode_384to386_bb4_var__u72_0_reg_386_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to386_bb4_var__u72_0_reg_386_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to386_bb4_var__u72_0_stall_in_reg_386_NO_SHIFT_REG),
	.valid_out(rnode_384to386_bb4_var__u72_0_valid_out_reg_386_NO_SHIFT_REG),
	.stall_out(rnode_384to386_bb4_var__u72_0_stall_out_reg_386_NO_SHIFT_REG),
	.data_in(local_bb4_var__u72),
	.data_out(rnode_384to386_bb4_var__u72_0_reg_386_NO_SHIFT_REG)
);

defparam rnode_384to386_bb4_var__u72_0_reg_386_fifo.DEPTH = 2;
defparam rnode_384to386_bb4_var__u72_0_reg_386_fifo.DATA_WIDTH = 1;
defparam rnode_384to386_bb4_var__u72_0_reg_386_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to386_bb4_var__u72_0_reg_386_fifo.IMPL = "shift_reg";

assign rnode_384to386_bb4_var__u72_0_reg_386_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u72_stall_in = 1'b0;
assign rnode_384to386_bb4_var__u72_0_NO_SHIFT_REG = rnode_384to386_bb4_var__u72_0_reg_386_NO_SHIFT_REG;
assign rnode_384to386_bb4_var__u72_0_stall_in_reg_386_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb4_var__u72_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i244_stall_local;
wire local_bb4_reduction_3_i244;

assign local_bb4_reduction_3_i244 = (rnode_383to384_bb4_cmp11_i231_4_NO_SHIFT_REG & local_bb4__not_i243);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i16_i262_stall_local;
wire [31:0] local_bb4_shr_i16_i262;

assign local_bb4_shr_i16_i262 = (local_bb4_conv3_i_i259 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i18_i264_stall_local;
wire [31:0] local_bb4_shl1_i18_i264;

assign local_bb4_shl1_i18_i264 = (local_bb4_conv3_i_i259 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u74_stall_local;
wire [31:0] local_bb4_var__u74;

assign local_bb4_var__u74 = (local_bb4_conv3_i_i259 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i_i272_stall_local;
wire [31:0] local_bb4_shl1_i_i272;

assign local_bb4_shl1_i_i272 = (local_bb4_conv3_i_i259 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb4__tr_i260_stall_local;
wire [31:0] local_bb4__tr_i260;
wire [63:0] local_bb4__tr_i260$ps;

assign local_bb4__tr_i260$ps = (local_bb4_var__u73 & 64'hFFFFFF);
assign local_bb4__tr_i260 = local_bb4__tr_i260$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_inc_i268_stall_local;
wire [31:0] local_bb4_inc_i268;

assign local_bb4_inc_i268 = ((rnode_385to386_bb4_add_i265_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp50_not_i273_stall_local;
wire local_bb4_cmp50_not_i273;

assign local_bb4_cmp50_not_i273 = ((rnode_385to386_bb4_add_i265_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4_and4_i225_stall_local;
wire [31:0] local_bb4_and4_i225;

assign local_bb4_and4_i225 = (rnode_387to388_bb4_xor_i224_0_NO_SHIFT_REG & 32'h80000000);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_385to387_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_385to387_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_385to387_bb4_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_385to387_bb4_reduction_0_i283_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_385to387_bb4_reduction_0_i283_0_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb4_reduction_0_i283_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb4_reduction_0_i283_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb4_reduction_0_i283_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_385to387_bb4_reduction_0_i283_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to387_bb4_reduction_0_i283_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to387_bb4_reduction_0_i283_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_385to387_bb4_reduction_0_i283_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_385to387_bb4_reduction_0_i283_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_384to385_bb4_reduction_0_i283_0_NO_SHIFT_REG),
	.data_out(rnode_385to387_bb4_reduction_0_i283_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_385to387_bb4_reduction_0_i283_0_reg_387_fifo.DEPTH = 2;
defparam rnode_385to387_bb4_reduction_0_i283_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_385to387_bb4_reduction_0_i283_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to387_bb4_reduction_0_i283_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_385to387_bb4_reduction_0_i283_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to387_bb4_reduction_0_i283_0_NO_SHIFT_REG = rnode_385to387_bb4_reduction_0_i283_0_reg_387_NO_SHIFT_REG;
assign rnode_385to387_bb4_reduction_0_i283_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_385to387_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__26_demorgan_i249_stall_local;
wire local_bb4__26_demorgan_i249;

assign local_bb4__26_demorgan_i249 = (rnode_383to384_bb4_cmp_i230_1_NO_SHIFT_REG | local_bb4_brmerge10_demorgan_i235);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge5_i240_stall_local;
wire local_bb4_brmerge5_i240;

assign local_bb4_brmerge5_i240 = (local_bb4_brmerge3_i239 | local_bb4_lnot17_not_i237);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i245_stall_local;
wire local_bb4_reduction_5_i245;

assign local_bb4_reduction_5_i245 = (rnode_383to384_bb4_lnot14_i232_0_NO_SHIFT_REG & local_bb4_reduction_3_i244);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i270_stall_local;
wire [31:0] local_bb4_shr_i_i270;

assign local_bb4_shr_i_i270 = ((local_bb4_var__u74 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i15_i261_stall_local;
wire [31:0] local_bb4_shl_i15_i261;

assign local_bb4_shl_i15_i261 = ((local_bb4__tr_i260 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb4_and48_i266_stall_local;
wire [31:0] local_bb4_and48_i266;

assign local_bb4_and48_i266 = ((local_bb4__tr_i260 & 32'hFFFFFF) & 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb4_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_reduction_0_i283_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb4_reduction_0_i283_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_reduction_0_i283_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_reduction_0_i283_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_reduction_0_i283_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_reduction_0_i283_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_reduction_0_i283_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_reduction_0_i283_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_reduction_0_i283_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_reduction_0_i283_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_385to387_bb4_reduction_0_i283_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb4_reduction_0_i283_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_reduction_0_i283_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_reduction_0_i283_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb4_reduction_0_i283_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_reduction_0_i283_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_reduction_0_i283_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_385to387_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_reduction_0_i283_0_NO_SHIFT_REG = rnode_387to388_bb4_reduction_0_i283_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_reduction_0_i283_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_mux_i242_stall_local;
wire local_bb4__mux_mux_mux_i242;

assign local_bb4__mux_mux_mux_i242 = (local_bb4_brmerge5_i240 & local_bb4__mux_mux_i241);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i246_stall_local;
wire local_bb4_reduction_6_i246;

assign local_bb4_reduction_6_i246 = (rnode_383to384_bb4_var__u70_0_NO_SHIFT_REG & local_bb4_reduction_5_i245);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i17_i263_stall_local;
wire [31:0] local_bb4_or_i17_i263;

assign local_bb4_or_i17_i263 = ((local_bb4_shl_i15_i261 & 32'hFFFF00) | (local_bb4_shr_i16_i262 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool49_i267_stall_local;
wire local_bb4_tobool49_i267;

assign local_bb4_tobool49_i267 = ((local_bb4_and48_i266 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i247_stall_local;
wire local_bb4__24_i247;

assign local_bb4__24_i247 = (rnode_383to384_bb4_cmp_i230_0_NO_SHIFT_REG ? local_bb4_reduction_6_i246 : local_bb4_brmerge10_demorgan_i235);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_i269_stall_local;
wire [31:0] local_bb4_shl_i_i269;

assign local_bb4_shl_i_i269 = ((local_bb4_or_i17_i263 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__31_i274_stall_local;
wire local_bb4__31_i274;

assign local_bb4__31_i274 = (local_bb4_tobool49_i267 & local_bb4_cmp50_not_i273);

// This section implements an unregistered operation.
// 
wire local_bb4__25_i248_stall_local;
wire local_bb4__25_i248;

assign local_bb4__25_i248 = (local_bb4__24_i247 ? rnode_383to384_bb4_lnot14_i232_1_NO_SHIFT_REG : local_bb4__mux_mux_mux_i242);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i271_stall_local;
wire [31:0] local_bb4_or_i_i271;

assign local_bb4_or_i_i271 = ((local_bb4_shl_i_i269 & 32'h1FFFFFE) | (local_bb4_shr_i_i270 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i275_stall_local;
wire [31:0] local_bb4__32_i275;

assign local_bb4__32_i275 = (local_bb4__31_i274 ? (local_bb4_shl1_i_i272 & 32'hFFFFFE00) : (local_bb4_shl1_i18_i264 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__36_i279_stall_local;
wire [31:0] local_bb4__36_i279;

assign local_bb4__36_i279 = (local_bb4__31_i274 ? (rnode_385to386_bb4_add_i265_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i250_stall_local;
wire local_bb4__27_i250;

assign local_bb4__27_i250 = (local_bb4__26_demorgan_i249 ? local_bb4__25_i248 : local_bb4__mux9_mux_i236);

// This section implements an unregistered operation.
// 
wire local_bb4__34_i277_stall_local;
wire [31:0] local_bb4__34_i277;

assign local_bb4__34_i277 = (local_bb4__31_i274 ? (local_bb4_or_i_i271 & 32'h1FFFFFF) : (local_bb4_or_i17_i263 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i276_stall_local;
wire [31:0] local_bb4__33_i276;

assign local_bb4__33_i276 = (local_bb4_tobool49_i267 ? (local_bb4__32_i275 & 32'hFFFFFF00) : (local_bb4_shl1_i18_i264 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__37_i280_stall_local;
wire [31:0] local_bb4__37_i280;

assign local_bb4__37_i280 = (local_bb4_tobool49_i267 ? (local_bb4__36_i279 & 32'h1FF) : (local_bb4_inc_i268 & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb4__29_i253_valid_out;
wire local_bb4__29_i253_stall_in;
wire local_bb4__29_i253_inputs_ready;
wire local_bb4__29_i253_stall_local;
wire local_bb4__29_i253;

assign local_bb4__29_i253_inputs_ready = (rnode_383to384_bb4_lnot14_i232_0_valid_out_0_NO_SHIFT_REG & rnode_383to384_bb4_var__u70_0_valid_out_NO_SHIFT_REG & rnode_383to384_bb4_lnot14_i232_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb4_lnot_i228_0_valid_out_0_NO_SHIFT_REG & rnode_383to384_bb4_cmp_i230_0_valid_out_0_NO_SHIFT_REG & rnode_383to384_bb4_cmp_i230_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb4_lnot14_i232_0_valid_out_2_NO_SHIFT_REG & rnode_383to384_bb4_cmp_i230_0_valid_out_2_NO_SHIFT_REG & rnode_383to384_bb4_cmp11_i231_0_valid_out_0_NO_SHIFT_REG & rnode_383to384_bb4_lnot17_i233_0_valid_out_0_NO_SHIFT_REG & rnode_383to384_bb4_cmp11_i231_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb4_cmp11_i231_0_valid_out_4_NO_SHIFT_REG & rnode_383to384_bb4_var__u71_0_valid_out_2_NO_SHIFT_REG & rnode_383to384_bb4_lnot17_i233_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb4_var__u71_0_valid_out_1_NO_SHIFT_REG & rnode_383to384_bb4_cmp11_i231_0_valid_out_3_NO_SHIFT_REG & rnode_383to384_bb4_cmp11_i231_0_valid_out_2_NO_SHIFT_REG & rnode_383to384_bb4_var__u71_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__29_i253 = (local_bb4__28_i252 | local_bb4__27_i250);
assign local_bb4__29_i253_valid_out = 1'b1;
assign rnode_383to384_bb4_lnot14_i232_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_var__u70_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot14_i232_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot_i228_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp_i230_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp_i230_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot14_i232_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp_i230_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot17_i233_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_var__u71_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_lnot17_i233_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_var__u71_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_cmp11_i231_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_383to384_bb4_var__u71_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__35_i278_stall_local;
wire [31:0] local_bb4__35_i278;

assign local_bb4__35_i278 = (local_bb4_tobool49_i267 ? (local_bb4__34_i277 & 32'h1FFFFFF) : (local_bb4_or_i17_i263 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp53_i281_stall_local;
wire local_bb4_cmp53_i281;

assign local_bb4_cmp53_i281 = ((local_bb4__37_i280 & 32'h3FF) > 32'h17D);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_384to385_bb4__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_384to385_bb4__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_384to385_bb4__29_i253_0_NO_SHIFT_REG;
 logic rnode_384to385_bb4__29_i253_0_reg_385_inputs_ready_NO_SHIFT_REG;
 logic rnode_384to385_bb4__29_i253_0_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4__29_i253_0_valid_out_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4__29_i253_0_stall_in_reg_385_NO_SHIFT_REG;
 logic rnode_384to385_bb4__29_i253_0_stall_out_reg_385_NO_SHIFT_REG;

acl_data_fifo rnode_384to385_bb4__29_i253_0_reg_385_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_384to385_bb4__29_i253_0_reg_385_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_384to385_bb4__29_i253_0_stall_in_reg_385_NO_SHIFT_REG),
	.valid_out(rnode_384to385_bb4__29_i253_0_valid_out_reg_385_NO_SHIFT_REG),
	.stall_out(rnode_384to385_bb4__29_i253_0_stall_out_reg_385_NO_SHIFT_REG),
	.data_in(local_bb4__29_i253),
	.data_out(rnode_384to385_bb4__29_i253_0_reg_385_NO_SHIFT_REG)
);

defparam rnode_384to385_bb4__29_i253_0_reg_385_fifo.DEPTH = 1;
defparam rnode_384to385_bb4__29_i253_0_reg_385_fifo.DATA_WIDTH = 1;
defparam rnode_384to385_bb4__29_i253_0_reg_385_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_384to385_bb4__29_i253_0_reg_385_fifo.IMPL = "shift_reg";

assign rnode_384to385_bb4__29_i253_0_reg_385_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__29_i253_stall_in = 1'b0;
assign rnode_384to385_bb4__29_i253_0_NO_SHIFT_REG = rnode_384to385_bb4__29_i253_0_reg_385_NO_SHIFT_REG;
assign rnode_384to385_bb4__29_i253_0_stall_in_reg_385_NO_SHIFT_REG = 1'b0;
assign rnode_384to385_bb4__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i286_stall_local;
wire [31:0] local_bb4_and75_i286;

assign local_bb4_and75_i286 = ((local_bb4__35_i278 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and83_i292_stall_local;
wire [31:0] local_bb4_and83_i292;

assign local_bb4_and83_i292 = ((local_bb4__35_i278 & 32'h1FFFFFF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i276_valid_out;
wire local_bb4__33_i276_stall_in;
wire local_bb4__37_i280_valid_out_1;
wire local_bb4__37_i280_stall_in_1;
wire local_bb4_and75_i286_valid_out;
wire local_bb4_and75_i286_stall_in;
wire local_bb4_and83_i292_valid_out;
wire local_bb4_and83_i292_stall_in;
wire local_bb4_or581_i282_valid_out;
wire local_bb4_or581_i282_stall_in;
wire local_bb4_or581_i282_inputs_ready;
wire local_bb4_or581_i282_stall_local;
wire local_bb4_or581_i282;

assign local_bb4_or581_i282_inputs_ready = (local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG & local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG & rnode_385to386_bb4_add_i265_0_valid_out_1_NO_SHIFT_REG & rnode_385to386_bb4_add_i265_0_valid_out_0_NO_SHIFT_REG & rnode_385to386_bb4_add_i265_0_valid_out_2_NO_SHIFT_REG & rnode_384to386_bb4_var__u72_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or581_i282 = (rnode_384to386_bb4_var__u72_0_NO_SHIFT_REG | local_bb4_cmp53_i281);
assign local_bb4__33_i276_valid_out = 1'b1;
assign local_bb4__37_i280_valid_out_1 = 1'b1;
assign local_bb4_and75_i286_valid_out = 1'b1;
assign local_bb4_and83_i292_valid_out = 1'b1;
assign local_bb4_or581_i282_valid_out = 1'b1;
assign local_bb4_mul_i_i258_stall_in_0 = 1'b0;
assign local_bb4_mul_i_i258_stall_in_1 = 1'b0;
assign rnode_385to386_bb4_add_i265_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb4_add_i265_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_385to386_bb4_add_i265_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_384to386_bb4_var__u72_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_385to387_bb4__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_385to387_bb4__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_385to387_bb4__29_i253_0_NO_SHIFT_REG;
 logic rnode_385to387_bb4__29_i253_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic rnode_385to387_bb4__29_i253_0_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb4__29_i253_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb4__29_i253_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_385to387_bb4__29_i253_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_385to387_bb4__29_i253_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_385to387_bb4__29_i253_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_385to387_bb4__29_i253_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_385to387_bb4__29_i253_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_385to387_bb4__29_i253_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in(rnode_384to385_bb4__29_i253_0_NO_SHIFT_REG),
	.data_out(rnode_385to387_bb4__29_i253_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_385to387_bb4__29_i253_0_reg_387_fifo.DEPTH = 2;
defparam rnode_385to387_bb4__29_i253_0_reg_387_fifo.DATA_WIDTH = 1;
defparam rnode_385to387_bb4__29_i253_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_385to387_bb4__29_i253_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_385to387_bb4__29_i253_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_384to385_bb4__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_385to387_bb4__29_i253_0_NO_SHIFT_REG = rnode_385to387_bb4__29_i253_0_reg_387_NO_SHIFT_REG;
assign rnode_385to387_bb4__29_i253_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_385to387_bb4__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb4__33_i276_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to387_bb4__33_i276_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4__33_i276_0_NO_SHIFT_REG;
 logic rnode_386to387_bb4__33_i276_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to387_bb4__33_i276_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4__33_i276_1_NO_SHIFT_REG;
 logic rnode_386to387_bb4__33_i276_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4__33_i276_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4__33_i276_0_valid_out_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4__33_i276_0_stall_in_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4__33_i276_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb4__33_i276_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb4__33_i276_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb4__33_i276_0_stall_in_0_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb4__33_i276_0_valid_out_0_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb4__33_i276_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in((local_bb4__33_i276 & 32'hFFFFFF00)),
	.data_out(rnode_386to387_bb4__33_i276_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb4__33_i276_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb4__33_i276_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb4__33_i276_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb4__33_i276_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb4__33_i276_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__33_i276_stall_in = 1'b0;
assign rnode_386to387_bb4__33_i276_0_stall_in_0_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb4__33_i276_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb4__33_i276_0_NO_SHIFT_REG = rnode_386to387_bb4__33_i276_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb4__33_i276_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb4__33_i276_1_NO_SHIFT_REG = rnode_386to387_bb4__33_i276_0_reg_387_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb4__37_i280_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4__37_i280_0_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4__37_i280_1_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4__37_i280_2_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4__37_i280_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_valid_out_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_stall_in_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4__37_i280_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb4__37_i280_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb4__37_i280_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb4__37_i280_0_stall_in_0_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb4__37_i280_0_valid_out_0_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb4__37_i280_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in((local_bb4__37_i280 & 32'h3FF)),
	.data_out(rnode_386to387_bb4__37_i280_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb4__37_i280_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb4__37_i280_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb4__37_i280_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb4__37_i280_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb4__37_i280_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__37_i280_stall_in_1 = 1'b0;
assign rnode_386to387_bb4__37_i280_0_stall_in_0_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb4__37_i280_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb4__37_i280_0_NO_SHIFT_REG = rnode_386to387_bb4__37_i280_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb4__37_i280_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb4__37_i280_1_NO_SHIFT_REG = rnode_386to387_bb4__37_i280_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb4__37_i280_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_386to387_bb4__37_i280_2_NO_SHIFT_REG = rnode_386to387_bb4__37_i280_0_reg_387_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb4_and75_i286_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and75_i286_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4_and75_i286_0_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and75_i286_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4_and75_i286_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and75_i286_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and75_i286_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and75_i286_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb4_and75_i286_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb4_and75_i286_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb4_and75_i286_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb4_and75_i286_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb4_and75_i286_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in((local_bb4_and75_i286 & 32'h7FFFFF)),
	.data_out(rnode_386to387_bb4_and75_i286_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb4_and75_i286_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb4_and75_i286_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb4_and75_i286_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb4_and75_i286_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb4_and75_i286_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and75_i286_stall_in = 1'b0;
assign rnode_386to387_bb4_and75_i286_0_NO_SHIFT_REG = rnode_386to387_bb4_and75_i286_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb4_and75_i286_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb4_and75_i286_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_386to387_bb4_and83_i292_0_valid_out_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and83_i292_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4_and83_i292_0_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and83_i292_0_reg_387_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_386to387_bb4_and83_i292_0_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and83_i292_0_valid_out_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and83_i292_0_stall_in_reg_387_NO_SHIFT_REG;
 logic rnode_386to387_bb4_and83_i292_0_stall_out_reg_387_NO_SHIFT_REG;

acl_data_fifo rnode_386to387_bb4_and83_i292_0_reg_387_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to387_bb4_and83_i292_0_reg_387_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to387_bb4_and83_i292_0_stall_in_reg_387_NO_SHIFT_REG),
	.valid_out(rnode_386to387_bb4_and83_i292_0_valid_out_reg_387_NO_SHIFT_REG),
	.stall_out(rnode_386to387_bb4_and83_i292_0_stall_out_reg_387_NO_SHIFT_REG),
	.data_in((local_bb4_and83_i292 & 32'h1)),
	.data_out(rnode_386to387_bb4_and83_i292_0_reg_387_NO_SHIFT_REG)
);

defparam rnode_386to387_bb4_and83_i292_0_reg_387_fifo.DEPTH = 1;
defparam rnode_386to387_bb4_and83_i292_0_reg_387_fifo.DATA_WIDTH = 32;
defparam rnode_386to387_bb4_and83_i292_0_reg_387_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to387_bb4_and83_i292_0_reg_387_fifo.IMPL = "shift_reg";

assign rnode_386to387_bb4_and83_i292_0_reg_387_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and83_i292_stall_in = 1'b0;
assign rnode_386to387_bb4_and83_i292_0_NO_SHIFT_REG = rnode_386to387_bb4_and83_i292_0_reg_387_NO_SHIFT_REG;
assign rnode_386to387_bb4_and83_i292_0_stall_in_reg_387_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb4_and83_i292_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_386to388_bb4_or581_i282_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_1_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_reg_388_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_valid_out_0_reg_388_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_stall_in_0_reg_388_NO_SHIFT_REG;
 logic rnode_386to388_bb4_or581_i282_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_386to388_bb4_or581_i282_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_386to388_bb4_or581_i282_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_386to388_bb4_or581_i282_0_stall_in_0_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_386to388_bb4_or581_i282_0_valid_out_0_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_386to388_bb4_or581_i282_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb4_or581_i282),
	.data_out(rnode_386to388_bb4_or581_i282_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_386to388_bb4_or581_i282_0_reg_388_fifo.DEPTH = 2;
defparam rnode_386to388_bb4_or581_i282_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_386to388_bb4_or581_i282_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_386to388_bb4_or581_i282_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_386to388_bb4_or581_i282_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or581_i282_stall_in = 1'b0;
assign rnode_386to388_bb4_or581_i282_0_stall_in_0_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_386to388_bb4_or581_i282_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_386to388_bb4_or581_i282_0_NO_SHIFT_REG = rnode_386to388_bb4_or581_i282_0_reg_388_NO_SHIFT_REG;
assign rnode_386to388_bb4_or581_i282_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_386to388_bb4_or581_i282_1_NO_SHIFT_REG = rnode_386to388_bb4_or581_i282_0_reg_388_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb4__29_i253_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4__29_i253_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb4__29_i253_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4__29_i253_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4__29_i253_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4__29_i253_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4__29_i253_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4__29_i253_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4__29_i253_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4__29_i253_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4__29_i253_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(rnode_385to387_bb4__29_i253_0_NO_SHIFT_REG),
	.data_out(rnode_387to388_bb4__29_i253_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4__29_i253_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4__29_i253_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb4__29_i253_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4__29_i253_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4__29_i253_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_385to387_bb4__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4__29_i253_0_NO_SHIFT_REG = rnode_387to388_bb4__29_i253_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4__29_i253_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i291_stall_local;
wire local_bb4_cmp77_i291;

assign local_bb4_cmp77_i291 = ((rnode_386to387_bb4__33_i276_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u75_stall_local;
wire local_bb4_var__u75;

assign local_bb4_var__u75 = ($signed((rnode_386to387_bb4__33_i276_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp68_i285_valid_out;
wire local_bb4_cmp68_i285_stall_in;
wire local_bb4_cmp68_i285_inputs_ready;
wire local_bb4_cmp68_i285_stall_local;
wire local_bb4_cmp68_i285;

assign local_bb4_cmp68_i285_inputs_ready = rnode_386to387_bb4__37_i280_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_cmp68_i285 = ((rnode_386to387_bb4__37_i280_0_NO_SHIFT_REG & 32'h3FF) < 32'h80);
assign local_bb4_cmp68_i285_valid_out = 1'b1;
assign rnode_386to387_bb4__37_i280_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i287_stall_local;
wire [31:0] local_bb4_sub_i287;

assign local_bb4_sub_i287 = ((rnode_386to387_bb4__37_i280_1_NO_SHIFT_REG & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp71_not_i302_valid_out;
wire local_bb4_cmp71_not_i302_stall_in;
wire local_bb4_cmp71_not_i302_inputs_ready;
wire local_bb4_cmp71_not_i302_stall_local;
wire local_bb4_cmp71_not_i302;

assign local_bb4_cmp71_not_i302_inputs_ready = rnode_386to387_bb4__37_i280_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_cmp71_not_i302 = ((rnode_386to387_bb4__37_i280_2_NO_SHIFT_REG & 32'h3FF) != 32'h7F);
assign local_bb4_cmp71_not_i302_valid_out = 1'b1;
assign rnode_386to387_bb4__37_i280_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool84_i293_stall_local;
wire local_bb4_tobool84_i293;

assign local_bb4_tobool84_i293 = ((rnode_386to387_bb4_and83_i292_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i284_stall_local;
wire local_bb4_reduction_2_i284;

assign local_bb4_reduction_2_i284 = (rnode_387to388_bb4_reduction_0_i283_0_NO_SHIFT_REG | rnode_386to388_bb4_or581_i282_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cond111_i310_stall_local;
wire [31:0] local_bb4_cond111_i310;

assign local_bb4_cond111_i310 = (rnode_386to388_bb4_or581_i282_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_cmp68_i285_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp68_i285_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp68_i285_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp68_i285_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp68_i285_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp68_i285_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp68_i285_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp68_i285_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_cmp68_i285_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_cmp68_i285_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_cmp68_i285_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_cmp68_i285_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_cmp68_i285_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb4_cmp68_i285),
	.data_out(rnode_387to388_bb4_cmp68_i285_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_cmp68_i285_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_cmp68_i285_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb4_cmp68_i285_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_cmp68_i285_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_cmp68_i285_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp68_i285_stall_in = 1'b0;
assign rnode_387to388_bb4_cmp68_i285_0_NO_SHIFT_REG = rnode_387to388_bb4_cmp68_i285_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_cmp68_i285_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_cmp68_i285_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and74_i288_stall_local;
wire [31:0] local_bb4_and74_i288;

assign local_bb4_and74_i288 = ((local_bb4_sub_i287 & 32'hFF800000) + 32'h40800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_cmp71_not_i302_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp71_not_i302_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp71_not_i302_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp71_not_i302_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp71_not_i302_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp71_not_i302_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp71_not_i302_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_cmp71_not_i302_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_cmp71_not_i302_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_cmp71_not_i302_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_cmp71_not_i302_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_cmp71_not_i302_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_cmp71_not_i302_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb4_cmp71_not_i302),
	.data_out(rnode_387to388_bb4_cmp71_not_i302_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_cmp71_not_i302_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_cmp71_not_i302_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb4_cmp71_not_i302_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_cmp71_not_i302_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_cmp71_not_i302_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp71_not_i302_stall_in = 1'b0;
assign rnode_387to388_bb4_cmp71_not_i302_0_NO_SHIFT_REG = rnode_387to388_bb4_cmp71_not_i302_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_cmp71_not_i302_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_cmp71_not_i302_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__39_i294_stall_local;
wire local_bb4__39_i294;

assign local_bb4__39_i294 = (local_bb4_tobool84_i293 & local_bb4_var__u75);

// This section implements an unregistered operation.
// 
wire local_bb4_conv101_i305_stall_local;
wire [31:0] local_bb4_conv101_i305;

assign local_bb4_conv101_i305[31:1] = 31'h0;
assign local_bb4_conv101_i305[0] = local_bb4_reduction_2_i284;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u76_stall_local;
wire [31:0] local_bb4_var__u76;

assign local_bb4_var__u76[31:1] = 31'h0;
assign local_bb4_var__u76[0] = rnode_387to388_bb4_cmp68_i285_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i289_stall_local;
wire [31:0] local_bb4_shl_i289;

assign local_bb4_shl_i289 = ((local_bb4_and74_i288 & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4__40_i295_valid_out;
wire local_bb4__40_i295_stall_in;
wire local_bb4__40_i295_inputs_ready;
wire local_bb4__40_i295_stall_local;
wire local_bb4__40_i295;

assign local_bb4__40_i295_inputs_ready = (rnode_386to387_bb4__33_i276_0_valid_out_0_NO_SHIFT_REG & rnode_386to387_bb4__33_i276_0_valid_out_1_NO_SHIFT_REG & rnode_386to387_bb4_and83_i292_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40_i295 = (local_bb4_cmp77_i291 | local_bb4__39_i294);
assign local_bb4__40_i295_valid_out = 1'b1;
assign rnode_386to387_bb4__33_i276_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb4__33_i276_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb4_and83_i292_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or76_i290_valid_out;
wire local_bb4_or76_i290_stall_in;
wire local_bb4_or76_i290_inputs_ready;
wire local_bb4_or76_i290_stall_local;
wire [31:0] local_bb4_or76_i290;

assign local_bb4_or76_i290_inputs_ready = (rnode_386to387_bb4__37_i280_0_valid_out_1_NO_SHIFT_REG & rnode_386to387_bb4_and75_i286_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or76_i290 = ((local_bb4_shl_i289 & 32'h7F800000) | (rnode_386to387_bb4_and75_i286_0_NO_SHIFT_REG & 32'h7FFFFF));
assign local_bb4_or76_i290_valid_out = 1'b1;
assign rnode_386to387_bb4__37_i280_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_386to387_bb4_and75_i286_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4__40_i295_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4__40_i295_0_stall_in_NO_SHIFT_REG;
 logic rnode_387to388_bb4__40_i295_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4__40_i295_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic rnode_387to388_bb4__40_i295_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4__40_i295_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4__40_i295_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4__40_i295_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4__40_i295_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4__40_i295_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4__40_i295_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4__40_i295_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4__40_i295_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in(local_bb4__40_i295),
	.data_out(rnode_387to388_bb4__40_i295_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4__40_i295_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4__40_i295_0_reg_388_fifo.DATA_WIDTH = 1;
defparam rnode_387to388_bb4__40_i295_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4__40_i295_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4__40_i295_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_i295_stall_in = 1'b0;
assign rnode_387to388_bb4__40_i295_0_NO_SHIFT_REG = rnode_387to388_bb4__40_i295_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4__40_i295_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4__40_i295_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_387to388_bb4_or76_i290_0_valid_out_NO_SHIFT_REG;
 logic rnode_387to388_bb4_or76_i290_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_or76_i290_0_NO_SHIFT_REG;
 logic rnode_387to388_bb4_or76_i290_0_reg_388_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_387to388_bb4_or76_i290_0_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_or76_i290_0_valid_out_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_or76_i290_0_stall_in_reg_388_NO_SHIFT_REG;
 logic rnode_387to388_bb4_or76_i290_0_stall_out_reg_388_NO_SHIFT_REG;

acl_data_fifo rnode_387to388_bb4_or76_i290_0_reg_388_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_387to388_bb4_or76_i290_0_reg_388_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_387to388_bb4_or76_i290_0_stall_in_reg_388_NO_SHIFT_REG),
	.valid_out(rnode_387to388_bb4_or76_i290_0_valid_out_reg_388_NO_SHIFT_REG),
	.stall_out(rnode_387to388_bb4_or76_i290_0_stall_out_reg_388_NO_SHIFT_REG),
	.data_in((local_bb4_or76_i290 & 32'h7FFFFFFF)),
	.data_out(rnode_387to388_bb4_or76_i290_0_reg_388_NO_SHIFT_REG)
);

defparam rnode_387to388_bb4_or76_i290_0_reg_388_fifo.DEPTH = 1;
defparam rnode_387to388_bb4_or76_i290_0_reg_388_fifo.DATA_WIDTH = 32;
defparam rnode_387to388_bb4_or76_i290_0_reg_388_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_387to388_bb4_or76_i290_0_reg_388_fifo.IMPL = "shift_reg";

assign rnode_387to388_bb4_or76_i290_0_reg_388_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or76_i290_stall_in = 1'b0;
assign rnode_387to388_bb4_or76_i290_0_NO_SHIFT_REG = rnode_387to388_bb4_or76_i290_0_reg_388_NO_SHIFT_REG;
assign rnode_387to388_bb4_or76_i290_0_stall_in_reg_388_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_or76_i290_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cond_i296_stall_local;
wire [31:0] local_bb4_cond_i296;

assign local_bb4_cond_i296[31:1] = 31'h0;
assign local_bb4_cond_i296[0] = rnode_387to388_bb4__40_i295_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add87_i297_stall_local;
wire [31:0] local_bb4_add87_i297;

assign local_bb4_add87_i297 = ((local_bb4_cond_i296 & 32'h1) + (rnode_387to388_bb4_or76_i290_0_NO_SHIFT_REG & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i298_stall_local;
wire [31:0] local_bb4_and88_i298;

assign local_bb4_and88_i298 = (local_bb4_add87_i297 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i300_stall_local;
wire [31:0] local_bb4_and90_i300;

assign local_bb4_and90_i300 = (local_bb4_add87_i297 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_or89_i299_stall_local;
wire [31:0] local_bb4_or89_i299;

assign local_bb4_or89_i299 = ((local_bb4_and88_i298 & 32'h7FFFFFFF) | (local_bb4_and4_i225 & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i301_stall_local;
wire local_bb4_cmp91_i301;

assign local_bb4_cmp91_i301 = ((local_bb4_and90_i300 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge14_i303_stall_local;
wire local_bb4_brmerge14_i303;

assign local_bb4_brmerge14_i303 = (local_bb4_cmp91_i301 | rnode_387to388_bb4_cmp71_not_i302_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_conv99_i304_stall_local;
wire [31:0] local_bb4_conv99_i304;

assign local_bb4_conv99_i304 = (local_bb4_brmerge14_i303 ? (local_bb4_var__u76 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or102_i306_stall_local;
wire [31:0] local_bb4_or102_i306;

assign local_bb4_or102_i306 = ((local_bb4_conv99_i304 & 32'h1) | (local_bb4_conv101_i305 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool103_i307_stall_local;
wire local_bb4_tobool103_i307;

assign local_bb4_tobool103_i307 = ((local_bb4_or102_i306 & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cond107_i308_stall_local;
wire [31:0] local_bb4_cond107_i308;

assign local_bb4_cond107_i308 = (local_bb4_tobool103_i307 ? (local_bb4_and4_i225 & 32'h80000000) : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and108_i309_stall_local;
wire [31:0] local_bb4_and108_i309;

assign local_bb4_and108_i309 = (local_bb4_cond107_i308 & local_bb4_or89_i299);

// This section implements an unregistered operation.
// 
wire local_bb4_or112_i311_stall_local;
wire [31:0] local_bb4_or112_i311;

assign local_bb4_or112_i311 = (local_bb4_and108_i309 | (local_bb4_cond111_i310 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u77_stall_local;
wire [31:0] local_bb4_var__u77;

assign local_bb4_var__u77 = local_bb4_or112_i311;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u78_stall_local;
wire [31:0] local_bb4_var__u78;

assign local_bb4_var__u78 = (rnode_387to388_bb4__29_i253_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb4_var__u77);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u79_stall_local;
wire [31:0] local_bb4_var__u79;

assign local_bb4_var__u79 = local_bb4_var__u78;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i193_stall_local;
wire [31:0] local_bb4_shr_i193;

assign local_bb4_shr_i193 = (local_bb4_var__u79 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i195_stall_local;
wire [31:0] local_bb4_xor_i195;

assign local_bb4_xor_i195 = (local_bb4_var__u39 ^ local_bb4_var__u79);

// This section implements an unregistered operation.
// 
wire local_bb4_and5_i_stall_local;
wire [31:0] local_bb4_and5_i;

assign local_bb4_and5_i = (local_bb4_var__u79 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i205_stall_local;
wire [31:0] local_bb4_or_i205;

assign local_bb4_or_i205 = ((local_bb4_and5_i & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i_valid_out;
wire local_bb4_shr2_i_stall_in;
wire local_bb4_xor_i195_valid_out;
wire local_bb4_xor_i195_stall_in;
wire local_bb4_and6_i_valid_out_1;
wire local_bb4_and6_i_stall_in_1;
wire local_bb4_conv1_i_i_valid_out;
wire local_bb4_conv1_i_i_stall_in;
wire local_bb4_var__u78_valid_out_1;
wire local_bb4_var__u78_stall_in_1;
wire local_bb4_shr_i193_valid_out;
wire local_bb4_shr_i193_stall_in;
wire local_bb4_and5_i_valid_out_1;
wire local_bb4_and5_i_stall_in_1;
wire local_bb4_conv_i_i_valid_out;
wire local_bb4_conv_i_i_stall_in;
wire local_bb4_conv_i_i_inputs_ready;
wire local_bb4_conv_i_i_stall_local;
wire [63:0] local_bb4_conv_i_i;

assign local_bb4_conv_i_i_inputs_ready = (rnode_387to388_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb4_xor_i224_0_valid_out_NO_SHIFT_REG & rnode_386to388_bb4_or581_i282_0_valid_out_1_NO_SHIFT_REG & rnode_387to388_bb4__29_i253_0_valid_out_NO_SHIFT_REG & rnode_386to388_bb4_or581_i282_0_valid_out_0_NO_SHIFT_REG & rnode_387to388_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb4_cmp68_i285_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb4_cmp71_not_i302_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb4__40_i295_0_valid_out_NO_SHIFT_REG & rnode_387to388_bb4_or76_i290_0_valid_out_NO_SHIFT_REG);
assign local_bb4_conv_i_i[63:32] = 32'h0;
assign local_bb4_conv_i_i[31:0] = ((local_bb4_or_i205 & 32'hFFFFFF) | 32'h800000);
assign local_bb4_shr2_i_valid_out = 1'b1;
assign local_bb4_xor_i195_valid_out = 1'b1;
assign local_bb4_and6_i_valid_out_1 = 1'b1;
assign local_bb4_conv1_i_i_valid_out = 1'b1;
assign local_bb4_var__u78_valid_out_1 = 1'b1;
assign local_bb4_shr_i193_valid_out = 1'b1;
assign local_bb4_and5_i_valid_out_1 = 1'b1;
assign local_bb4_conv_i_i_valid_out = 1'b1;
assign rnode_387to388_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to388_bb4_or581_i282_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_386to388_bb4_or581_i282_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_cmp68_i285_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_cmp71_not_i302_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4__40_i295_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_387to388_bb4_or76_i290_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_shr2_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr2_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_shr2_i_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr2_i_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_shr2_i_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr2_i_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr2_i_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr2_i_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_shr2_i_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_shr2_i_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_shr2_i_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_shr2_i_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_shr2_i_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb4_shr2_i & 32'h1FF)),
	.data_out(rnode_388to389_bb4_shr2_i_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_shr2_i_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_shr2_i_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb4_shr2_i_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_shr2_i_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_shr2_i_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr2_i_stall_in = 1'b0;
assign rnode_388to389_bb4_shr2_i_0_NO_SHIFT_REG = rnode_388to389_bb4_shr2_i_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_shr2_i_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_shr2_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb4_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_xor_i195_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_xor_i195_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_xor_i195_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_xor_i195_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_xor_i195_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_xor_i195_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_xor_i195_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_xor_i195_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_xor_i195_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_xor_i195_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_xor_i195_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i195),
	.data_out(rnode_388to389_bb4_xor_i195_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_xor_i195_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_xor_i195_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb4_xor_i195_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_xor_i195_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_xor_i195_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i195_stall_in = 1'b0;
assign rnode_388to389_bb4_xor_i195_0_NO_SHIFT_REG = rnode_388to389_bb4_xor_i195_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_xor_i195_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_and6_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_and6_i_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_and6_i_1_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_and6_i_2_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_and6_i_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_valid_out_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_stall_in_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and6_i_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_and6_i_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_and6_i_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_and6_i_0_stall_in_0_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_and6_i_0_valid_out_0_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_and6_i_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb4_and6_i & 32'h7FFFFF)),
	.data_out(rnode_388to389_bb4_and6_i_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_and6_i_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_and6_i_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb4_and6_i_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_and6_i_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_and6_i_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and6_i_stall_in_1 = 1'b0;
assign rnode_388to389_bb4_and6_i_0_stall_in_0_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_and6_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_and6_i_0_NO_SHIFT_REG = rnode_388to389_bb4_and6_i_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_and6_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_and6_i_1_NO_SHIFT_REG = rnode_388to389_bb4_and6_i_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_and6_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_and6_i_2_NO_SHIFT_REG = rnode_388to389_bb4_and6_i_0_reg_389_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_var__u78_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb4_var__u78_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_var__u78_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_var__u78_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_var__u78_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_var__u78_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_var__u78_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_var__u78_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_var__u78_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_var__u78_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_var__u78_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_var__u78_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_var__u78_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in(local_bb4_var__u78),
	.data_out(rnode_388to389_bb4_var__u78_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_var__u78_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_var__u78_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb4_var__u78_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_var__u78_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_var__u78_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u78_stall_in_1 = 1'b0;
assign rnode_388to389_bb4_var__u78_0_NO_SHIFT_REG = rnode_388to389_bb4_var__u78_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_var__u78_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_var__u78_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_shr_i193_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr_i193_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_shr_i193_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr_i193_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_shr_i193_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr_i193_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr_i193_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_shr_i193_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_shr_i193_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_shr_i193_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_shr_i193_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_shr_i193_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_shr_i193_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb4_shr_i193 & 32'h1FF)),
	.data_out(rnode_388to389_bb4_shr_i193_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_shr_i193_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_shr_i193_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb4_shr_i193_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_shr_i193_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_shr_i193_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr_i193_stall_in = 1'b0;
assign rnode_388to389_bb4_shr_i193_0_NO_SHIFT_REG = rnode_388to389_bb4_shr_i193_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_shr_i193_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_shr_i193_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_388to389_bb4_and5_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and5_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_and5_i_0_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and5_i_0_reg_389_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_388to389_bb4_and5_i_0_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and5_i_0_valid_out_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and5_i_0_stall_in_reg_389_NO_SHIFT_REG;
 logic rnode_388to389_bb4_and5_i_0_stall_out_reg_389_NO_SHIFT_REG;

acl_data_fifo rnode_388to389_bb4_and5_i_0_reg_389_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_388to389_bb4_and5_i_0_reg_389_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_388to389_bb4_and5_i_0_stall_in_reg_389_NO_SHIFT_REG),
	.valid_out(rnode_388to389_bb4_and5_i_0_valid_out_reg_389_NO_SHIFT_REG),
	.stall_out(rnode_388to389_bb4_and5_i_0_stall_out_reg_389_NO_SHIFT_REG),
	.data_in((local_bb4_and5_i & 32'h7FFFFF)),
	.data_out(rnode_388to389_bb4_and5_i_0_reg_389_NO_SHIFT_REG)
);

defparam rnode_388to389_bb4_and5_i_0_reg_389_fifo.DEPTH = 1;
defparam rnode_388to389_bb4_and5_i_0_reg_389_fifo.DATA_WIDTH = 32;
defparam rnode_388to389_bb4_and5_i_0_reg_389_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_388to389_bb4_and5_i_0_reg_389_fifo.IMPL = "shift_reg";

assign rnode_388to389_bb4_and5_i_0_reg_389_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and5_i_stall_in_1 = 1'b0;
assign rnode_388to389_bb4_and5_i_0_NO_SHIFT_REG = rnode_388to389_bb4_and5_i_0_reg_389_NO_SHIFT_REG;
assign rnode_388to389_bb4_and5_i_0_stall_in_reg_389_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_and5_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_mul_i_i_inputs_ready;
 reg local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG;
wire local_bb4_mul_i_i_stall_in_0;
 reg local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i_stall_in_1;
wire local_bb4_mul_i_i_output_regs_ready;
wire [63:0] local_bb4_mul_i_i;
 reg local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul_i_i_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i_causedstall;

acl_int_mult int_module_local_bb4_mul_i_i (
	.clock(clock),
	.dataa(((local_bb4_conv1_i_i & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb4_conv_i_i & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb4_mul_i_i_output_regs_ready),
	.result(local_bb4_mul_i_i)
);

defparam int_module_local_bb4_mul_i_i.INPUT1_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i.INPUT2_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i.OUTPUT_WIDTH = 64;
defparam int_module_local_bb4_mul_i_i.LATENCY = 3;
defparam int_module_local_bb4_mul_i_i.SIGNED = 0;

assign local_bb4_mul_i_i_inputs_ready = 1'b1;
assign local_bb4_mul_i_i_output_regs_ready = 1'b1;
assign local_bb4_conv1_i_i_stall_in = 1'b0;
assign local_bb4_conv_i_i_stall_in = 1'b0;
assign local_bb4_mul_i_i_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i_output_regs_ready)
		begin
			local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i_output_regs_ready)
		begin
			local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul_i_i_stall_in_0))
			begin
				local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_mul_i_i_stall_in_1))
			begin
				local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and3_i_stall_local;
wire [31:0] local_bb4_and3_i;

assign local_bb4_and3_i = ((rnode_388to389_bb4_shr2_i_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_389to392_bb4_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to392_bb4_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_389to392_bb4_xor_i195_0_NO_SHIFT_REG;
 logic rnode_389to392_bb4_xor_i195_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to392_bb4_xor_i195_0_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb4_xor_i195_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb4_xor_i195_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_389to392_bb4_xor_i195_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_389to392_bb4_xor_i195_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to392_bb4_xor_i195_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to392_bb4_xor_i195_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_389to392_bb4_xor_i195_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_389to392_bb4_xor_i195_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_388to389_bb4_xor_i195_0_NO_SHIFT_REG),
	.data_out(rnode_389to392_bb4_xor_i195_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_389to392_bb4_xor_i195_0_reg_392_fifo.DEPTH = 3;
defparam rnode_389to392_bb4_xor_i195_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_389to392_bb4_xor_i195_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to392_bb4_xor_i195_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_389to392_bb4_xor_i195_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_388to389_bb4_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_389to392_bb4_xor_i195_0_NO_SHIFT_REG = rnode_389to392_bb4_xor_i195_0_reg_392_NO_SHIFT_REG;
assign rnode_389to392_bb4_xor_i195_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_389to392_bb4_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_i_stall_local;
wire local_bb4_lnot17_i;

assign local_bb4_lnot17_i = ((rnode_388to389_bb4_and6_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u80_stall_local;
wire [31:0] local_bb4_var__u80;

assign local_bb4_var__u80 = rnode_388to389_bb4_var__u78_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i194_stall_local;
wire [31:0] local_bb4_and_i194;

assign local_bb4_and_i194 = ((rnode_388to389_bb4_shr_i193_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i_stall_local;
wire local_bb4_lnot14_i;

assign local_bb4_lnot14_i = ((rnode_388to389_bb4_and5_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_conv3_i_i_stall_local;
wire [31:0] local_bb4_conv3_i_i;
wire [63:0] local_bb4_conv3_i_i$ps;

assign local_bb4_conv3_i_i$ps = (local_bb4_mul_i_i & 64'hFFFFFFFFFFFF);
assign local_bb4_conv3_i_i = local_bb4_conv3_i_i$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u81_stall_local;
wire [63:0] local_bb4_var__u81;

assign local_bb4_var__u81 = ((local_bb4_mul_i_i & 64'hFFFFFFFFFFFF) >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot8_i_stall_local;
wire local_bb4_lnot8_i;

assign local_bb4_lnot8_i = ((local_bb4_and3_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_i_stall_local;
wire local_bb4_cmp11_i;

assign local_bb4_cmp11_i = ((local_bb4_and3_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u82_stall_local;
wire [31:0] local_bb4_var__u82;

assign local_bb4_var__u82 = ((local_bb4_and3_i & 32'hFF) | (rnode_388to389_bb4_and6_i_1_NO_SHIFT_REG & 32'h7FFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_xor_i195_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_xor_i195_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_xor_i195_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_xor_i195_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_xor_i195_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_xor_i195_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_xor_i195_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_xor_i195_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_xor_i195_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_xor_i195_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_xor_i195_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_389to392_bb4_xor_i195_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb4_xor_i195_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_xor_i195_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_xor_i195_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_392to393_bb4_xor_i195_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_xor_i195_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_xor_i195_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to392_bb4_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_xor_i195_0_NO_SHIFT_REG = rnode_392to393_bb4_xor_i195_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_xor_i195_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_not_i_stall_local;
wire local_bb4_lnot17_not_i;

assign local_bb4_lnot17_not_i = (local_bb4_lnot17_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_stall_local;
wire [31:0] local_bb4_and_i;

assign local_bb4_and_i = (local_bb4_var__u80 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i_stall_local;
wire [31:0] local_bb4_and10_i;

assign local_bb4_and10_i = (local_bb4_var__u80 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i196_stall_local;
wire local_bb4_lnot_i196;

assign local_bb4_lnot_i196 = ((local_bb4_and_i194 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i197_stall_local;
wire local_bb4_cmp_i197;

assign local_bb4_cmp_i197 = ((local_bb4_and_i194 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u83_stall_local;
wire [31:0] local_bb4_var__u83;

assign local_bb4_var__u83 = ((rnode_388to389_bb4_and6_i_2_NO_SHIFT_REG & 32'h7FFFFF) | (local_bb4_and_i194 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i206_stall_local;
wire [31:0] local_bb4_add_i206;

assign local_bb4_add_i206 = ((local_bb4_and3_i & 32'hFF) + (local_bb4_and_i194 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_not_i_stall_local;
wire local_bb4_lnot14_not_i;

assign local_bb4_lnot14_not_i = (local_bb4_lnot14_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i16_i_stall_local;
wire [31:0] local_bb4_shr_i16_i;

assign local_bb4_shr_i16_i = (local_bb4_conv3_i_i >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i18_i_stall_local;
wire [31:0] local_bb4_shl1_i18_i;

assign local_bb4_shl1_i18_i = (local_bb4_conv3_i_i << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u84_stall_local;
wire [31:0] local_bb4_var__u84;

assign local_bb4_var__u84 = (local_bb4_conv3_i_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i_i_stall_local;
wire [31:0] local_bb4_shl1_i_i;

assign local_bb4_shl1_i_i = (local_bb4_conv3_i_i << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb4__tr_i_stall_local;
wire [31:0] local_bb4__tr_i;
wire [63:0] local_bb4__tr_i$ps;

assign local_bb4__tr_i$ps = (local_bb4_var__u81 & 64'hFFFFFF);
assign local_bb4__tr_i = local_bb4__tr_i$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge8_demorgan_i_stall_local;
wire local_bb4_brmerge8_demorgan_i;

assign local_bb4_brmerge8_demorgan_i = (local_bb4_cmp11_i & local_bb4_lnot17_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_not_i_stall_local;
wire local_bb4_cmp11_not_i;

assign local_bb4_cmp11_not_i = (local_bb4_cmp11_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u85_stall_local;
wire local_bb4_var__u85;

assign local_bb4_var__u85 = ((local_bb4_var__u82 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and4_i_stall_local;
wire [31:0] local_bb4_and4_i;

assign local_bb4_and4_i = (rnode_392to393_bb4_xor_i195_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i1_stall_local;
wire [31:0] local_bb4_shr_i1;

assign local_bb4_shr_i1 = ((local_bb4_and_i & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i_stall_local;
wire local_bb4_cmp13_i;

assign local_bb4_cmp13_i = ((local_bb4_and10_i & 32'hFFFF) > (local_bb4_and12_i & 32'hFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i212_stall_local;
wire local_bb4_reduction_0_i212;

assign local_bb4_reduction_0_i212 = (local_bb4_lnot_i196 | local_bb4_lnot8_i);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u86_stall_local;
wire local_bb4_var__u86;

assign local_bb4_var__u86 = (local_bb4_cmp_i197 | local_bb4_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u87_stall_local;
wire local_bb4_var__u87;

assign local_bb4_var__u87 = ((local_bb4_var__u83 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i203_stall_local;
wire local_bb4__28_i203;

assign local_bb4__28_i203 = (local_bb4_cmp_i197 & local_bb4_lnot14_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i207_stall_local;
wire [31:0] local_bb4_shr_i_i207;

assign local_bb4_shr_i_i207 = ((local_bb4_var__u84 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i15_i_stall_local;
wire [31:0] local_bb4_shl_i15_i;

assign local_bb4_shl_i15_i = ((local_bb4__tr_i & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb4_and48_i_stall_local;
wire [31:0] local_bb4_and48_i;

assign local_bb4_and48_i = ((local_bb4__tr_i & 32'hFFFFFF) & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge10_demorgan_i_stall_local;
wire local_bb4_brmerge10_demorgan_i;

assign local_bb4_brmerge10_demorgan_i = (local_bb4_brmerge8_demorgan_i & local_bb4_lnot_i196);

// This section implements an unregistered operation.
// 
wire local_bb4__mux9_mux_i_stall_local;
wire local_bb4__mux9_mux_i;

assign local_bb4__mux9_mux_i = (local_bb4_brmerge8_demorgan_i ^ local_bb4_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge3_i_stall_local;
wire local_bb4_brmerge3_i;

assign local_bb4_brmerge3_i = (local_bb4_var__u85 | local_bb4_cmp11_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_i_stall_local;
wire local_bb4__mux_mux_i;

assign local_bb4__mux_mux_i = (local_bb4_var__u85 | local_bb4_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb4__not_i_stall_local;
wire local_bb4__not_i;

assign local_bb4__not_i = (local_bb4_var__u85 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i3_stall_local;
wire local_bb4_cmp_i3;

assign local_bb4_cmp_i3 = ((local_bb4_shr_i1 & 32'h7FFF) > (local_bb4_shr3_i & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i_stall_local;
wire local_bb4_cmp8_i;

assign local_bb4_cmp8_i = ((local_bb4_shr_i1 & 32'h7FFF) == (local_bb4_shr3_i & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_or_i17_i_stall_local;
wire [31:0] local_bb4_or_i17_i;

assign local_bb4_or_i17_i = ((local_bb4_shl_i15_i & 32'hFFFF00) | (local_bb4_shr_i16_i & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool49_i_stall_local;
wire local_bb4_tobool49_i;

assign local_bb4_tobool49_i = ((local_bb4_and48_i & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__26_demorgan_i_stall_local;
wire local_bb4__26_demorgan_i;

assign local_bb4__26_demorgan_i = (local_bb4_cmp_i197 | local_bb4_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge5_i_stall_local;
wire local_bb4_brmerge5_i;

assign local_bb4_brmerge5_i = (local_bb4_brmerge3_i | local_bb4_lnot17_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i198_stall_local;
wire local_bb4_reduction_3_i198;

assign local_bb4_reduction_3_i198 = (local_bb4_cmp11_i & local_bb4__not_i);

// This section implements an unregistered operation.
// 
wire local_bb4___i4_stall_local;
wire local_bb4___i4;

assign local_bb4___i4 = (local_bb4_cmp8_i & local_bb4_cmp13_i);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_i_stall_local;
wire [31:0] local_bb4_shl_i_i;

assign local_bb4_shl_i_i = ((local_bb4_or_i17_i & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_mux_i_stall_local;
wire local_bb4__mux_mux_mux_i;

assign local_bb4__mux_mux_mux_i = (local_bb4_brmerge5_i & local_bb4__mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i199_stall_local;
wire local_bb4_reduction_5_i199;

assign local_bb4_reduction_5_i199 = (local_bb4_lnot14_i & local_bb4_reduction_3_i198);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u52_valid_out_2;
wire local_bb4_var__u52_stall_in_2;
wire local_bb4__21_i_valid_out;
wire local_bb4__21_i_stall_in;
wire local_bb4_var__u80_valid_out_2;
wire local_bb4_var__u80_stall_in_2;
wire local_bb4__21_i_inputs_ready;
wire local_bb4__21_i_stall_local;
wire local_bb4__21_i;

assign local_bb4__21_i_inputs_ready = (rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_valid_out_0_NO_SHIFT_REG & rnode_388to389_bb4_var__u78_0_valid_out_NO_SHIFT_REG);
assign local_bb4__21_i = (local_bb4_cmp_i3 | local_bb4___i4);
assign local_bb4_var__u52_valid_out_2 = 1'b1;
assign local_bb4__21_i_valid_out = 1'b1;
assign local_bb4_var__u80_valid_out_2 = 1'b1;
assign rnode_388to389_bb4_sum_312_pop9_c1_ene6_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_var__u78_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i208_stall_local;
wire [31:0] local_bb4_or_i_i208;

assign local_bb4_or_i_i208 = ((local_bb4_shl_i_i & 32'h1FFFFFE) | (local_bb4_shr_i_i207 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i200_stall_local;
wire local_bb4_reduction_6_i200;

assign local_bb4_reduction_6_i200 = (local_bb4_var__u87 & local_bb4_reduction_5_i199);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb4_var__u52_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u52_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_var__u52_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u52_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u52_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_var__u52_1_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u52_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_var__u52_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u52_0_valid_out_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u52_0_stall_in_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u52_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb4_var__u52_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb4_var__u52_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb4_var__u52_0_stall_in_0_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb4_var__u52_0_valid_out_0_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb4_var__u52_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb4_var__u52),
	.data_out(rnode_389to390_bb4_var__u52_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb4_var__u52_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb4_var__u52_0_reg_390_fifo.DATA_WIDTH = 32;
defparam rnode_389to390_bb4_var__u52_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb4_var__u52_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb4_var__u52_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u52_stall_in_2 = 1'b0;
assign rnode_389to390_bb4_var__u52_0_stall_in_0_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_var__u52_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4_var__u52_0_NO_SHIFT_REG = rnode_389to390_bb4_var__u52_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb4_var__u52_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4_var__u52_1_NO_SHIFT_REG = rnode_389to390_bb4_var__u52_0_reg_390_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb4__21_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_1_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_valid_out_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_stall_in_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4__21_i_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb4__21_i_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb4__21_i_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb4__21_i_0_stall_in_0_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb4__21_i_0_valid_out_0_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb4__21_i_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb4__21_i),
	.data_out(rnode_389to390_bb4__21_i_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb4__21_i_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb4__21_i_0_reg_390_fifo.DATA_WIDTH = 1;
defparam rnode_389to390_bb4__21_i_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb4__21_i_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb4__21_i_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i_stall_in = 1'b0;
assign rnode_389to390_bb4__21_i_0_stall_in_0_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4__21_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4__21_i_0_NO_SHIFT_REG = rnode_389to390_bb4__21_i_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb4__21_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4__21_i_1_NO_SHIFT_REG = rnode_389to390_bb4__21_i_0_reg_390_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb4_var__u80_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u80_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_var__u80_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u80_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u80_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_var__u80_1_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u80_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to390_bb4_var__u80_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u80_0_valid_out_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u80_0_stall_in_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u80_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb4_var__u80_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb4_var__u80_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb4_var__u80_0_stall_in_0_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb4_var__u80_0_valid_out_0_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb4_var__u80_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb4_var__u80),
	.data_out(rnode_389to390_bb4_var__u80_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb4_var__u80_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb4_var__u80_0_reg_390_fifo.DATA_WIDTH = 32;
defparam rnode_389to390_bb4_var__u80_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb4_var__u80_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb4_var__u80_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u80_stall_in_2 = 1'b0;
assign rnode_389to390_bb4_var__u80_0_stall_in_0_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_var__u80_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4_var__u80_0_NO_SHIFT_REG = rnode_389to390_bb4_var__u80_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb4_var__u80_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4_var__u80_1_NO_SHIFT_REG = rnode_389to390_bb4_var__u80_0_reg_390_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__24_i201_stall_local;
wire local_bb4__24_i201;

assign local_bb4__24_i201 = (local_bb4_cmp_i197 ? local_bb4_reduction_6_i200 : local_bb4_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i_stall_local;
wire [31:0] local_bb4__22_i;

assign local_bb4__22_i = (rnode_389to390_bb4__21_i_0_NO_SHIFT_REG ? rnode_389to390_bb4_var__u52_0_NO_SHIFT_REG : rnode_389to390_bb4_var__u80_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i_stall_local;
wire [31:0] local_bb4__23_i;

assign local_bb4__23_i = (rnode_389to390_bb4__21_i_1_NO_SHIFT_REG ? rnode_389to390_bb4_var__u80_1_NO_SHIFT_REG : rnode_389to390_bb4_var__u52_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__25_i_stall_local;
wire local_bb4__25_i;

assign local_bb4__25_i = (local_bb4__24_i201 ? local_bb4_lnot14_i : local_bb4__mux_mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i_stall_local;
wire [31:0] local_bb4_shr18_i;

assign local_bb4_shr18_i = (local_bb4__22_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i_stall_local;
wire [31:0] local_bb4_shr16_i;

assign local_bb4_shr16_i = (local_bb4__23_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i202_stall_local;
wire local_bb4__27_i202;

assign local_bb4__27_i202 = (local_bb4__26_demorgan_i ? local_bb4__25_i : local_bb4__mux9_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i_stall_local;
wire [31:0] local_bb4_and19_i;

assign local_bb4_and19_i = ((local_bb4_shr18_i & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i_stall_local;
wire [31:0] local_bb4_sub_i;

assign local_bb4_sub_i = ((local_bb4_shr16_i & 32'h1FF) - (local_bb4_shr18_i & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i206_valid_out;
wire local_bb4_add_i206_stall_in;
wire local_bb4_reduction_0_i212_valid_out;
wire local_bb4_reduction_0_i212_stall_in;
wire local_bb4_var__u86_valid_out;
wire local_bb4_var__u86_stall_in;
wire local_bb4__29_i204_valid_out;
wire local_bb4__29_i204_stall_in;
wire local_bb4__29_i204_inputs_ready;
wire local_bb4__29_i204_stall_local;
wire local_bb4__29_i204;

assign local_bb4__29_i204_inputs_ready = (rnode_388to389_bb4_shr2_i_0_valid_out_NO_SHIFT_REG & rnode_388to389_bb4_and6_i_0_valid_out_1_NO_SHIFT_REG & rnode_388to389_bb4_and6_i_0_valid_out_0_NO_SHIFT_REG & rnode_388to389_bb4_and6_i_0_valid_out_2_NO_SHIFT_REG & rnode_388to389_bb4_shr_i193_0_valid_out_NO_SHIFT_REG & rnode_388to389_bb4_and5_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4__29_i204 = (local_bb4__28_i203 | local_bb4__27_i202);
assign local_bb4_add_i206_valid_out = 1'b1;
assign local_bb4_reduction_0_i212_valid_out = 1'b1;
assign local_bb4_var__u86_valid_out = 1'b1;
assign local_bb4__29_i204_valid_out = 1'b1;
assign rnode_388to389_bb4_shr2_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_and6_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_and6_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_and6_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_shr_i193_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_388to389_bb4_and5_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i_stall_local;
wire local_bb4_lnot23_i;

assign local_bb4_lnot23_i = ((local_bb4_and19_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i_stall_local;
wire local_bb4_cmp27_i;

assign local_bb4_cmp27_i = ((local_bb4_and19_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and68_i_stall_local;
wire [31:0] local_bb4_and68_i;

assign local_bb4_and68_i = (local_bb4_sub_i & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_389to391_bb4_add_i206_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb4_add_i206_0_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb4_add_i206_1_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb4_add_i206_2_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_389to391_bb4_add_i206_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_valid_out_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_stall_in_0_reg_391_NO_SHIFT_REG;
 logic rnode_389to391_bb4_add_i206_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_389to391_bb4_add_i206_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to391_bb4_add_i206_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to391_bb4_add_i206_0_stall_in_0_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_389to391_bb4_add_i206_0_valid_out_0_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_389to391_bb4_add_i206_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb4_add_i206 & 32'h1FF)),
	.data_out(rnode_389to391_bb4_add_i206_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_389to391_bb4_add_i206_0_reg_391_fifo.DEPTH = 2;
defparam rnode_389to391_bb4_add_i206_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_389to391_bb4_add_i206_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to391_bb4_add_i206_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_389to391_bb4_add_i206_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add_i206_stall_in = 1'b0;
assign rnode_389to391_bb4_add_i206_0_stall_in_0_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb4_add_i206_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_389to391_bb4_add_i206_0_NO_SHIFT_REG = rnode_389to391_bb4_add_i206_0_reg_391_NO_SHIFT_REG;
assign rnode_389to391_bb4_add_i206_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_389to391_bb4_add_i206_1_NO_SHIFT_REG = rnode_389to391_bb4_add_i206_0_reg_391_NO_SHIFT_REG;
assign rnode_389to391_bb4_add_i206_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_389to391_bb4_add_i206_2_NO_SHIFT_REG = rnode_389to391_bb4_add_i206_0_reg_391_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to390_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_389to390_bb4_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4_reduction_0_i212_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to390_bb4_reduction_0_i212_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_reduction_0_i212_0_valid_out_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_reduction_0_i212_0_stall_in_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_reduction_0_i212_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb4_reduction_0_i212_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb4_reduction_0_i212_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb4_reduction_0_i212_0_stall_in_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb4_reduction_0_i212_0_valid_out_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb4_reduction_0_i212_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_0_i212),
	.data_out(rnode_389to390_bb4_reduction_0_i212_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb4_reduction_0_i212_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb4_reduction_0_i212_0_reg_390_fifo.DATA_WIDTH = 1;
defparam rnode_389to390_bb4_reduction_0_i212_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb4_reduction_0_i212_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb4_reduction_0_i212_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_0_i212_stall_in = 1'b0;
assign rnode_389to390_bb4_reduction_0_i212_0_NO_SHIFT_REG = rnode_389to390_bb4_reduction_0_i212_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb4_reduction_0_i212_0_stall_in_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb4_var__u86_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u86_0_stall_in_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u86_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u86_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u86_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u86_0_valid_out_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u86_0_stall_in_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4_var__u86_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb4_var__u86_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb4_var__u86_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb4_var__u86_0_stall_in_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb4_var__u86_0_valid_out_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb4_var__u86_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb4_var__u86),
	.data_out(rnode_389to390_bb4_var__u86_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb4_var__u86_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb4_var__u86_0_reg_390_fifo.DATA_WIDTH = 1;
defparam rnode_389to390_bb4_var__u86_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb4_var__u86_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb4_var__u86_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u86_stall_in = 1'b0;
assign rnode_389to390_bb4_var__u86_0_NO_SHIFT_REG = rnode_389to390_bb4_var__u86_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb4_var__u86_0_stall_in_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_var__u86_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_389to390_bb4__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_389to390_bb4__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_389to390_bb4__29_i204_0_NO_SHIFT_REG;
 logic rnode_389to390_bb4__29_i204_0_reg_390_inputs_ready_NO_SHIFT_REG;
 logic rnode_389to390_bb4__29_i204_0_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4__29_i204_0_valid_out_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4__29_i204_0_stall_in_reg_390_NO_SHIFT_REG;
 logic rnode_389to390_bb4__29_i204_0_stall_out_reg_390_NO_SHIFT_REG;

acl_data_fifo rnode_389to390_bb4__29_i204_0_reg_390_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_389to390_bb4__29_i204_0_reg_390_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_389to390_bb4__29_i204_0_stall_in_reg_390_NO_SHIFT_REG),
	.valid_out(rnode_389to390_bb4__29_i204_0_valid_out_reg_390_NO_SHIFT_REG),
	.stall_out(rnode_389to390_bb4__29_i204_0_stall_out_reg_390_NO_SHIFT_REG),
	.data_in(local_bb4__29_i204),
	.data_out(rnode_389to390_bb4__29_i204_0_reg_390_NO_SHIFT_REG)
);

defparam rnode_389to390_bb4__29_i204_0_reg_390_fifo.DEPTH = 1;
defparam rnode_389to390_bb4__29_i204_0_reg_390_fifo.DATA_WIDTH = 1;
defparam rnode_389to390_bb4__29_i204_0_reg_390_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_389to390_bb4__29_i204_0_reg_390_fifo.IMPL = "shift_reg";

assign rnode_389to390_bb4__29_i204_0_reg_390_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__29_i204_stall_in = 1'b0;
assign rnode_389to390_bb4__29_i204_0_NO_SHIFT_REG = rnode_389to390_bb4__29_i204_0_reg_390_NO_SHIFT_REG;
assign rnode_389to390_bb4__29_i204_0_stall_in_reg_390_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp69_i_stall_local;
wire local_bb4_cmp69_i;

assign local_bb4_cmp69_i = ((local_bb4_and68_i & 32'hFF) > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_inc_i_stall_local;
wire [31:0] local_bb4_inc_i;

assign local_bb4_inc_i = ((rnode_389to391_bb4_add_i206_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp50_not_i_stall_local;
wire local_bb4_cmp50_not_i;

assign local_bb4_cmp50_not_i = ((rnode_389to391_bb4_add_i206_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_390to392_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to392_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_390to392_bb4_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_390to392_bb4_reduction_0_i212_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_390to392_bb4_reduction_0_i212_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_reduction_0_i212_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_reduction_0_i212_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_reduction_0_i212_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_390to392_bb4_reduction_0_i212_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to392_bb4_reduction_0_i212_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to392_bb4_reduction_0_i212_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_390to392_bb4_reduction_0_i212_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_390to392_bb4_reduction_0_i212_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_389to390_bb4_reduction_0_i212_0_NO_SHIFT_REG),
	.data_out(rnode_390to392_bb4_reduction_0_i212_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_390to392_bb4_reduction_0_i212_0_reg_392_fifo.DEPTH = 2;
defparam rnode_390to392_bb4_reduction_0_i212_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_390to392_bb4_reduction_0_i212_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to392_bb4_reduction_0_i212_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_390to392_bb4_reduction_0_i212_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4_reduction_0_i212_0_NO_SHIFT_REG = rnode_390to392_bb4_reduction_0_i212_0_reg_392_NO_SHIFT_REG;
assign rnode_390to392_bb4_reduction_0_i212_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4_var__u86_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb4_var__u86_0_stall_in_NO_SHIFT_REG;
 logic rnode_390to391_bb4_var__u86_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_var__u86_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic rnode_390to391_bb4_var__u86_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_var__u86_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_var__u86_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_var__u86_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4_var__u86_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4_var__u86_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4_var__u86_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4_var__u86_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4_var__u86_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in(rnode_389to390_bb4_var__u86_0_NO_SHIFT_REG),
	.data_out(rnode_390to391_bb4_var__u86_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4_var__u86_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4_var__u86_0_reg_391_fifo.DATA_WIDTH = 1;
defparam rnode_390to391_bb4_var__u86_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4_var__u86_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4_var__u86_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4_var__u86_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_var__u86_0_NO_SHIFT_REG = rnode_390to391_bb4_var__u86_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_var__u86_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_var__u86_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_390to392_bb4__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to392_bb4__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_390to392_bb4__29_i204_0_NO_SHIFT_REG;
 logic rnode_390to392_bb4__29_i204_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_390to392_bb4__29_i204_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4__29_i204_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4__29_i204_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4__29_i204_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_390to392_bb4__29_i204_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to392_bb4__29_i204_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to392_bb4__29_i204_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_390to392_bb4__29_i204_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_390to392_bb4__29_i204_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_389to390_bb4__29_i204_0_NO_SHIFT_REG),
	.data_out(rnode_390to392_bb4__29_i204_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_390to392_bb4__29_i204_0_reg_392_fifo.DEPTH = 2;
defparam rnode_390to392_bb4__29_i204_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_390to392_bb4__29_i204_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to392_bb4__29_i204_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_390to392_bb4__29_i204_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_389to390_bb4__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4__29_i204_0_NO_SHIFT_REG = rnode_390to392_bb4__29_i204_0_reg_392_NO_SHIFT_REG;
assign rnode_390to392_bb4__29_i204_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_align_0_i_stall_local;
wire [31:0] local_bb4_align_0_i;

assign local_bb4_align_0_i = (local_bb4_cmp69_i ? 32'h1F : (local_bb4_and68_i & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i209_stall_local;
wire local_bb4__31_i209;

assign local_bb4__31_i209 = (local_bb4_tobool49_i & local_bb4_cmp50_not_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_reduction_0_i212_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4_reduction_0_i212_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_reduction_0_i212_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_reduction_0_i212_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_reduction_0_i212_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_reduction_0_i212_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_reduction_0_i212_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_reduction_0_i212_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_reduction_0_i212_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_reduction_0_i212_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_390to392_bb4_reduction_0_i212_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb4_reduction_0_i212_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_reduction_0_i212_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_reduction_0_i212_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4_reduction_0_i212_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_reduction_0_i212_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_reduction_0_i212_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_reduction_0_i212_0_NO_SHIFT_REG = rnode_392to393_bb4_reduction_0_i212_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_reduction_0_i212_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_var__u86_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb4_var__u86_0_stall_in_NO_SHIFT_REG;
 logic rnode_391to392_bb4_var__u86_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_var__u86_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_391to392_bb4_var__u86_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_var__u86_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_var__u86_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_var__u86_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_var__u86_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_var__u86_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_var__u86_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_var__u86_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_var__u86_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(rnode_390to391_bb4_var__u86_0_NO_SHIFT_REG),
	.data_out(rnode_391to392_bb4_var__u86_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_var__u86_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_var__u86_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_391to392_bb4_var__u86_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_var__u86_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_var__u86_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4_var__u86_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_var__u86_0_NO_SHIFT_REG = rnode_391to392_bb4_var__u86_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_var__u86_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_var__u86_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4__29_i204_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4__29_i204_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4__29_i204_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__29_i204_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__29_i204_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__29_i204_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4__29_i204_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4__29_i204_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4__29_i204_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4__29_i204_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4__29_i204_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(rnode_390to392_bb4__29_i204_0_NO_SHIFT_REG),
	.data_out(rnode_392to393_bb4__29_i204_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4__29_i204_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4__29_i204_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4__29_i204_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4__29_i204_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4__29_i204_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4__29_i204_0_NO_SHIFT_REG = rnode_392to393_bb4__29_i204_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4__29_i204_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and93_i_stall_local;
wire [31:0] local_bb4_and93_i;

assign local_bb4_and93_i = ((local_bb4_align_0_i & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and95_i_stall_local;
wire [31:0] local_bb4_and95_i;

assign local_bb4_and95_i = ((local_bb4_align_0_i & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and115_i_stall_local;
wire [31:0] local_bb4_and115_i;

assign local_bb4_and115_i = ((local_bb4_align_0_i & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and130_i_stall_local;
wire [31:0] local_bb4_and130_i;

assign local_bb4_and130_i = ((local_bb4_align_0_i & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i_valid_out_1;
wire local_bb4__22_i_stall_in_1;
wire local_bb4__23_i_valid_out_1;
wire local_bb4__23_i_stall_in_1;
wire local_bb4_shr16_i_valid_out_1;
wire local_bb4_shr16_i_stall_in_1;
wire local_bb4_lnot23_i_valid_out;
wire local_bb4_lnot23_i_stall_in;
wire local_bb4_cmp27_i_valid_out;
wire local_bb4_cmp27_i_stall_in;
wire local_bb4_and93_i_valid_out;
wire local_bb4_and93_i_stall_in;
wire local_bb4_and95_i_valid_out;
wire local_bb4_and95_i_stall_in;
wire local_bb4_and115_i_valid_out;
wire local_bb4_and115_i_stall_in;
wire local_bb4_and130_i_valid_out;
wire local_bb4_and130_i_stall_in;
wire local_bb4_and149_i_valid_out;
wire local_bb4_and149_i_stall_in;
wire local_bb4_and149_i_inputs_ready;
wire local_bb4_and149_i_stall_local;
wire [31:0] local_bb4_and149_i;

assign local_bb4_and149_i_inputs_ready = (rnode_389to390_bb4__21_i_0_valid_out_0_NO_SHIFT_REG & rnode_389to390_bb4_var__u52_0_valid_out_0_NO_SHIFT_REG & rnode_389to390_bb4_var__u80_0_valid_out_0_NO_SHIFT_REG & rnode_389to390_bb4__21_i_0_valid_out_1_NO_SHIFT_REG & rnode_389to390_bb4_var__u80_0_valid_out_1_NO_SHIFT_REG & rnode_389to390_bb4_var__u52_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_and149_i = ((local_bb4_align_0_i & 32'hFF) & 32'h3);
assign local_bb4__22_i_valid_out_1 = 1'b1;
assign local_bb4__23_i_valid_out_1 = 1'b1;
assign local_bb4_shr16_i_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i_valid_out = 1'b1;
assign local_bb4_cmp27_i_valid_out = 1'b1;
assign local_bb4_and93_i_valid_out = 1'b1;
assign local_bb4_and95_i_valid_out = 1'b1;
assign local_bb4_and115_i_valid_out = 1'b1;
assign local_bb4_and130_i_valid_out = 1'b1;
assign local_bb4_and149_i_valid_out = 1'b1;
assign rnode_389to390_bb4__21_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_var__u52_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_var__u80_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4__21_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_var__u80_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_389to390_bb4_var__u52_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__32_i210_stall_local;
wire [31:0] local_bb4__32_i210;

assign local_bb4__32_i210 = (local_bb4__31_i209 ? (local_bb4_shl1_i_i & 32'hFFFFFE00) : (local_bb4_shl1_i18_i & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__34_i_stall_local;
wire [31:0] local_bb4__34_i;

assign local_bb4__34_i = (local_bb4__31_i209 ? (local_bb4_or_i_i208 & 32'h1FFFFFF) : (local_bb4_or_i17_i & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__36_i_stall_local;
wire [31:0] local_bb4__36_i;

assign local_bb4__36_i = (local_bb4__31_i209 ? (rnode_389to391_bb4_add_i206_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4__22_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4__22_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4__22_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4__22_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_390to391_bb4__22_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4__22_i_1_NO_SHIFT_REG;
 logic rnode_390to391_bb4__22_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4__22_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4__22_i_0_valid_out_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4__22_i_0_stall_in_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4__22_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4__22_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4__22_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4__22_i_0_stall_in_0_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4__22_i_0_valid_out_0_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4__22_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in(local_bb4__22_i),
	.data_out(rnode_390to391_bb4__22_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4__22_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4__22_i_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb4__22_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4__22_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4__22_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i_stall_in_1 = 1'b0;
assign rnode_390to391_bb4__22_i_0_stall_in_0_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4__22_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4__22_i_0_NO_SHIFT_REG = rnode_390to391_bb4__22_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4__22_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4__22_i_1_NO_SHIFT_REG = rnode_390to391_bb4__22_i_0_reg_391_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4__23_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4__23_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4__23_i_1_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4__23_i_2_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4__23_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_valid_out_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_stall_in_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4__23_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4__23_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4__23_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4__23_i_0_stall_in_0_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4__23_i_0_valid_out_0_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4__23_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in(local_bb4__23_i),
	.data_out(rnode_390to391_bb4__23_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4__23_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4__23_i_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb4__23_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4__23_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4__23_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i_stall_in_1 = 1'b0;
assign rnode_390to391_bb4__23_i_0_stall_in_0_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4__23_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4__23_i_0_NO_SHIFT_REG = rnode_390to391_bb4__23_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4__23_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4__23_i_1_NO_SHIFT_REG = rnode_390to391_bb4__23_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4__23_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4__23_i_2_NO_SHIFT_REG = rnode_390to391_bb4__23_i_0_reg_391_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_390to392_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_390to392_bb4_shr16_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_390to392_bb4_shr16_i_0_NO_SHIFT_REG;
 logic rnode_390to392_bb4_shr16_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_390to392_bb4_shr16_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_390to392_bb4_shr16_i_1_NO_SHIFT_REG;
 logic rnode_390to392_bb4_shr16_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to392_bb4_shr16_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_shr16_i_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_shr16_i_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_shr16_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_390to392_bb4_shr16_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to392_bb4_shr16_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to392_bb4_shr16_i_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_390to392_bb4_shr16_i_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_390to392_bb4_shr16_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i & 32'h1FF)),
	.data_out(rnode_390to392_bb4_shr16_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_390to392_bb4_shr16_i_0_reg_392_fifo.DEPTH = 2;
defparam rnode_390to392_bb4_shr16_i_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_390to392_bb4_shr16_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to392_bb4_shr16_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_390to392_bb4_shr16_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i_stall_in_1 = 1'b0;
assign rnode_390to392_bb4_shr16_i_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4_shr16_i_0_NO_SHIFT_REG = rnode_390to392_bb4_shr16_i_0_reg_392_NO_SHIFT_REG;
assign rnode_390to392_bb4_shr16_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4_shr16_i_1_NO_SHIFT_REG = rnode_390to392_bb4_shr16_i_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb4_lnot23_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_390to391_bb4_lnot23_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_lnot23_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic rnode_390to391_bb4_lnot23_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_lnot23_i_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_lnot23_i_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_lnot23_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4_lnot23_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4_lnot23_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4_lnot23_i_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4_lnot23_i_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4_lnot23_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i),
	.data_out(rnode_390to391_bb4_lnot23_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4_lnot23_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4_lnot23_i_0_reg_391_fifo.DATA_WIDTH = 1;
defparam rnode_390to391_bb4_lnot23_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4_lnot23_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4_lnot23_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i_stall_in = 1'b0;
assign rnode_390to391_bb4_lnot23_i_0_NO_SHIFT_REG = rnode_390to391_bb4_lnot23_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_lnot23_i_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_390to392_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_1_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_2_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_390to392_bb4_cmp27_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_390to392_bb4_cmp27_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to392_bb4_cmp27_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to392_bb4_cmp27_i_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_390to392_bb4_cmp27_i_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_390to392_bb4_cmp27_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i),
	.data_out(rnode_390to392_bb4_cmp27_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_390to392_bb4_cmp27_i_0_reg_392_fifo.DEPTH = 2;
defparam rnode_390to392_bb4_cmp27_i_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_390to392_bb4_cmp27_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to392_bb4_cmp27_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_390to392_bb4_cmp27_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i_stall_in = 1'b0;
assign rnode_390to392_bb4_cmp27_i_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4_cmp27_i_0_NO_SHIFT_REG = rnode_390to392_bb4_cmp27_i_0_reg_392_NO_SHIFT_REG;
assign rnode_390to392_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4_cmp27_i_1_NO_SHIFT_REG = rnode_390to392_bb4_cmp27_i_0_reg_392_NO_SHIFT_REG;
assign rnode_390to392_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4_cmp27_i_2_NO_SHIFT_REG = rnode_390to392_bb4_cmp27_i_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4_and93_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and93_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and93_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and93_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and93_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and93_i_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and93_i_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and93_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4_and93_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4_and93_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4_and93_i_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4_and93_i_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4_and93_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb4_and93_i & 32'h1C)),
	.data_out(rnode_390to391_bb4_and93_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4_and93_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4_and93_i_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb4_and93_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4_and93_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4_and93_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and93_i_stall_in = 1'b0;
assign rnode_390to391_bb4_and93_i_0_NO_SHIFT_REG = rnode_390to391_bb4_and93_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_and93_i_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and93_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4_and95_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and95_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and95_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and95_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and95_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and95_i_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and95_i_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and95_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4_and95_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4_and95_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4_and95_i_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4_and95_i_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4_and95_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb4_and95_i & 32'h10)),
	.data_out(rnode_390to391_bb4_and95_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4_and95_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4_and95_i_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb4_and95_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4_and95_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4_and95_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and95_i_stall_in = 1'b0;
assign rnode_390to391_bb4_and95_i_0_NO_SHIFT_REG = rnode_390to391_bb4_and95_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_and95_i_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and95_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4_and115_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and115_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and115_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and115_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and115_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and115_i_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and115_i_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and115_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4_and115_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4_and115_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4_and115_i_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4_and115_i_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4_and115_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb4_and115_i & 32'h8)),
	.data_out(rnode_390to391_bb4_and115_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4_and115_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4_and115_i_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb4_and115_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4_and115_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4_and115_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and115_i_stall_in = 1'b0;
assign rnode_390to391_bb4_and115_i_0_NO_SHIFT_REG = rnode_390to391_bb4_and115_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_and115_i_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and115_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4_and130_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and130_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and130_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and130_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and130_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and130_i_0_valid_out_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and130_i_0_stall_in_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and130_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4_and130_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4_and130_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4_and130_i_0_stall_in_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4_and130_i_0_valid_out_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4_and130_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb4_and130_i & 32'h4)),
	.data_out(rnode_390to391_bb4_and130_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4_and130_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4_and130_i_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb4_and130_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4_and130_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4_and130_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and130_i_stall_in = 1'b0;
assign rnode_390to391_bb4_and130_i_0_NO_SHIFT_REG = rnode_390to391_bb4_and130_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_and130_i_0_stall_in_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and130_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_390to391_bb4_and149_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and149_i_0_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and149_i_1_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and149_i_2_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_reg_391_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_390to391_bb4_and149_i_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_valid_out_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_stall_in_0_reg_391_NO_SHIFT_REG;
 logic rnode_390to391_bb4_and149_i_0_stall_out_reg_391_NO_SHIFT_REG;

acl_data_fifo rnode_390to391_bb4_and149_i_0_reg_391_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_390to391_bb4_and149_i_0_reg_391_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_390to391_bb4_and149_i_0_stall_in_0_reg_391_NO_SHIFT_REG),
	.valid_out(rnode_390to391_bb4_and149_i_0_valid_out_0_reg_391_NO_SHIFT_REG),
	.stall_out(rnode_390to391_bb4_and149_i_0_stall_out_reg_391_NO_SHIFT_REG),
	.data_in((local_bb4_and149_i & 32'h3)),
	.data_out(rnode_390to391_bb4_and149_i_0_reg_391_NO_SHIFT_REG)
);

defparam rnode_390to391_bb4_and149_i_0_reg_391_fifo.DEPTH = 1;
defparam rnode_390to391_bb4_and149_i_0_reg_391_fifo.DATA_WIDTH = 32;
defparam rnode_390to391_bb4_and149_i_0_reg_391_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_390to391_bb4_and149_i_0_reg_391_fifo.IMPL = "shift_reg";

assign rnode_390to391_bb4_and149_i_0_reg_391_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and149_i_stall_in = 1'b0;
assign rnode_390to391_bb4_and149_i_0_stall_in_0_reg_391_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and149_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4_and149_i_0_NO_SHIFT_REG = rnode_390to391_bb4_and149_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_and149_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4_and149_i_1_NO_SHIFT_REG = rnode_390to391_bb4_and149_i_0_reg_391_NO_SHIFT_REG;
assign rnode_390to391_bb4_and149_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_390to391_bb4_and149_i_2_NO_SHIFT_REG = rnode_390to391_bb4_and149_i_0_reg_391_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__33_i211_stall_local;
wire [31:0] local_bb4__33_i211;

assign local_bb4__33_i211 = (local_bb4_tobool49_i ? (local_bb4__32_i210 & 32'hFFFFFF00) : (local_bb4_shl1_i18_i & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__35_i_stall_local;
wire [31:0] local_bb4__35_i;

assign local_bb4__35_i = (local_bb4_tobool49_i ? (local_bb4__34_i & 32'h1FFFFFF) : (local_bb4_or_i17_i & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__37_i_stall_local;
wire [31:0] local_bb4__37_i;

assign local_bb4__37_i = (local_bb4_tobool49_i ? (local_bb4__36_i & 32'h1FF) : (local_bb4_inc_i & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i_stall_local;
wire [31:0] local_bb4_and21_i;

assign local_bb4_and21_i = (rnode_390to391_bb4__22_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i_valid_out;
wire local_bb4_and20_i_stall_in;
wire local_bb4_and20_i_inputs_ready;
wire local_bb4_and20_i_stall_local;
wire [31:0] local_bb4_and20_i;

assign local_bb4_and20_i_inputs_ready = rnode_390to391_bb4__23_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i = (rnode_390to391_bb4__23_i_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i_valid_out = 1'b1;
assign rnode_390to391_bb4__23_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i_valid_out;
wire local_bb4_and35_i_stall_in;
wire local_bb4_and35_i_inputs_ready;
wire local_bb4_and35_i_stall_local;
wire [31:0] local_bb4_and35_i;

assign local_bb4_and35_i_inputs_ready = rnode_390to391_bb4__23_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i = (rnode_390to391_bb4__23_i_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i_valid_out = 1'b1;
assign rnode_390to391_bb4__23_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i_stall_local;
wire [31:0] local_bb4_xor_i;

assign local_bb4_xor_i = (rnode_390to391_bb4__23_i_2_NO_SHIFT_REG ^ rnode_390to391_bb4__22_i_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i_stall_local;
wire [31:0] local_bb4_and17_i;

assign local_bb4_and17_i = ((rnode_390to392_bb4_shr16_i_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_392to394_bb4_shr16_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to394_bb4_shr16_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to394_bb4_shr16_i_0_NO_SHIFT_REG;
 logic rnode_392to394_bb4_shr16_i_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to394_bb4_shr16_i_0_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_shr16_i_0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_shr16_i_0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_shr16_i_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_392to394_bb4_shr16_i_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to394_bb4_shr16_i_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to394_bb4_shr16_i_0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_392to394_bb4_shr16_i_0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_392to394_bb4_shr16_i_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in((rnode_390to392_bb4_shr16_i_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_392to394_bb4_shr16_i_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_392to394_bb4_shr16_i_0_reg_394_fifo.DEPTH = 2;
defparam rnode_392to394_bb4_shr16_i_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_392to394_bb4_shr16_i_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to394_bb4_shr16_i_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_392to394_bb4_shr16_i_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_390to392_bb4_shr16_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_shr16_i_0_NO_SHIFT_REG = rnode_392to394_bb4_shr16_i_0_reg_394_NO_SHIFT_REG;
assign rnode_392to394_bb4_shr16_i_0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_shr16_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp96_i_stall_local;
wire local_bb4_cmp96_i;

assign local_bb4_cmp96_i = ((rnode_390to391_bb4_and95_i_0_NO_SHIFT_REG & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp116_i_stall_local;
wire local_bb4_cmp116_i;

assign local_bb4_cmp116_i = ((rnode_390to391_bb4_and115_i_0_NO_SHIFT_REG & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp131_not_i_stall_local;
wire local_bb4_cmp131_not_i;

assign local_bb4_cmp131_not_i = ((rnode_390to391_bb4_and130_i_0_NO_SHIFT_REG & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i_stall_local;
wire local_bb4_Pivot20_i;

assign local_bb4_Pivot20_i = ((rnode_390to391_bb4_and149_i_1_NO_SHIFT_REG & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i_stall_local;
wire local_bb4_SwitchLeaf_i;

assign local_bb4_SwitchLeaf_i = ((rnode_390to391_bb4_and149_i_2_NO_SHIFT_REG & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i214_stall_local;
wire [31:0] local_bb4_and75_i214;

assign local_bb4_and75_i214 = ((local_bb4__35_i & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i211_valid_out;
wire local_bb4__33_i211_stall_in;
wire local_bb4__37_i_valid_out;
wire local_bb4__37_i_stall_in;
wire local_bb4_and75_i214_valid_out;
wire local_bb4_and75_i214_stall_in;
wire local_bb4_and83_i_valid_out;
wire local_bb4_and83_i_stall_in;
wire local_bb4_and83_i_inputs_ready;
wire local_bb4_and83_i_stall_local;
wire [31:0] local_bb4_and83_i;

assign local_bb4_and83_i_inputs_ready = (local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG & rnode_389to391_bb4_add_i206_0_valid_out_1_NO_SHIFT_REG & rnode_389to391_bb4_add_i206_0_valid_out_0_NO_SHIFT_REG & rnode_389to391_bb4_add_i206_0_valid_out_2_NO_SHIFT_REG & local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG);
assign local_bb4_and83_i = ((local_bb4__35_i & 32'h1FFFFFF) & 32'h1);
assign local_bb4__33_i211_valid_out = 1'b1;
assign local_bb4__37_i_valid_out = 1'b1;
assign local_bb4_and75_i214_valid_out = 1'b1;
assign local_bb4_and83_i_valid_out = 1'b1;
assign local_bb4_mul_i_i_stall_in_0 = 1'b0;
assign rnode_389to391_bb4_add_i206_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb4_add_i206_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_389to391_bb4_add_i206_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign local_bb4_mul_i_i_stall_in_1 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i_stall_local;
wire local_bb4_lnot33_not_i;

assign local_bb4_lnot33_not_i = ((local_bb4_and21_i & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or64_i_stall_local;
wire [31:0] local_bb4_or64_i;

assign local_bb4_or64_i = ((local_bb4_and21_i & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and20_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and20_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and20_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and20_i_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and20_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and20_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and20_i_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and20_i_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and20_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_and20_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_and20_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_and20_i_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_and20_i_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_and20_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i & 32'h7FFFFF)),
	.data_out(rnode_391to392_bb4_and20_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_and20_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_and20_i_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb4_and20_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_and20_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_and20_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i_stall_in = 1'b0;
assign rnode_391to392_bb4_and20_i_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4_and20_i_0_NO_SHIFT_REG = rnode_391to392_bb4_and20_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4_and20_i_1_NO_SHIFT_REG = rnode_391to392_bb4_and20_i_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and35_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and35_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and35_i_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and35_i_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and35_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_and35_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_and35_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_and35_i_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_and35_i_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_and35_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i & 32'h80000000)),
	.data_out(rnode_391to392_bb4_and35_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_and35_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_and35_i_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb4_and35_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_and35_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_and35_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i_stall_in = 1'b0;
assign rnode_391to392_bb4_and35_i_0_NO_SHIFT_REG = rnode_391to392_bb4_and35_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_and35_i_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp37_i_stall_local;
wire local_bb4_cmp37_i;

assign local_bb4_cmp37_i = ($signed(local_bb4_xor_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor_lobit_i_stall_local;
wire [31:0] local_bb4_xor_lobit_i;

assign local_bb4_xor_lobit_i = ($signed(local_bb4_xor_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and36_lobit_i_stall_local;
wire [31:0] local_bb4_and36_lobit_i;

assign local_bb4_and36_lobit_i = (local_bb4_xor_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i_stall_local;
wire local_bb4_lnot_i;

assign local_bb4_lnot_i = ((local_bb4_and17_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i5_stall_local;
wire local_bb4_cmp25_i5;

assign local_bb4_cmp25_i5 = ((local_bb4_and17_i & 32'hFF) == 32'hFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4__33_i211_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4__33_i211_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__33_i211_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4__33_i211_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4__33_i211_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__33_i211_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4__33_i211_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__33_i211_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4__33_i211_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4__33_i211_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4__33_i211_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4__33_i211_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4__33_i211_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4__33_i211_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4__33_i211_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4__33_i211_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb4__33_i211 & 32'hFFFFFF00)),
	.data_out(rnode_391to392_bb4__33_i211_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4__33_i211_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4__33_i211_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb4__33_i211_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4__33_i211_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4__33_i211_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__33_i211_stall_in = 1'b0;
assign rnode_391to392_bb4__33_i211_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4__33_i211_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4__33_i211_0_NO_SHIFT_REG = rnode_391to392_bb4__33_i211_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4__33_i211_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4__33_i211_1_NO_SHIFT_REG = rnode_391to392_bb4__33_i211_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4__37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__37_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__37_i_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__37_i_2_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__37_i_3_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4__37_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4__37_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4__37_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4__37_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4__37_i_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4__37_i_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4__37_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb4__37_i & 32'h3FF)),
	.data_out(rnode_391to392_bb4__37_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4__37_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4__37_i_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb4__37_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4__37_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4__37_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__37_i_stall_in = 1'b0;
assign rnode_391to392_bb4__37_i_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4__37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4__37_i_0_NO_SHIFT_REG = rnode_391to392_bb4__37_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4__37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4__37_i_1_NO_SHIFT_REG = rnode_391to392_bb4__37_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4__37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4__37_i_2_NO_SHIFT_REG = rnode_391to392_bb4__37_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4__37_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4__37_i_3_NO_SHIFT_REG = rnode_391to392_bb4__37_i_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_391to393_bb4_and75_i214_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to393_bb4_and75_i214_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to393_bb4_and75_i214_0_NO_SHIFT_REG;
 logic rnode_391to393_bb4_and75_i214_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to393_bb4_and75_i214_0_reg_393_NO_SHIFT_REG;
 logic rnode_391to393_bb4_and75_i214_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_391to393_bb4_and75_i214_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_391to393_bb4_and75_i214_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_391to393_bb4_and75_i214_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to393_bb4_and75_i214_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to393_bb4_and75_i214_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_391to393_bb4_and75_i214_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_391to393_bb4_and75_i214_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in((local_bb4_and75_i214 & 32'h7FFFFF)),
	.data_out(rnode_391to393_bb4_and75_i214_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_391to393_bb4_and75_i214_0_reg_393_fifo.DEPTH = 2;
defparam rnode_391to393_bb4_and75_i214_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_391to393_bb4_and75_i214_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to393_bb4_and75_i214_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_391to393_bb4_and75_i214_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and75_i214_stall_in = 1'b0;
assign rnode_391to393_bb4_and75_i214_0_NO_SHIFT_REG = rnode_391to393_bb4_and75_i214_0_reg_393_NO_SHIFT_REG;
assign rnode_391to393_bb4_and75_i214_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_391to393_bb4_and75_i214_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_and83_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and83_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and83_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and83_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and83_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and83_i_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and83_i_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and83_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_and83_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_and83_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_and83_i_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_and83_i_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_and83_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb4_and83_i & 32'h1)),
	.data_out(rnode_391to392_bb4_and83_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_and83_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_and83_i_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb4_and83_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_and83_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_and83_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and83_i_stall_in = 1'b0;
assign rnode_391to392_bb4_and83_i_0_NO_SHIFT_REG = rnode_391to392_bb4_and83_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_and83_i_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and83_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shl65_i_stall_local;
wire [31:0] local_bb4_shl65_i;

assign local_bb4_shl65_i = ((local_bb4_or64_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i_stall_local;
wire local_bb4_lnot30_i;

assign local_bb4_lnot30_i = ((rnode_391to392_bb4_and20_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i6_stall_local;
wire [31:0] local_bb4_or_i6;

assign local_bb4_or_i6 = ((rnode_391to392_bb4_and20_i_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_392to394_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to394_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and35_i_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to394_bb4_and35_i_0_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and35_i_0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and35_i_0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and35_i_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_392to394_bb4_and35_i_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to394_bb4_and35_i_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to394_bb4_and35_i_0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_392to394_bb4_and35_i_0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_392to394_bb4_and35_i_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in((rnode_391to392_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_392to394_bb4_and35_i_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_392to394_bb4_and35_i_0_reg_394_fifo.DEPTH = 2;
defparam rnode_392to394_bb4_and35_i_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_392to394_bb4_and35_i_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to394_bb4_and35_i_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_392to394_bb4_and35_i_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_and35_i_0_NO_SHIFT_REG = rnode_392to394_bb4_and35_i_0_reg_394_NO_SHIFT_REG;
assign rnode_392to394_bb4_and35_i_0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i_stall_local;
wire local_bb4_cmp25_not_i;

assign local_bb4_cmp25_not_i = (local_bb4_cmp25_i5 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u88_stall_local;
wire local_bb4_var__u88;

assign local_bb4_var__u88 = (local_bb4_cmp25_i5 | rnode_390to392_bb4_cmp27_i_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i_stall_local;
wire local_bb4_cmp77_i;

assign local_bb4_cmp77_i = ((rnode_391to392_bb4__33_i211_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u89_stall_local;
wire local_bb4_var__u89;

assign local_bb4_var__u89 = ($signed((rnode_391to392_bb4__33_i211_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp53_i_stall_local;
wire local_bb4_cmp53_i;

assign local_bb4_cmp53_i = ((rnode_391to392_bb4__37_i_0_NO_SHIFT_REG & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp68_i_valid_out;
wire local_bb4_cmp68_i_stall_in;
wire local_bb4_cmp68_i_inputs_ready;
wire local_bb4_cmp68_i_stall_local;
wire local_bb4_cmp68_i;

assign local_bb4_cmp68_i_inputs_ready = rnode_391to392_bb4__37_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp68_i = ((rnode_391to392_bb4__37_i_1_NO_SHIFT_REG & 32'h3FF) < 32'h80);
assign local_bb4_cmp68_i_valid_out = 1'b1;
assign rnode_391to392_bb4__37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i215_stall_local;
wire [31:0] local_bb4_sub_i215;

assign local_bb4_sub_i215 = ((rnode_391to392_bb4__37_i_2_NO_SHIFT_REG & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp71_not_i_valid_out;
wire local_bb4_cmp71_not_i_stall_in;
wire local_bb4_cmp71_not_i_inputs_ready;
wire local_bb4_cmp71_not_i_stall_local;
wire local_bb4_cmp71_not_i;

assign local_bb4_cmp71_not_i_inputs_ready = rnode_391to392_bb4__37_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4_cmp71_not_i = ((rnode_391to392_bb4__37_i_3_NO_SHIFT_REG & 32'h3FF) != 32'h7F);
assign local_bb4_cmp71_not_i_valid_out = 1'b1;
assign rnode_391to392_bb4__37_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool84_i_stall_local;
wire local_bb4_tobool84_i;

assign local_bb4_tobool84_i = ((rnode_391to392_bb4_and83_i_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i_stall_local;
wire [31:0] local_bb4__28_i;

assign local_bb4__28_i = (rnode_390to391_bb4_lnot23_i_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl65_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i_stall_local;
wire local_bb4_lnot30_not_i;

assign local_bb4_lnot30_not_i = (local_bb4_lnot30_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i7_stall_local;
wire [31:0] local_bb4_shl_i7;

assign local_bb4_shl_i7 = ((local_bb4_or_i6 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and35_i_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_and35_i_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and35_i_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and35_i_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and35_i_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_and35_i_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_and35_i_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_and35_i_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_and35_i_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_and35_i_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in((rnode_392to394_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_394to395_bb4_and35_i_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_and35_i_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_and35_i_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_394to395_bb4_and35_i_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_and35_i_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_and35_i_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_392to394_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_and35_i_0_NO_SHIFT_REG = rnode_394to395_bb4_and35_i_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_and35_i_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i_stall_local;
wire local_bb4_or_cond_i;

assign local_bb4_or_cond_i = (local_bb4_lnot30_i | local_bb4_cmp25_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or581_i_valid_out;
wire local_bb4_or581_i_stall_in;
wire local_bb4_or581_i_inputs_ready;
wire local_bb4_or581_i_stall_local;
wire local_bb4_or581_i;

assign local_bb4_or581_i_inputs_ready = (rnode_391to392_bb4_var__u86_0_valid_out_NO_SHIFT_REG & rnode_391to392_bb4__37_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_or581_i = (rnode_391to392_bb4_var__u86_0_NO_SHIFT_REG | local_bb4_cmp53_i);
assign local_bb4_or581_i_valid_out = 1'b1;
assign rnode_391to392_bb4_var__u86_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4__37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_cmp68_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp68_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp68_i_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp68_i_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp68_i_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp68_i_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp68_i_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp68_i_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_cmp68_i_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_cmp68_i_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_cmp68_i_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_cmp68_i_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_cmp68_i_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb4_cmp68_i),
	.data_out(rnode_392to393_bb4_cmp68_i_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_cmp68_i_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_cmp68_i_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4_cmp68_i_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_cmp68_i_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_cmp68_i_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp68_i_stall_in = 1'b0;
assign rnode_392to393_bb4_cmp68_i_0_NO_SHIFT_REG = rnode_392to393_bb4_cmp68_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_cmp68_i_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_cmp68_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and74_i_stall_local;
wire [31:0] local_bb4_and74_i;

assign local_bb4_and74_i = ((local_bb4_sub_i215 & 32'hFF800000) + 32'h40800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_cmp71_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp71_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp71_not_i_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp71_not_i_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp71_not_i_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp71_not_i_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp71_not_i_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_cmp71_not_i_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_cmp71_not_i_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_cmp71_not_i_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_cmp71_not_i_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_cmp71_not_i_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_cmp71_not_i_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb4_cmp71_not_i),
	.data_out(rnode_392to393_bb4_cmp71_not_i_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_cmp71_not_i_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_cmp71_not_i_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4_cmp71_not_i_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_cmp71_not_i_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_cmp71_not_i_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp71_not_i_stall_in = 1'b0;
assign rnode_392to393_bb4_cmp71_not_i_0_NO_SHIFT_REG = rnode_392to393_bb4_cmp71_not_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_cmp71_not_i_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_cmp71_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__39_i_stall_local;
wire local_bb4__39_i;

assign local_bb4__39_i = (local_bb4_tobool84_i & local_bb4_var__u89);

// This section implements an unregistered operation.
// 
wire local_bb4_and72_i_stall_local;
wire [31:0] local_bb4_and72_i;

assign local_bb4_and72_i = ((local_bb4__28_i & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i_stall_local;
wire [31:0] local_bb4_and75_i;

assign local_bb4_and75_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and78_i_stall_local;
wire [31:0] local_bb4_and78_i;

assign local_bb4_and78_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr94_i_stall_local;
wire [31:0] local_bb4_shr94_i;

assign local_bb4_shr94_i = ((local_bb4__28_i & 32'h7FFFFF8) >> (rnode_390to391_bb4_and93_i_0_NO_SHIFT_REG & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i_stall_local;
wire [31:0] local_bb4_and90_i;

assign local_bb4_and90_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and87_i_stall_local;
wire [31:0] local_bb4_and87_i;

assign local_bb4_and87_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and84_i_stall_local;
wire [31:0] local_bb4_and84_i;

assign local_bb4_and84_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u90_stall_local;
wire [31:0] local_bb4_var__u90;

assign local_bb4_var__u90 = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i_stall_local;
wire local_bb4_or_cond_not_i;

assign local_bb4_or_cond_not_i = (local_bb4_cmp25_i5 & local_bb4_lnot30_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i_stall_local;
wire [31:0] local_bb4__27_i;

assign local_bb4__27_i = (local_bb4_lnot_i ? 32'h0 : ((local_bb4_shl_i7 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i_stall_local;
wire local_bb4_reduction_8_i;

assign local_bb4_reduction_8_i = (rnode_390to392_bb4_cmp27_i_1_NO_SHIFT_REG & local_bb4_or_cond_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_or581_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_1_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_valid_out_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_stall_in_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_or581_i_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_or581_i_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_or581_i_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_or581_i_0_stall_in_0_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_or581_i_0_valid_out_0_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_or581_i_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb4_or581_i),
	.data_out(rnode_392to393_bb4_or581_i_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_or581_i_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_or581_i_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4_or581_i_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_or581_i_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_or581_i_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or581_i_stall_in = 1'b0;
assign rnode_392to393_bb4_or581_i_0_stall_in_0_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_or581_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4_or581_i_0_NO_SHIFT_REG = rnode_392to393_bb4_or581_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_or581_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4_or581_i_1_NO_SHIFT_REG = rnode_392to393_bb4_or581_i_0_reg_393_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u91_stall_local;
wire [31:0] local_bb4_var__u91;

assign local_bb4_var__u91[31:1] = 31'h0;
assign local_bb4_var__u91[0] = rnode_392to393_bb4_cmp68_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i216_valid_out;
wire local_bb4_shl_i216_stall_in;
wire local_bb4_shl_i216_inputs_ready;
wire local_bb4_shl_i216_stall_local;
wire [31:0] local_bb4_shl_i216;

assign local_bb4_shl_i216_inputs_ready = rnode_391to392_bb4__37_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shl_i216 = ((local_bb4_and74_i & 32'hFF800000) & 32'h7F800000);
assign local_bb4_shl_i216_valid_out = 1'b1;
assign rnode_391to392_bb4__37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__40_i_valid_out;
wire local_bb4__40_i_stall_in;
wire local_bb4__40_i_inputs_ready;
wire local_bb4__40_i_stall_local;
wire local_bb4__40_i;

assign local_bb4__40_i_inputs_ready = (rnode_391to392_bb4__33_i211_0_valid_out_0_NO_SHIFT_REG & rnode_391to392_bb4__33_i211_0_valid_out_1_NO_SHIFT_REG & rnode_391to392_bb4_and83_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40_i = (local_bb4_cmp77_i | local_bb4__39_i);
assign local_bb4__40_i_valid_out = 1'b1;
assign rnode_391to392_bb4__33_i211_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4__33_i211_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and83_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and72_tr_i_stall_local;
wire [7:0] local_bb4_and72_tr_i;
wire [31:0] local_bb4_and72_tr_i$ps;

assign local_bb4_and72_tr_i$ps = (local_bb4_and72_i & 32'hFFFFFF);
assign local_bb4_and72_tr_i = local_bb4_and72_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp76_i_stall_local;
wire local_bb4_cmp76_i;

assign local_bb4_cmp76_i = ((local_bb4_and75_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp79_i_stall_local;
wire local_bb4_cmp79_i;

assign local_bb4_cmp79_i = ((local_bb4_and78_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and142_i_stall_local;
wire [31:0] local_bb4_and142_i;

assign local_bb4_and142_i = (local_bb4_shr94_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr150_i_stall_local;
wire [31:0] local_bb4_shr150_i;

assign local_bb4_shr150_i = (local_bb4_shr94_i >> (rnode_390to391_bb4_and149_i_0_NO_SHIFT_REG & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u92_stall_local;
wire [31:0] local_bb4_var__u92;

assign local_bb4_var__u92 = (local_bb4_shr94_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and146_i_stall_local;
wire [31:0] local_bb4_and146_i;

assign local_bb4_and146_i = (local_bb4_shr94_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i_stall_local;
wire local_bb4_cmp91_i;

assign local_bb4_cmp91_i = ((local_bb4_and90_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp88_i_stall_local;
wire local_bb4_cmp88_i;

assign local_bb4_cmp88_i = ((local_bb4_and87_i & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp85_i_stall_local;
wire local_bb4_cmp85_i;

assign local_bb4_cmp85_i = ((local_bb4_and84_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u93_stall_local;
wire local_bb4_var__u93;

assign local_bb4_var__u93 = ((local_bb4_var__u90 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i213_stall_local;
wire local_bb4_reduction_2_i213;

assign local_bb4_reduction_2_i213 = (rnode_392to393_bb4_reduction_0_i212_0_NO_SHIFT_REG | rnode_392to393_bb4_or581_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cond111_i_stall_local;
wire [31:0] local_bb4_cond111_i;

assign local_bb4_cond111_i = (rnode_392to393_bb4_or581_i_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_shl_i216_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_shl_i216_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_shl_i216_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_shl_i216_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_shl_i216_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_shl_i216_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_shl_i216_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_shl_i216_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_shl_i216_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_shl_i216_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_shl_i216_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_shl_i216_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_shl_i216_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in((local_bb4_shl_i216 & 32'h7F800000)),
	.data_out(rnode_392to393_bb4_shl_i216_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_shl_i216_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_shl_i216_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_392to393_bb4_shl_i216_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_shl_i216_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_shl_i216_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shl_i216_stall_in = 1'b0;
assign rnode_392to393_bb4_shl_i216_0_NO_SHIFT_REG = rnode_392to393_bb4_shl_i216_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_shl_i216_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_shl_i216_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4__40_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4__40_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4__40_i_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4__40_i_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4__40_i_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__40_i_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__40_i_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__40_i_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4__40_i_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4__40_i_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4__40_i_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4__40_i_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4__40_i_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb4__40_i),
	.data_out(rnode_392to393_bb4__40_i_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4__40_i_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4__40_i_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4__40_i_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4__40_i_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4__40_i_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_i_stall_in = 1'b0;
assign rnode_392to393_bb4__40_i_0_NO_SHIFT_REG = rnode_392to393_bb4__40_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4__40_i_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4__40_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_frombool74_i_stall_local;
wire [7:0] local_bb4_frombool74_i;

assign local_bb4_frombool74_i = (local_bb4_and72_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u94_stall_local;
wire [31:0] local_bb4_var__u94;

assign local_bb4_var__u94 = ((local_bb4_and146_i & 32'h3FFFFFFF) | local_bb4_shr94_i);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i_stall_local;
wire local_bb4__31_v_i;

assign local_bb4__31_v_i = (local_bb4_cmp96_i ? local_bb4_cmp79_i : local_bb4_cmp91_i);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i_stall_local;
wire local_bb4__30_v_i;

assign local_bb4__30_v_i = (local_bb4_cmp96_i ? local_bb4_cmp76_i : local_bb4_cmp88_i);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool109_i_stall_local;
wire [7:0] local_bb4_frombool109_i;

assign local_bb4_frombool109_i[7:1] = 7'h0;
assign local_bb4_frombool109_i[0] = local_bb4_cmp85_i;

// This section implements an unregistered operation.
// 
wire local_bb4_or107_i_stall_local;
wire [31:0] local_bb4_or107_i;

assign local_bb4_or107_i[31:1] = 31'h0;
assign local_bb4_or107_i[0] = local_bb4_var__u93;

// This section implements an unregistered operation.
// 
wire local_bb4_conv101_i_stall_local;
wire [31:0] local_bb4_conv101_i;

assign local_bb4_conv101_i[31:1] = 31'h0;
assign local_bb4_conv101_i[0] = local_bb4_reduction_2_i213;

// This section implements an unregistered operation.
// 
wire local_bb4_or76_i_stall_local;
wire [31:0] local_bb4_or76_i;

assign local_bb4_or76_i = ((rnode_392to393_bb4_shl_i216_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_391to393_bb4_and75_i214_0_NO_SHIFT_REG & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond_i217_stall_local;
wire [31:0] local_bb4_cond_i217;

assign local_bb4_cond_i217[31:1] = 31'h0;
assign local_bb4_cond_i217[0] = rnode_392to393_bb4__40_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or1596_i_stall_local;
wire [31:0] local_bb4_or1596_i;

assign local_bb4_or1596_i = (local_bb4_var__u94 | (local_bb4_and142_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i_stall_local;
wire [7:0] local_bb4__31_i;

assign local_bb4__31_i[7:1] = 7'h0;
assign local_bb4__31_i[0] = local_bb4__31_v_i;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i_stall_local;
wire [7:0] local_bb4__30_i;

assign local_bb4__30_i[7:1] = 7'h0;
assign local_bb4__30_i[0] = local_bb4__30_v_i;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i_stall_local;
wire [7:0] local_bb4__29_i;

assign local_bb4__29_i = (local_bb4_cmp96_i ? (local_bb4_frombool74_i & 8'h1) : (local_bb4_frombool109_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i_stall_local;
wire [31:0] local_bb4__32_i;

assign local_bb4__32_i = (local_bb4_cmp96_i ? 32'h0 : (local_bb4_or107_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_add87_i_stall_local;
wire [31:0] local_bb4_add87_i;

assign local_bb4_add87_i = ((local_bb4_cond_i217 & 32'h1) + (local_bb4_or76_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_or162_i_stall_local;
wire [31:0] local_bb4_or162_i;

assign local_bb4_or162_i = (local_bb4_or1596_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1237_i_stall_local;
wire [7:0] local_bb4_or1237_i;

assign local_bb4_or1237_i = ((local_bb4__30_i & 8'h1) | (local_bb4__29_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i_stall_local;
wire [7:0] local_bb4__33_i;

assign local_bb4__33_i = (local_bb4_cmp116_i ? (local_bb4__29_i & 8'h1) : (local_bb4__31_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i_stall_local;
wire [31:0] local_bb4_and88_i;

assign local_bb4_and88_i = (local_bb4_add87_i & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i218_stall_local;
wire [31:0] local_bb4_and90_i218;

assign local_bb4_and90_i218 = (local_bb4_add87_i & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i_stall_local;
wire [31:0] local_bb4__37_v_i;

assign local_bb4__37_v_i = (local_bb4_Pivot20_i ? 32'h0 : (local_bb4_or162_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or123_i_stall_local;
wire [31:0] local_bb4_or123_i;

assign local_bb4_or123_i[31:8] = 24'h0;
assign local_bb4_or123_i[7:0] = (local_bb4_or1237_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u95_stall_local;
wire [7:0] local_bb4_var__u95;

assign local_bb4_var__u95 = ((local_bb4__33_i & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or89_i_stall_local;
wire [31:0] local_bb4_or89_i;

assign local_bb4_or89_i = ((local_bb4_and88_i & 32'h7FFFFFFF) | (local_bb4_and4_i & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i219_stall_local;
wire local_bb4_cmp91_i219;

assign local_bb4_cmp91_i219 = ((local_bb4_and90_i218 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i_stall_local;
wire [31:0] local_bb4__39_v_i;

assign local_bb4__39_v_i = (local_bb4_SwitchLeaf_i ? (local_bb4_var__u92 & 32'h1) : (local_bb4__37_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i_stall_local;
wire [31:0] local_bb4_or124_i;

assign local_bb4_or124_i = (local_bb4_cmp116_i ? 32'h0 : (local_bb4_or123_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv135_i_stall_local;
wire [31:0] local_bb4_conv135_i;

assign local_bb4_conv135_i[31:8] = 24'h0;
assign local_bb4_conv135_i[7:0] = (local_bb4_var__u95 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge14_i_stall_local;
wire local_bb4_brmerge14_i;

assign local_bb4_brmerge14_i = (local_bb4_cmp91_i219 | rnode_392to393_bb4_cmp71_not_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i_stall_local;
wire [31:0] local_bb4_reduction_3_i;

assign local_bb4_reduction_3_i = ((local_bb4__32_i & 32'h1) | (local_bb4_or124_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or136_i_stall_local;
wire [31:0] local_bb4_or136_i;

assign local_bb4_or136_i = (local_bb4_cmp131_not_i ? (local_bb4_conv135_i & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_conv99_i_stall_local;
wire [31:0] local_bb4_conv99_i;

assign local_bb4_conv99_i = (local_bb4_brmerge14_i ? (local_bb4_var__u91 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i_stall_local;
wire [31:0] local_bb4_reduction_5_i;

assign local_bb4_reduction_5_i = (local_bb4_shr150_i | (local_bb4_reduction_3_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i_stall_local;
wire [31:0] local_bb4_reduction_4_i;

assign local_bb4_reduction_4_i = ((local_bb4_or136_i & 32'h1) | (local_bb4__39_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or102_i_stall_local;
wire [31:0] local_bb4_or102_i;

assign local_bb4_or102_i = ((local_bb4_conv99_i & 32'h1) | (local_bb4_conv101_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i_stall_local;
wire [31:0] local_bb4_reduction_6_i;

assign local_bb4_reduction_6_i = ((local_bb4_reduction_4_i & 32'h1) | local_bb4_reduction_5_i);

// This section implements an unregistered operation.
// 
wire local_bb4_tobool103_i_stall_local;
wire local_bb4_tobool103_i;

assign local_bb4_tobool103_i = ((local_bb4_or102_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i_valid_out;
wire local_bb4_lnot33_not_i_stall_in;
wire local_bb4_cmp37_i_valid_out;
wire local_bb4_cmp37_i_stall_in;
wire local_bb4_and36_lobit_i_valid_out;
wire local_bb4_and36_lobit_i_stall_in;
wire local_bb4_xor188_i_valid_out;
wire local_bb4_xor188_i_stall_in;
wire local_bb4_xor188_i_inputs_ready;
wire local_bb4_xor188_i_stall_local;
wire [31:0] local_bb4_xor188_i;

assign local_bb4_xor188_i_inputs_ready = (rnode_390to391_bb4__22_i_0_valid_out_0_NO_SHIFT_REG & rnode_390to391_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG & rnode_390to391_bb4_and93_i_0_valid_out_NO_SHIFT_REG & rnode_390to391_bb4_and149_i_0_valid_out_0_NO_SHIFT_REG & rnode_390to391_bb4_and95_i_0_valid_out_NO_SHIFT_REG & rnode_390to391_bb4_and149_i_0_valid_out_2_NO_SHIFT_REG & rnode_390to391_bb4_and115_i_0_valid_out_NO_SHIFT_REG & rnode_390to391_bb4_and130_i_0_valid_out_NO_SHIFT_REG & rnode_390to391_bb4_and149_i_0_valid_out_1_NO_SHIFT_REG & rnode_390to391_bb4__23_i_0_valid_out_2_NO_SHIFT_REG & rnode_390to391_bb4__22_i_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor188_i = (local_bb4_reduction_6_i ^ local_bb4_xor_lobit_i);
assign local_bb4_lnot33_not_i_valid_out = 1'b1;
assign local_bb4_cmp37_i_valid_out = 1'b1;
assign local_bb4_and36_lobit_i_valid_out = 1'b1;
assign local_bb4_xor188_i_valid_out = 1'b1;
assign rnode_390to391_bb4__22_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_lnot23_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and93_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and149_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and95_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and149_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and115_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and130_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4_and149_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4__23_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_390to391_bb4__22_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cond107_i_stall_local;
wire [31:0] local_bb4_cond107_i;

assign local_bb4_cond107_i = (local_bb4_tobool103_i ? (local_bb4_and4_i & 32'h80000000) : 32'hFFFFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb4_lnot33_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_391to392_bb4_lnot33_not_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_lnot33_not_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_391to392_bb4_lnot33_not_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_lnot33_not_i_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_lnot33_not_i_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_lnot33_not_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_lnot33_not_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_lnot33_not_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_lnot33_not_i_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_lnot33_not_i_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_lnot33_not_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i),
	.data_out(rnode_391to392_bb4_lnot33_not_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_lnot33_not_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_lnot33_not_i_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_391to392_bb4_lnot33_not_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_lnot33_not_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_lnot33_not_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i_stall_in = 1'b0;
assign rnode_391to392_bb4_lnot33_not_i_0_NO_SHIFT_REG = rnode_391to392_bb4_lnot33_not_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_lnot33_not_i_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_valid_out_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_stall_in_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_cmp37_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_cmp37_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_cmp37_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_cmp37_i_0_stall_in_0_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_cmp37_i_0_valid_out_0_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_cmp37_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(local_bb4_cmp37_i),
	.data_out(rnode_391to392_bb4_cmp37_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_cmp37_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_cmp37_i_0_reg_392_fifo.DATA_WIDTH = 1;
defparam rnode_391to392_bb4_cmp37_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_cmp37_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_cmp37_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp37_i_stall_in = 1'b0;
assign rnode_391to392_bb4_cmp37_i_0_stall_in_0_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4_cmp37_i_0_NO_SHIFT_REG = rnode_391to392_bb4_cmp37_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4_cmp37_i_1_NO_SHIFT_REG = rnode_391to392_bb4_cmp37_i_0_reg_392_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and36_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and36_lobit_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and36_lobit_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_and36_lobit_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and36_lobit_i_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and36_lobit_i_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_and36_lobit_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_and36_lobit_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_and36_lobit_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_and36_lobit_i_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_and36_lobit_i_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_and36_lobit_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in((local_bb4_and36_lobit_i & 32'h1)),
	.data_out(rnode_391to392_bb4_and36_lobit_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_and36_lobit_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_and36_lobit_i_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb4_and36_lobit_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_and36_lobit_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_and36_lobit_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and36_lobit_i_stall_in = 1'b0;
assign rnode_391to392_bb4_and36_lobit_i_0_NO_SHIFT_REG = rnode_391to392_bb4_and36_lobit_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_and36_lobit_i_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_391to392_bb4_xor188_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_391to392_bb4_xor188_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_xor188_i_0_NO_SHIFT_REG;
 logic rnode_391to392_bb4_xor188_i_0_reg_392_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_391to392_bb4_xor188_i_0_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_xor188_i_0_valid_out_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_xor188_i_0_stall_in_reg_392_NO_SHIFT_REG;
 logic rnode_391to392_bb4_xor188_i_0_stall_out_reg_392_NO_SHIFT_REG;

acl_data_fifo rnode_391to392_bb4_xor188_i_0_reg_392_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_391to392_bb4_xor188_i_0_reg_392_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_391to392_bb4_xor188_i_0_stall_in_reg_392_NO_SHIFT_REG),
	.valid_out(rnode_391to392_bb4_xor188_i_0_valid_out_reg_392_NO_SHIFT_REG),
	.stall_out(rnode_391to392_bb4_xor188_i_0_stall_out_reg_392_NO_SHIFT_REG),
	.data_in(local_bb4_xor188_i),
	.data_out(rnode_391to392_bb4_xor188_i_0_reg_392_NO_SHIFT_REG)
);

defparam rnode_391to392_bb4_xor188_i_0_reg_392_fifo.DEPTH = 1;
defparam rnode_391to392_bb4_xor188_i_0_reg_392_fifo.DATA_WIDTH = 32;
defparam rnode_391to392_bb4_xor188_i_0_reg_392_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_391to392_bb4_xor188_i_0_reg_392_fifo.IMPL = "shift_reg";

assign rnode_391to392_bb4_xor188_i_0_reg_392_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor188_i_stall_in = 1'b0;
assign rnode_391to392_bb4_xor188_i_0_NO_SHIFT_REG = rnode_391to392_bb4_xor188_i_0_reg_392_NO_SHIFT_REG;
assign rnode_391to392_bb4_xor188_i_0_stall_in_reg_392_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_xor188_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and108_i_stall_local;
wire [31:0] local_bb4_and108_i;

assign local_bb4_and108_i = (local_bb4_cond107_i & local_bb4_or89_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i_stall_local;
wire local_bb4_brmerge_not_i;

assign local_bb4_brmerge_not_i = (rnode_390to392_bb4_cmp27_i_0_NO_SHIFT_REG & rnode_391to392_bb4_lnot33_not_i_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_392to394_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_2_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_valid_out_0_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_stall_in_0_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_cmp37_i_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_392to394_bb4_cmp37_i_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to394_bb4_cmp37_i_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to394_bb4_cmp37_i_0_stall_in_0_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_392to394_bb4_cmp37_i_0_valid_out_0_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_392to394_bb4_cmp37_i_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in(rnode_391to392_bb4_cmp37_i_1_NO_SHIFT_REG),
	.data_out(rnode_392to394_bb4_cmp37_i_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_392to394_bb4_cmp37_i_0_reg_394_fifo.DEPTH = 2;
defparam rnode_392to394_bb4_cmp37_i_0_reg_394_fifo.DATA_WIDTH = 1;
defparam rnode_392to394_bb4_cmp37_i_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to394_bb4_cmp37_i_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_392to394_bb4_cmp37_i_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_391to392_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_cmp37_i_0_stall_in_0_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_392to394_bb4_cmp37_i_0_NO_SHIFT_REG = rnode_392to394_bb4_cmp37_i_0_reg_394_NO_SHIFT_REG;
assign rnode_392to394_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_392to394_bb4_cmp37_i_1_NO_SHIFT_REG = rnode_392to394_bb4_cmp37_i_0_reg_394_NO_SHIFT_REG;
assign rnode_392to394_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_392to394_bb4_cmp37_i_2_NO_SHIFT_REG = rnode_392to394_bb4_cmp37_i_0_reg_394_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i8_stall_local;
wire [31:0] local_bb4_add_i8;

assign local_bb4_add_i8 = ((local_bb4__27_i & 32'h7FFFFF8) | (rnode_391to392_bb4_and36_lobit_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or112_i_stall_local;
wire [31:0] local_bb4_or112_i;

assign local_bb4_or112_i = (local_bb4_and108_i | (local_bb4_cond111_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4__24_i_stall_local;
wire local_bb4__24_i;

assign local_bb4__24_i = (local_bb4_or_cond_not_i | local_bb4_brmerge_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i_stall_local;
wire local_bb4_brmerge_not_not_i;

assign local_bb4_brmerge_not_not_i = (local_bb4_brmerge_not_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp37_i_stall_local;
wire local_bb4_not_cmp37_i;

assign local_bb4_not_cmp37_i = (rnode_392to394_bb4_cmp37_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add192_i_stall_local;
wire [31:0] local_bb4_add192_i;

assign local_bb4_add192_i = ((local_bb4_add_i8 & 32'h7FFFFF9) + rnode_391to392_bb4_xor188_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u96_valid_out;
wire local_bb4_var__u96_stall_in;
wire local_bb4_var__u96_inputs_ready;
wire local_bb4_var__u96_stall_local;
wire [31:0] local_bb4_var__u96;

assign local_bb4_var__u96_inputs_ready = (rnode_392to393_bb4_xor_i195_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb4__29_i204_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb4_or581_i_0_valid_out_1_NO_SHIFT_REG & rnode_392to393_bb4_or581_i_0_valid_out_0_NO_SHIFT_REG & rnode_392to393_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb4_cmp68_i_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb4_cmp71_not_i_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb4_shl_i216_0_valid_out_NO_SHIFT_REG & rnode_391to393_bb4_and75_i214_0_valid_out_NO_SHIFT_REG & rnode_392to393_bb4__40_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_var__u96 = (rnode_392to393_bb4__29_i204_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb4_or112_i);
assign local_bb4_var__u96_valid_out = 1'b1;
assign rnode_392to393_bb4_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_or581_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_or581_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_cmp68_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_cmp71_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_shl_i216_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to393_bb4_and75_i214_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4__40_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i_stall_local;
wire local_bb4_reduction_7_i;

assign local_bb4_reduction_7_i = (local_bb4_cmp25_i5 & local_bb4_brmerge_not_not_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb4_var__u96_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_var__u96_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_var__u96_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_var__u96_2_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_var__u96_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_valid_out_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_stall_in_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u96_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb4_var__u96_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb4_var__u96_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb4_var__u96_0_stall_in_0_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb4_var__u96_0_valid_out_0_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb4_var__u96_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in(local_bb4_var__u96),
	.data_out(rnode_393to394_bb4_var__u96_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb4_var__u96_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb4_var__u96_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb4_var__u96_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb4_var__u96_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb4_var__u96_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u96_stall_in = 1'b0;
assign rnode_393to394_bb4_var__u96_0_stall_in_0_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_var__u96_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_var__u96_0_NO_SHIFT_REG = rnode_393to394_bb4_var__u96_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_var__u96_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_var__u96_1_NO_SHIFT_REG = rnode_393to394_bb4_var__u96_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_var__u96_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_var__u96_2_NO_SHIFT_REG = rnode_393to394_bb4_var__u96_0_reg_394_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i_stall_local;
wire local_bb4_reduction_9_i;

assign local_bb4_reduction_9_i = (local_bb4_reduction_7_i & local_bb4_reduction_8_i);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i11_stall_local;
wire [31:0] local_bb4_and_i11;

assign local_bb4_and_i11 = (rnode_393to394_bb4_var__u96_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i17_stall_local;
wire [31:0] local_bb4_and10_i17;

assign local_bb4_and10_i17 = (rnode_393to394_bb4_var__u96_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_var__u96_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u96_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_var__u96_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u96_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u96_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_var__u96_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u96_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_var__u96_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u96_0_valid_out_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u96_0_stall_in_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u96_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_var__u96_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_var__u96_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_var__u96_0_stall_in_0_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_var__u96_0_valid_out_0_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_var__u96_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(rnode_393to394_bb4_var__u96_2_NO_SHIFT_REG),
	.data_out(rnode_394to395_bb4_var__u96_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_var__u96_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_var__u96_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_394to395_bb4_var__u96_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_var__u96_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_var__u96_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_var__u96_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u96_0_stall_in_0_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u96_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4_var__u96_0_NO_SHIFT_REG = rnode_394to395_bb4_var__u96_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_var__u96_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4_var__u96_1_NO_SHIFT_REG = rnode_394to395_bb4_var__u96_0_reg_395_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i_valid_out_2;
wire local_bb4_and17_i_stall_in_2;
wire local_bb4_var__u88_valid_out;
wire local_bb4_var__u88_stall_in;
wire local_bb4_add192_i_valid_out;
wire local_bb4_add192_i_stall_in;
wire local_bb4__26_i_valid_out;
wire local_bb4__26_i_stall_in;
wire local_bb4__26_i_inputs_ready;
wire local_bb4__26_i_stall_local;
wire local_bb4__26_i;

assign local_bb4__26_i_inputs_ready = (rnode_390to392_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG & rnode_390to392_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG & rnode_391to392_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_391to392_bb4_xor188_i_0_valid_out_NO_SHIFT_REG & rnode_391to392_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG & rnode_390to392_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG & rnode_391to392_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG & rnode_390to392_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG & rnode_391to392_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG & rnode_391to392_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i = (local_bb4_reduction_9_i ? rnode_391to392_bb4_cmp37_i_0_NO_SHIFT_REG : local_bb4__24_i);
assign local_bb4_and17_i_valid_out_2 = 1'b1;
assign local_bb4_var__u88_valid_out = 1'b1;
assign local_bb4_add192_i_valid_out = 1'b1;
assign local_bb4__26_i_valid_out = 1'b1;
assign rnode_390to392_bb4_shr16_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4_cmp27_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and36_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_xor188_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and20_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4_cmp27_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_lnot33_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_390to392_bb4_cmp27_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_and20_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_391to392_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i12_stall_local;
wire [31:0] local_bb4_shr_i12;

assign local_bb4_shr_i12 = ((local_bb4_and_i11 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i19_stall_local;
wire local_bb4_cmp13_i19;

assign local_bb4_cmp13_i19 = ((local_bb4_and10_i17 & 32'hFFFF) > (local_bb4_and12_i18 & 32'hFFFF));

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_392to394_bb4_and17_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and17_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_392to394_bb4_and17_i_0_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and17_i_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to394_bb4_and17_i_0_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and17_i_0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and17_i_0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_392to394_bb4_and17_i_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_392to394_bb4_and17_i_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to394_bb4_and17_i_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to394_bb4_and17_i_0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_392to394_bb4_and17_i_0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_392to394_bb4_and17_i_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i & 32'hFF)),
	.data_out(rnode_392to394_bb4_and17_i_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_392to394_bb4_and17_i_0_reg_394_fifo.DEPTH = 2;
defparam rnode_392to394_bb4_and17_i_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_392to394_bb4_and17_i_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to394_bb4_and17_i_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_392to394_bb4_and17_i_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i_stall_in_2 = 1'b0;
assign rnode_392to394_bb4_and17_i_0_NO_SHIFT_REG = rnode_392to394_bb4_and17_i_0_reg_394_NO_SHIFT_REG;
assign rnode_392to394_bb4_and17_i_0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_and17_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_var__u88_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4_var__u88_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4_var__u88_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_var__u88_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4_var__u88_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_var__u88_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_var__u88_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_var__u88_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_var__u88_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_var__u88_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_var__u88_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_var__u88_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_var__u88_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb4_var__u88),
	.data_out(rnode_392to393_bb4_var__u88_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_var__u88_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_var__u88_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4_var__u88_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_var__u88_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_var__u88_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u88_stall_in = 1'b0;
assign rnode_392to393_bb4_var__u88_0_NO_SHIFT_REG = rnode_392to393_bb4_var__u88_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_var__u88_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_var__u88_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_add192_i_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_add192_i_1_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_add192_i_2_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_add192_i_3_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_392to393_bb4_add192_i_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_valid_out_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_stall_in_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4_add192_i_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4_add192_i_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4_add192_i_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4_add192_i_0_stall_in_0_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4_add192_i_0_valid_out_0_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4_add192_i_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb4_add192_i),
	.data_out(rnode_392to393_bb4_add192_i_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4_add192_i_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4_add192_i_0_reg_393_fifo.DATA_WIDTH = 32;
defparam rnode_392to393_bb4_add192_i_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4_add192_i_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4_add192_i_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add192_i_stall_in = 1'b0;
assign rnode_392to393_bb4_add192_i_0_stall_in_0_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4_add192_i_0_NO_SHIFT_REG = rnode_392to393_bb4_add192_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4_add192_i_1_NO_SHIFT_REG = rnode_392to393_bb4_add192_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4_add192_i_2_NO_SHIFT_REG = rnode_392to393_bb4_add192_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4_add192_i_3_NO_SHIFT_REG = rnode_392to393_bb4_add192_i_0_reg_393_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_392to393_bb4__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_392to393_bb4__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_392to393_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_392to393_bb4__26_i_0_reg_393_inputs_ready_NO_SHIFT_REG;
 logic rnode_392to393_bb4__26_i_0_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__26_i_0_valid_out_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__26_i_0_stall_in_reg_393_NO_SHIFT_REG;
 logic rnode_392to393_bb4__26_i_0_stall_out_reg_393_NO_SHIFT_REG;

acl_data_fifo rnode_392to393_bb4__26_i_0_reg_393_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_392to393_bb4__26_i_0_reg_393_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_392to393_bb4__26_i_0_stall_in_reg_393_NO_SHIFT_REG),
	.valid_out(rnode_392to393_bb4__26_i_0_valid_out_reg_393_NO_SHIFT_REG),
	.stall_out(rnode_392to393_bb4__26_i_0_stall_out_reg_393_NO_SHIFT_REG),
	.data_in(local_bb4__26_i),
	.data_out(rnode_392to393_bb4__26_i_0_reg_393_NO_SHIFT_REG)
);

defparam rnode_392to393_bb4__26_i_0_reg_393_fifo.DEPTH = 1;
defparam rnode_392to393_bb4__26_i_0_reg_393_fifo.DATA_WIDTH = 1;
defparam rnode_392to393_bb4__26_i_0_reg_393_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_392to393_bb4__26_i_0_reg_393_fifo.IMPL = "shift_reg";

assign rnode_392to393_bb4__26_i_0_reg_393_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i_stall_in = 1'b0;
assign rnode_392to393_bb4__26_i_0_NO_SHIFT_REG = rnode_392to393_bb4__26_i_0_reg_393_NO_SHIFT_REG;
assign rnode_392to393_bb4__26_i_0_stall_in_reg_393_NO_SHIFT_REG = 1'b0;
assign rnode_392to393_bb4__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i15_stall_local;
wire local_bb4_cmp_i15;

assign local_bb4_cmp_i15 = ((local_bb4_shr_i12 & 32'h7FFF) > (local_bb4_shr3_i14 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i16_stall_local;
wire local_bb4_cmp8_i16;

assign local_bb4_cmp8_i16 = ((local_bb4_shr_i12 & 32'h7FFF) == (local_bb4_shr3_i14 & 32'h7FFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb4_var__u88_0_valid_out_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u88_0_stall_in_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u88_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u88_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u88_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u88_0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u88_0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_var__u88_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb4_var__u88_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb4_var__u88_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb4_var__u88_0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb4_var__u88_0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb4_var__u88_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in(rnode_392to393_bb4_var__u88_0_NO_SHIFT_REG),
	.data_out(rnode_393to394_bb4_var__u88_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb4_var__u88_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb4_var__u88_0_reg_394_fifo.DATA_WIDTH = 1;
defparam rnode_393to394_bb4_var__u88_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb4_var__u88_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb4_var__u88_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4_var__u88_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_var__u88_0_NO_SHIFT_REG = rnode_393to394_bb4_var__u88_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_var__u88_0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_var__u88_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and193_i_valid_out;
wire local_bb4_and193_i_stall_in;
wire local_bb4_and193_i_inputs_ready;
wire local_bb4_and193_i_stall_local;
wire [31:0] local_bb4_and193_i;

assign local_bb4_and193_i_inputs_ready = rnode_392to393_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and193_i = (rnode_392to393_bb4_add192_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and193_i_valid_out = 1'b1;
assign rnode_392to393_bb4_add192_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and195_i_valid_out;
wire local_bb4_and195_i_stall_in;
wire local_bb4_and195_i_inputs_ready;
wire local_bb4_and195_i_stall_local;
wire [31:0] local_bb4_and195_i;

assign local_bb4_and195_i_inputs_ready = rnode_392to393_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and195_i = (rnode_392to393_bb4_add192_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and195_i_valid_out = 1'b1;
assign rnode_392to393_bb4_add192_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and198_i_valid_out;
wire local_bb4_and198_i_stall_in;
wire local_bb4_and198_i_inputs_ready;
wire local_bb4_and198_i_stall_local;
wire [31:0] local_bb4_and198_i;

assign local_bb4_and198_i_inputs_ready = rnode_392to393_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and198_i = (rnode_392to393_bb4_add192_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and198_i_valid_out = 1'b1;
assign rnode_392to393_bb4_add192_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and201_i_stall_local;
wire [31:0] local_bb4_and201_i;

assign local_bb4_and201_i = (rnode_392to393_bb4_add192_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_393to395_bb4__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_393to395_bb4__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_393to395_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_393to395_bb4__26_i_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic rnode_393to395_bb4__26_i_0_reg_395_NO_SHIFT_REG;
 logic rnode_393to395_bb4__26_i_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_393to395_bb4__26_i_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_393to395_bb4__26_i_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_393to395_bb4__26_i_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to395_bb4__26_i_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to395_bb4__26_i_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_393to395_bb4__26_i_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_393to395_bb4__26_i_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(rnode_392to393_bb4__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_393to395_bb4__26_i_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_393to395_bb4__26_i_0_reg_395_fifo.DEPTH = 2;
defparam rnode_393to395_bb4__26_i_0_reg_395_fifo.DATA_WIDTH = 1;
defparam rnode_393to395_bb4__26_i_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to395_bb4__26_i_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_393to395_bb4__26_i_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_392to393_bb4__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_393to395_bb4__26_i_0_NO_SHIFT_REG = rnode_393to395_bb4__26_i_0_reg_395_NO_SHIFT_REG;
assign rnode_393to395_bb4__26_i_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_393to395_bb4__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4___i20_stall_local;
wire local_bb4___i20;

assign local_bb4___i20 = (local_bb4_cmp8_i16 & local_bb4_cmp13_i19);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_var__u88_0_valid_out_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u88_0_stall_in_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u88_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u88_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u88_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u88_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u88_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u88_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_var__u88_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_var__u88_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_var__u88_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_var__u88_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_var__u88_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(rnode_393to394_bb4_var__u88_0_NO_SHIFT_REG),
	.data_out(rnode_394to395_bb4_var__u88_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_var__u88_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_var__u88_0_reg_395_fifo.DATA_WIDTH = 1;
defparam rnode_394to395_bb4_var__u88_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_var__u88_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_var__u88_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_var__u88_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u88_0_NO_SHIFT_REG = rnode_394to395_bb4_var__u88_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_var__u88_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u88_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and193_i_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and193_i_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and193_i_2_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and193_i_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_valid_out_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_stall_in_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and193_i_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb4_and193_i_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb4_and193_i_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb4_and193_i_0_stall_in_0_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb4_and193_i_0_valid_out_0_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb4_and193_i_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in((local_bb4_and193_i & 32'hFFFFFFF)),
	.data_out(rnode_393to394_bb4_and193_i_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb4_and193_i_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb4_and193_i_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb4_and193_i_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb4_and193_i_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb4_and193_i_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and193_i_stall_in = 1'b0;
assign rnode_393to394_bb4_and193_i_0_stall_in_0_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_and193_i_0_NO_SHIFT_REG = rnode_393to394_bb4_and193_i_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_and193_i_1_NO_SHIFT_REG = rnode_393to394_bb4_and193_i_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4_and193_i_2_NO_SHIFT_REG = rnode_393to394_bb4_and193_i_0_reg_394_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb4_and195_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and195_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and195_i_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and195_i_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and195_i_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and195_i_0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and195_i_0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and195_i_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb4_and195_i_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb4_and195_i_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb4_and195_i_0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb4_and195_i_0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb4_and195_i_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in((local_bb4_and195_i & 32'h1F)),
	.data_out(rnode_393to394_bb4_and195_i_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb4_and195_i_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb4_and195_i_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb4_and195_i_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb4_and195_i_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb4_and195_i_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and195_i_stall_in = 1'b0;
assign rnode_393to394_bb4_and195_i_0_NO_SHIFT_REG = rnode_393to394_bb4_and195_i_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_and195_i_0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and195_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb4_and198_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and198_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and198_i_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and198_i_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4_and198_i_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and198_i_0_valid_out_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and198_i_0_stall_in_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4_and198_i_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb4_and198_i_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb4_and198_i_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb4_and198_i_0_stall_in_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb4_and198_i_0_valid_out_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb4_and198_i_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in((local_bb4_and198_i & 32'h1)),
	.data_out(rnode_393to394_bb4_and198_i_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb4_and198_i_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb4_and198_i_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb4_and198_i_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb4_and198_i_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb4_and198_i_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and198_i_stall_in = 1'b0;
assign rnode_393to394_bb4_and198_i_0_NO_SHIFT_REG = rnode_393to394_bb4_and198_i_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4_and198_i_0_stall_in_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and198_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i_stall_local;
wire [31:0] local_bb4_shr_i_i;

assign local_bb4_shr_i_i = ((local_bb4_and201_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4__26_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_valid_out_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_stall_in_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__26_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4__26_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4__26_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4__26_i_0_stall_in_0_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4__26_i_0_valid_out_0_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4__26_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(rnode_393to395_bb4__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_395to396_bb4__26_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4__26_i_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4__26_i_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_395to396_bb4__26_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4__26_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4__26_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_393to395_bb4__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__26_i_0_stall_in_0_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__26_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__26_i_0_NO_SHIFT_REG = rnode_395to396_bb4__26_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4__26_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__26_i_1_NO_SHIFT_REG = rnode_395to396_bb4__26_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4__26_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__26_i_2_NO_SHIFT_REG = rnode_395to396_bb4__26_i_0_reg_396_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u53_valid_out_2;
wire local_bb4_var__u53_stall_in_2;
wire local_bb4__21_i21_valid_out;
wire local_bb4__21_i21_stall_in;
wire local_bb4__21_i21_inputs_ready;
wire local_bb4__21_i21_stall_local;
wire local_bb4__21_i21;

assign local_bb4__21_i21_inputs_ready = (rnode_393to394_bb4_t_313_pop8_c1_ene4_0_valid_out_0_NO_SHIFT_REG & rnode_393to394_bb4_var__u96_0_valid_out_1_NO_SHIFT_REG & rnode_393to394_bb4_var__u96_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__21_i21 = (local_bb4_cmp_i15 | local_bb4___i20);
assign local_bb4_var__u53_valid_out_2 = 1'b1;
assign local_bb4__21_i21_valid_out = 1'b1;
assign rnode_393to394_bb4_t_313_pop8_c1_ene4_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_var__u96_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_var__u96_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr216_i_stall_local;
wire [31:0] local_bb4_shr216_i;

assign local_bb4_shr216_i = ((rnode_393to394_bb4_and193_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i_stall_local;
wire [31:0] local_bb4__pre_i;

assign local_bb4__pre_i = ((rnode_393to394_bb4_and195_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i_stall_local;
wire [31:0] local_bb4_or_i_i;

assign local_bb4_or_i_i = ((local_bb4_shr_i_i & 32'h3FFFFFF) | (local_bb4_and201_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond292_i_stall_local;
wire [31:0] local_bb4_cond292_i;

assign local_bb4_cond292_i = (rnode_395to396_bb4__26_i_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u97_stall_local;
wire [31:0] local_bb4_var__u97;

assign local_bb4_var__u97[31:1] = 31'h0;
assign local_bb4_var__u97[0] = rnode_395to396_bb4__26_i_2_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_var__u53_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u53_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_var__u53_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u53_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u53_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_var__u53_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u53_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_var__u53_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u53_0_valid_out_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u53_0_stall_in_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_var__u53_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_var__u53_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_var__u53_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_var__u53_0_stall_in_0_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_var__u53_0_valid_out_0_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_var__u53_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(local_bb4_var__u53),
	.data_out(rnode_394to395_bb4_var__u53_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_var__u53_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_var__u53_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_394to395_bb4_var__u53_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_var__u53_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_var__u53_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u53_stall_in_2 = 1'b0;
assign rnode_394to395_bb4_var__u53_0_stall_in_0_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u53_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4_var__u53_0_NO_SHIFT_REG = rnode_394to395_bb4_var__u53_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_var__u53_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4_var__u53_1_NO_SHIFT_REG = rnode_394to395_bb4_var__u53_0_reg_395_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4__21_i21_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_valid_out_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_stall_in_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4__21_i21_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4__21_i21_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4__21_i21_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4__21_i21_0_stall_in_0_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4__21_i21_0_valid_out_0_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4__21_i21_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(local_bb4__21_i21),
	.data_out(rnode_394to395_bb4__21_i21_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4__21_i21_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4__21_i21_0_reg_395_fifo.DATA_WIDTH = 1;
defparam rnode_394to395_bb4__21_i21_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4__21_i21_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4__21_i21_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i21_stall_in = 1'b0;
assign rnode_394to395_bb4__21_i21_0_stall_in_0_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4__21_i21_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4__21_i21_0_NO_SHIFT_REG = rnode_394to395_bb4__21_i21_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4__21_i21_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4__21_i21_1_NO_SHIFT_REG = rnode_394to395_bb4__21_i21_0_reg_395_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or219_i_stall_local;
wire [31:0] local_bb4_or219_i;

assign local_bb4_or219_i = ((local_bb4_shr216_i & 32'h7FFFFFF) | (rnode_393to394_bb4_and198_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool213_i_stall_local;
wire local_bb4_tobool213_i;

assign local_bb4_tobool213_i = ((local_bb4__pre_i & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i_stall_local;
wire [31:0] local_bb4_shr1_i_i;

assign local_bb4_shr1_i_i = ((local_bb4_or_i_i & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i_stall_local;
wire [31:0] local_bb4_lnot_ext_i;

assign local_bb4_lnot_ext_i = ((local_bb4_var__u97 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i22_stall_local;
wire [31:0] local_bb4__22_i22;

assign local_bb4__22_i22 = (rnode_394to395_bb4__21_i21_0_NO_SHIFT_REG ? rnode_394to395_bb4_var__u53_0_NO_SHIFT_REG : rnode_394to395_bb4_var__u96_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i23_stall_local;
wire [31:0] local_bb4__23_i23;

assign local_bb4__23_i23 = (rnode_394to395_bb4__21_i21_1_NO_SHIFT_REG ? rnode_394to395_bb4_var__u96_1_NO_SHIFT_REG : rnode_394to395_bb4_var__u53_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i_stall_local;
wire local_bb4__40_demorgan_i;

assign local_bb4__40_demorgan_i = (rnode_392to394_bb4_cmp37_i_0_NO_SHIFT_REG | local_bb4_tobool213_i);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i_stall_local;
wire local_bb4__42_i;

assign local_bb4__42_i = (local_bb4_tobool213_i & local_bb4_not_cmp37_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i_stall_local;
wire [31:0] local_bb4_or2_i_i;

assign local_bb4_or2_i_i = ((local_bb4_shr1_i_i & 32'h1FFFFFF) | (local_bb4_or_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i26_stall_local;
wire [31:0] local_bb4_shr18_i26;

assign local_bb4_shr18_i26 = (local_bb4__22_i22 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i24_stall_local;
wire [31:0] local_bb4_shr16_i24;

assign local_bb4_shr16_i24 = (local_bb4__23_i23 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4__43_i_stall_local;
wire [31:0] local_bb4__43_i;

assign local_bb4__43_i = (local_bb4__42_i ? 32'h0 : (local_bb4__pre_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i_stall_local;
wire [31:0] local_bb4_shr3_i_i;

assign local_bb4_shr3_i_i = ((local_bb4_or2_i_i & 32'h7FFFFFF) >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i27_stall_local;
wire [31:0] local_bb4_and19_i27;

assign local_bb4_and19_i27 = ((local_bb4_shr18_i26 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i56_stall_local;
wire [31:0] local_bb4_sub_i56;

assign local_bb4_sub_i56 = ((local_bb4_shr16_i24 & 32'h1FF) - (local_bb4_shr18_i26 & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i_stall_local;
wire [31:0] local_bb4_or4_i_i;

assign local_bb4_or4_i_i = ((local_bb4_shr3_i_i & 32'h7FFFFF) | (local_bb4_or2_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i31_stall_local;
wire local_bb4_lnot23_i31;

assign local_bb4_lnot23_i31 = ((local_bb4_and19_i27 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i33_stall_local;
wire local_bb4_cmp27_i33;

assign local_bb4_cmp27_i33 = ((local_bb4_and19_i27 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and68_i57_stall_local;
wire [31:0] local_bb4_and68_i57;

assign local_bb4_and68_i57 = (local_bb4_sub_i56 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i_stall_local;
wire [31:0] local_bb4_shr5_i_i;

assign local_bb4_shr5_i_i = ((local_bb4_or4_i_i & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp69_i58_stall_local;
wire local_bb4_cmp69_i58;

assign local_bb4_cmp69_i58 = ((local_bb4_and68_i57 & 32'hFF) > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i_stall_local;
wire [31:0] local_bb4_or6_i_i;

assign local_bb4_or6_i_i = ((local_bb4_shr5_i_i & 32'h7FFFF) | (local_bb4_or4_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__22_i22_valid_out_1;
wire local_bb4__22_i22_stall_in_1;
wire local_bb4__23_i23_valid_out_1;
wire local_bb4__23_i23_stall_in_1;
wire local_bb4_shr16_i24_valid_out_1;
wire local_bb4_shr16_i24_stall_in_1;
wire local_bb4_lnot23_i31_valid_out;
wire local_bb4_lnot23_i31_stall_in;
wire local_bb4_cmp27_i33_valid_out;
wire local_bb4_cmp27_i33_stall_in;
wire local_bb4_align_0_i59_valid_out;
wire local_bb4_align_0_i59_stall_in;
wire local_bb4_align_0_i59_inputs_ready;
wire local_bb4_align_0_i59_stall_local;
wire [31:0] local_bb4_align_0_i59;

assign local_bb4_align_0_i59_inputs_ready = (rnode_394to395_bb4__21_i21_0_valid_out_0_NO_SHIFT_REG & rnode_394to395_bb4_var__u53_0_valid_out_0_NO_SHIFT_REG & rnode_394to395_bb4_var__u96_0_valid_out_0_NO_SHIFT_REG & rnode_394to395_bb4__21_i21_0_valid_out_1_NO_SHIFT_REG & rnode_394to395_bb4_var__u53_0_valid_out_1_NO_SHIFT_REG & rnode_394to395_bb4_var__u96_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_align_0_i59 = (local_bb4_cmp69_i58 ? 32'h1F : (local_bb4_and68_i57 & 32'hFF));
assign local_bb4__22_i22_valid_out_1 = 1'b1;
assign local_bb4__23_i23_valid_out_1 = 1'b1;
assign local_bb4_shr16_i24_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i31_valid_out = 1'b1;
assign local_bb4_cmp27_i33_valid_out = 1'b1;
assign local_bb4_align_0_i59_valid_out = 1'b1;
assign rnode_394to395_bb4__21_i21_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u53_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u96_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4__21_i21_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u53_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u96_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i_stall_local;
wire [31:0] local_bb4_shr7_i_i;

assign local_bb4_shr7_i_i = ((local_bb4_or6_i_i & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i_stall_local;
wire [31:0] local_bb4_or6_masked_i_i;

assign local_bb4_or6_masked_i_i = ((local_bb4_or6_i_i & 32'h7FFFFFF) & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4__22_i22_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__22_i22_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4__22_i22_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__22_i22_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__22_i22_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4__22_i22_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__22_i22_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4__22_i22_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__22_i22_0_valid_out_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__22_i22_0_stall_in_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__22_i22_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4__22_i22_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4__22_i22_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4__22_i22_0_stall_in_0_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4__22_i22_0_valid_out_0_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4__22_i22_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(local_bb4__22_i22),
	.data_out(rnode_395to396_bb4__22_i22_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4__22_i22_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4__22_i22_0_reg_396_fifo.DATA_WIDTH = 32;
defparam rnode_395to396_bb4__22_i22_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4__22_i22_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4__22_i22_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i22_stall_in_1 = 1'b0;
assign rnode_395to396_bb4__22_i22_0_stall_in_0_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__22_i22_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__22_i22_0_NO_SHIFT_REG = rnode_395to396_bb4__22_i22_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4__22_i22_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__22_i22_1_NO_SHIFT_REG = rnode_395to396_bb4__22_i22_0_reg_396_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4__23_i23_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4__23_i23_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4__23_i23_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4__23_i23_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4__23_i23_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_valid_out_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_stall_in_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__23_i23_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4__23_i23_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4__23_i23_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4__23_i23_0_stall_in_0_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4__23_i23_0_valid_out_0_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4__23_i23_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(local_bb4__23_i23),
	.data_out(rnode_395to396_bb4__23_i23_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4__23_i23_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4__23_i23_0_reg_396_fifo.DATA_WIDTH = 32;
defparam rnode_395to396_bb4__23_i23_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4__23_i23_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4__23_i23_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i23_stall_in_1 = 1'b0;
assign rnode_395to396_bb4__23_i23_0_stall_in_0_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__23_i23_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__23_i23_0_NO_SHIFT_REG = rnode_395to396_bb4__23_i23_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4__23_i23_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__23_i23_1_NO_SHIFT_REG = rnode_395to396_bb4__23_i23_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4__23_i23_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__23_i23_2_NO_SHIFT_REG = rnode_395to396_bb4__23_i23_0_reg_396_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_395to397_bb4_shr16_i24_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to397_bb4_shr16_i24_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_395to397_bb4_shr16_i24_0_NO_SHIFT_REG;
 logic rnode_395to397_bb4_shr16_i24_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to397_bb4_shr16_i24_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_395to397_bb4_shr16_i24_1_NO_SHIFT_REG;
 logic rnode_395to397_bb4_shr16_i24_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to397_bb4_shr16_i24_0_reg_397_NO_SHIFT_REG;
 logic rnode_395to397_bb4_shr16_i24_0_valid_out_0_reg_397_NO_SHIFT_REG;
 logic rnode_395to397_bb4_shr16_i24_0_stall_in_0_reg_397_NO_SHIFT_REG;
 logic rnode_395to397_bb4_shr16_i24_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_395to397_bb4_shr16_i24_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to397_bb4_shr16_i24_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to397_bb4_shr16_i24_0_stall_in_0_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_395to397_bb4_shr16_i24_0_valid_out_0_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_395to397_bb4_shr16_i24_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i24 & 32'h1FF)),
	.data_out(rnode_395to397_bb4_shr16_i24_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_395to397_bb4_shr16_i24_0_reg_397_fifo.DEPTH = 2;
defparam rnode_395to397_bb4_shr16_i24_0_reg_397_fifo.DATA_WIDTH = 32;
defparam rnode_395to397_bb4_shr16_i24_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to397_bb4_shr16_i24_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_395to397_bb4_shr16_i24_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i24_stall_in_1 = 1'b0;
assign rnode_395to397_bb4_shr16_i24_0_stall_in_0_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_395to397_bb4_shr16_i24_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to397_bb4_shr16_i24_0_NO_SHIFT_REG = rnode_395to397_bb4_shr16_i24_0_reg_397_NO_SHIFT_REG;
assign rnode_395to397_bb4_shr16_i24_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to397_bb4_shr16_i24_1_NO_SHIFT_REG = rnode_395to397_bb4_shr16_i24_0_reg_397_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_lnot23_i31_0_valid_out_NO_SHIFT_REG;
 logic rnode_395to396_bb4_lnot23_i31_0_stall_in_NO_SHIFT_REG;
 logic rnode_395to396_bb4_lnot23_i31_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_lnot23_i31_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to396_bb4_lnot23_i31_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_lnot23_i31_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_lnot23_i31_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_lnot23_i31_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_lnot23_i31_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_lnot23_i31_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_lnot23_i31_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_lnot23_i31_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_lnot23_i31_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i31),
	.data_out(rnode_395to396_bb4_lnot23_i31_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_lnot23_i31_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_lnot23_i31_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_395to396_bb4_lnot23_i31_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_lnot23_i31_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_lnot23_i31_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i31_stall_in = 1'b0;
assign rnode_395to396_bb4_lnot23_i31_0_NO_SHIFT_REG = rnode_395to396_bb4_lnot23_i31_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_lnot23_i31_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_lnot23_i31_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_395to397_bb4_cmp27_i33_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_1_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_2_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_reg_397_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_valid_out_0_reg_397_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_stall_in_0_reg_397_NO_SHIFT_REG;
 logic rnode_395to397_bb4_cmp27_i33_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_395to397_bb4_cmp27_i33_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to397_bb4_cmp27_i33_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to397_bb4_cmp27_i33_0_stall_in_0_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_395to397_bb4_cmp27_i33_0_valid_out_0_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_395to397_bb4_cmp27_i33_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i33),
	.data_out(rnode_395to397_bb4_cmp27_i33_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_395to397_bb4_cmp27_i33_0_reg_397_fifo.DEPTH = 2;
defparam rnode_395to397_bb4_cmp27_i33_0_reg_397_fifo.DATA_WIDTH = 1;
defparam rnode_395to397_bb4_cmp27_i33_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to397_bb4_cmp27_i33_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_395to397_bb4_cmp27_i33_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i33_stall_in = 1'b0;
assign rnode_395to397_bb4_cmp27_i33_0_stall_in_0_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_395to397_bb4_cmp27_i33_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to397_bb4_cmp27_i33_0_NO_SHIFT_REG = rnode_395to397_bb4_cmp27_i33_0_reg_397_NO_SHIFT_REG;
assign rnode_395to397_bb4_cmp27_i33_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to397_bb4_cmp27_i33_1_NO_SHIFT_REG = rnode_395to397_bb4_cmp27_i33_0_reg_397_NO_SHIFT_REG;
assign rnode_395to397_bb4_cmp27_i33_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_395to397_bb4_cmp27_i33_2_NO_SHIFT_REG = rnode_395to397_bb4_cmp27_i33_0_reg_397_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_align_0_i59_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_align_0_i59_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_align_0_i59_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_align_0_i59_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_align_0_i59_3_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_align_0_i59_4_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_align_0_i59_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_valid_out_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_stall_in_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_align_0_i59_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_align_0_i59_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_align_0_i59_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_align_0_i59_0_stall_in_0_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_align_0_i59_0_valid_out_0_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_align_0_i59_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in((local_bb4_align_0_i59 & 32'hFF)),
	.data_out(rnode_395to396_bb4_align_0_i59_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_align_0_i59_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_align_0_i59_0_reg_396_fifo.DATA_WIDTH = 32;
defparam rnode_395to396_bb4_align_0_i59_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_align_0_i59_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_align_0_i59_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_align_0_i59_stall_in = 1'b0;
assign rnode_395to396_bb4_align_0_i59_0_stall_in_0_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_align_0_i59_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_align_0_i59_0_NO_SHIFT_REG = rnode_395to396_bb4_align_0_i59_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_align_0_i59_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_align_0_i59_1_NO_SHIFT_REG = rnode_395to396_bb4_align_0_i59_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_align_0_i59_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_align_0_i59_2_NO_SHIFT_REG = rnode_395to396_bb4_align_0_i59_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_align_0_i59_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_align_0_i59_3_NO_SHIFT_REG = rnode_395to396_bb4_align_0_i59_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_align_0_i59_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_align_0_i59_4_NO_SHIFT_REG = rnode_395to396_bb4_align_0_i59_0_reg_396_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i_stall_local;
wire [31:0] local_bb4_neg_i_i;

assign local_bb4_neg_i_i = ((local_bb4_or6_masked_i_i & 32'h7FFFFFF) | (local_bb4_shr7_i_i & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i29_stall_local;
wire [31:0] local_bb4_and21_i29;

assign local_bb4_and21_i29 = (rnode_395to396_bb4__22_i22_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i28_valid_out;
wire local_bb4_and20_i28_stall_in;
wire local_bb4_and20_i28_inputs_ready;
wire local_bb4_and20_i28_stall_local;
wire [31:0] local_bb4_and20_i28;

assign local_bb4_and20_i28_inputs_ready = rnode_395to396_bb4__23_i23_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i28 = (rnode_395to396_bb4__23_i23_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i28_valid_out = 1'b1;
assign rnode_395to396_bb4__23_i23_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i34_valid_out;
wire local_bb4_and35_i34_stall_in;
wire local_bb4_and35_i34_inputs_ready;
wire local_bb4_and35_i34_stall_local;
wire [31:0] local_bb4_and35_i34;

assign local_bb4_and35_i34_inputs_ready = rnode_395to396_bb4__23_i23_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i34 = (rnode_395to396_bb4__23_i23_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i34_valid_out = 1'b1;
assign rnode_395to396_bb4__23_i23_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i35_stall_local;
wire [31:0] local_bb4_xor_i35;

assign local_bb4_xor_i35 = (rnode_395to396_bb4__23_i23_2_NO_SHIFT_REG ^ rnode_395to396_bb4__22_i22_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i25_stall_local;
wire [31:0] local_bb4_and17_i25;

assign local_bb4_and17_i25 = ((rnode_395to397_bb4_shr16_i24_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_397to399_bb4_shr16_i24_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to399_bb4_shr16_i24_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_397to399_bb4_shr16_i24_0_NO_SHIFT_REG;
 logic rnode_397to399_bb4_shr16_i24_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_397to399_bb4_shr16_i24_0_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_shr16_i24_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_shr16_i24_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_shr16_i24_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_397to399_bb4_shr16_i24_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to399_bb4_shr16_i24_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to399_bb4_shr16_i24_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_397to399_bb4_shr16_i24_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_397to399_bb4_shr16_i24_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in((rnode_395to397_bb4_shr16_i24_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_397to399_bb4_shr16_i24_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_397to399_bb4_shr16_i24_0_reg_399_fifo.DEPTH = 2;
defparam rnode_397to399_bb4_shr16_i24_0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_397to399_bb4_shr16_i24_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to399_bb4_shr16_i24_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_397to399_bb4_shr16_i24_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_395to397_bb4_shr16_i24_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_shr16_i24_0_NO_SHIFT_REG = rnode_397to399_bb4_shr16_i24_0_reg_399_NO_SHIFT_REG;
assign rnode_397to399_bb4_shr16_i24_0_stall_in_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_shr16_i24_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and93_i67_stall_local;
wire [31:0] local_bb4_and93_i67;

assign local_bb4_and93_i67 = ((rnode_395to396_bb4_align_0_i59_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and95_i69_stall_local;
wire [31:0] local_bb4_and95_i69;

assign local_bb4_and95_i69 = ((rnode_395to396_bb4_align_0_i59_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and115_i85_stall_local;
wire [31:0] local_bb4_and115_i85;

assign local_bb4_and115_i85 = ((rnode_395to396_bb4_align_0_i59_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and130_i91_stall_local;
wire [31:0] local_bb4_and130_i91;

assign local_bb4_and130_i91 = ((rnode_395to396_bb4_align_0_i59_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and149_i96_stall_local;
wire [31:0] local_bb4_and149_i96;

assign local_bb4_and149_i96 = ((rnode_395to396_bb4_align_0_i59_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i9_stall_local;
wire [31:0] local_bb4_and_i_i9;

assign local_bb4_and_i_i9 = ((local_bb4_neg_i_i & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i40_stall_local;
wire local_bb4_lnot33_not_i40;

assign local_bb4_lnot33_not_i40 = ((local_bb4_and21_i29 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or64_i53_stall_local;
wire [31:0] local_bb4_or64_i53;

assign local_bb4_or64_i53 = ((local_bb4_and21_i29 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_and20_i28_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and20_i28_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_and20_i28_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and20_i28_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and20_i28_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_and20_i28_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and20_i28_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_and20_i28_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and20_i28_0_valid_out_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and20_i28_0_stall_in_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and20_i28_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_and20_i28_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_and20_i28_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_and20_i28_0_stall_in_0_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_and20_i28_0_valid_out_0_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_and20_i28_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i28 & 32'h7FFFFF)),
	.data_out(rnode_396to397_bb4_and20_i28_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_and20_i28_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_and20_i28_0_reg_397_fifo.DATA_WIDTH = 32;
defparam rnode_396to397_bb4_and20_i28_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_and20_i28_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_and20_i28_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i28_stall_in = 1'b0;
assign rnode_396to397_bb4_and20_i28_0_stall_in_0_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_and20_i28_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_and20_i28_0_NO_SHIFT_REG = rnode_396to397_bb4_and20_i28_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_and20_i28_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_and20_i28_1_NO_SHIFT_REG = rnode_396to397_bb4_and20_i28_0_reg_397_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_and35_i34_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and35_i34_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_and35_i34_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and35_i34_0_valid_out_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and35_i34_0_stall_in_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and35_i34_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_and35_i34_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_and35_i34_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_and35_i34_0_stall_in_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_and35_i34_0_valid_out_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_and35_i34_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i34 & 32'h80000000)),
	.data_out(rnode_396to397_bb4_and35_i34_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_and35_i34_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_and35_i34_0_reg_397_fifo.DATA_WIDTH = 32;
defparam rnode_396to397_bb4_and35_i34_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_and35_i34_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_and35_i34_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i34_stall_in = 1'b0;
assign rnode_396to397_bb4_and35_i34_0_NO_SHIFT_REG = rnode_396to397_bb4_and35_i34_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_and35_i34_0_stall_in_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp37_i36_stall_local;
wire local_bb4_cmp37_i36;

assign local_bb4_cmp37_i36 = ($signed(local_bb4_xor_i35) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor_lobit_i109_stall_local;
wire [31:0] local_bb4_xor_lobit_i109;

assign local_bb4_xor_lobit_i109 = ($signed(local_bb4_xor_i35) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and36_lobit_i111_stall_local;
wire [31:0] local_bb4_and36_lobit_i111;

assign local_bb4_and36_lobit_i111 = (local_bb4_xor_i35 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i30_stall_local;
wire local_bb4_lnot_i30;

assign local_bb4_lnot_i30 = ((local_bb4_and17_i25 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i32_stall_local;
wire local_bb4_cmp25_i32;

assign local_bb4_cmp25_i32 = ((local_bb4_and17_i25 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp96_i70_stall_local;
wire local_bb4_cmp96_i70;

assign local_bb4_cmp96_i70 = ((local_bb4_and95_i69 & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp116_i86_stall_local;
wire local_bb4_cmp116_i86;

assign local_bb4_cmp116_i86 = ((local_bb4_and115_i85 & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp131_not_i93_stall_local;
wire local_bb4_cmp131_not_i93;

assign local_bb4_cmp131_not_i93 = ((local_bb4_and130_i91 & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i98_stall_local;
wire local_bb4_Pivot20_i98;

assign local_bb4_Pivot20_i98 = ((local_bb4_and149_i96 & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i99_stall_local;
wire local_bb4_SwitchLeaf_i99;

assign local_bb4_SwitchLeaf_i99 = ((local_bb4_and149_i96 & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i9_valid_out;
wire local_bb4__and_i_i9_stall_in;
wire local_bb4__and_i_i9_inputs_ready;
wire local_bb4__and_i_i9_stall_local;
wire [31:0] local_bb4__and_i_i9;

thirtysix_six_comp local_bb4__and_i_i9_popcnt_instance (
	.data((local_bb4_and_i_i9 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i9)
);


assign local_bb4__and_i_i9_inputs_ready = rnode_392to393_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i9_valid_out = 1'b1;
assign rnode_392to393_bb4_add192_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shl65_i54_stall_local;
wire [31:0] local_bb4_shl65_i54;

assign local_bb4_shl65_i54 = ((local_bb4_or64_i53 & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i38_stall_local;
wire local_bb4_lnot30_i38;

assign local_bb4_lnot30_i38 = ((rnode_396to397_bb4_and20_i28_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i50_stall_local;
wire [31:0] local_bb4_or_i50;

assign local_bb4_or_i50 = ((rnode_396to397_bb4_and20_i28_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_397to399_bb4_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_397to399_bb4_and35_i34_0_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and35_i34_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_397to399_bb4_and35_i34_0_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and35_i34_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and35_i34_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and35_i34_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_397to399_bb4_and35_i34_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to399_bb4_and35_i34_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to399_bb4_and35_i34_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_397to399_bb4_and35_i34_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_397to399_bb4_and35_i34_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in((rnode_396to397_bb4_and35_i34_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_397to399_bb4_and35_i34_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_397to399_bb4_and35_i34_0_reg_399_fifo.DEPTH = 2;
defparam rnode_397to399_bb4_and35_i34_0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_397to399_bb4_and35_i34_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to399_bb4_and35_i34_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_397to399_bb4_and35_i34_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_and35_i34_0_NO_SHIFT_REG = rnode_397to399_bb4_and35_i34_0_reg_399_NO_SHIFT_REG;
assign rnode_397to399_bb4_and35_i34_0_stall_in_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i37_stall_local;
wire local_bb4_cmp25_not_i37;

assign local_bb4_cmp25_not_i37 = (local_bb4_cmp25_i32 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u98_stall_local;
wire local_bb4_var__u98;

assign local_bb4_var__u98 = (local_bb4_cmp25_i32 | rnode_395to397_bb4_cmp27_i33_2_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_393to394_bb4__and_i_i9_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4__and_i_i9_0_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4__and_i_i9_1_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4__and_i_i9_2_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_reg_394_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_393to394_bb4__and_i_i9_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_valid_out_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_stall_in_0_reg_394_NO_SHIFT_REG;
 logic rnode_393to394_bb4__and_i_i9_0_stall_out_reg_394_NO_SHIFT_REG;

acl_data_fifo rnode_393to394_bb4__and_i_i9_0_reg_394_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_393to394_bb4__and_i_i9_0_reg_394_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_393to394_bb4__and_i_i9_0_stall_in_0_reg_394_NO_SHIFT_REG),
	.valid_out(rnode_393to394_bb4__and_i_i9_0_valid_out_0_reg_394_NO_SHIFT_REG),
	.stall_out(rnode_393to394_bb4__and_i_i9_0_stall_out_reg_394_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i9 & 32'h3F)),
	.data_out(rnode_393to394_bb4__and_i_i9_0_reg_394_NO_SHIFT_REG)
);

defparam rnode_393to394_bb4__and_i_i9_0_reg_394_fifo.DEPTH = 1;
defparam rnode_393to394_bb4__and_i_i9_0_reg_394_fifo.DATA_WIDTH = 32;
defparam rnode_393to394_bb4__and_i_i9_0_reg_394_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_393to394_bb4__and_i_i9_0_reg_394_fifo.IMPL = "shift_reg";

assign rnode_393to394_bb4__and_i_i9_0_reg_394_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i9_stall_in = 1'b0;
assign rnode_393to394_bb4__and_i_i9_0_stall_in_0_reg_394_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4__and_i_i9_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4__and_i_i9_0_NO_SHIFT_REG = rnode_393to394_bb4__and_i_i9_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4__and_i_i9_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4__and_i_i9_1_NO_SHIFT_REG = rnode_393to394_bb4__and_i_i9_0_reg_394_NO_SHIFT_REG;
assign rnode_393to394_bb4__and_i_i9_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_393to394_bb4__and_i_i9_2_NO_SHIFT_REG = rnode_393to394_bb4__and_i_i9_0_reg_394_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__28_i55_stall_local;
wire [31:0] local_bb4__28_i55;

assign local_bb4__28_i55 = (rnode_395to396_bb4_lnot23_i31_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl65_i54 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i42_stall_local;
wire local_bb4_lnot30_not_i42;

assign local_bb4_lnot30_not_i42 = (local_bb4_lnot30_i38 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i51_stall_local;
wire [31:0] local_bb4_shl_i51;

assign local_bb4_shl_i51 = ((local_bb4_or_i50 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_399to400_bb4_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4_and35_i34_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and35_i34_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4_and35_i34_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and35_i34_0_valid_out_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and35_i34_0_stall_in_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and35_i34_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_399to400_bb4_and35_i34_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to400_bb4_and35_i34_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to400_bb4_and35_i34_0_stall_in_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_399to400_bb4_and35_i34_0_valid_out_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_399to400_bb4_and35_i34_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in((rnode_397to399_bb4_and35_i34_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_399to400_bb4_and35_i34_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_399to400_bb4_and35_i34_0_reg_400_fifo.DEPTH = 1;
defparam rnode_399to400_bb4_and35_i34_0_reg_400_fifo.DATA_WIDTH = 32;
defparam rnode_399to400_bb4_and35_i34_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to400_bb4_and35_i34_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_399to400_bb4_and35_i34_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_397to399_bb4_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_and35_i34_0_NO_SHIFT_REG = rnode_399to400_bb4_and35_i34_0_reg_400_NO_SHIFT_REG;
assign rnode_399to400_bb4_and35_i34_0_stall_in_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i39_stall_local;
wire local_bb4_or_cond_i39;

assign local_bb4_or_cond_i39 = (local_bb4_lnot30_i38 | local_bb4_cmp25_not_i37);

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i_stall_local;
wire [31:0] local_bb4_and9_i_i;

assign local_bb4_and9_i_i = ((rnode_393to394_bb4__and_i_i9_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and203_i_stall_local;
wire [31:0] local_bb4_and203_i;

assign local_bb4_and203_i = ((rnode_393to394_bb4__and_i_i9_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i_stall_local;
wire [31:0] local_bb4_and206_i;

assign local_bb4_and206_i = ((rnode_393to394_bb4__and_i_i9_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_and72_i60_stall_local;
wire [31:0] local_bb4_and72_i60;

assign local_bb4_and72_i60 = ((local_bb4__28_i55 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i63_stall_local;
wire [31:0] local_bb4_and75_i63;

assign local_bb4_and75_i63 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and78_i65_stall_local;
wire [31:0] local_bb4_and78_i65;

assign local_bb4_and78_i65 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr94_i68_stall_local;
wire [31:0] local_bb4_shr94_i68;

assign local_bb4_shr94_i68 = ((local_bb4__28_i55 & 32'h7FFFFF8) >> (local_bb4_and93_i67 & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i71_stall_local;
wire [31:0] local_bb4_and90_i71;

assign local_bb4_and90_i71 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and87_i72_stall_local;
wire [31:0] local_bb4_and87_i72;

assign local_bb4_and87_i72 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and84_i73_stall_local;
wire [31:0] local_bb4_and84_i73;

assign local_bb4_and84_i73 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u99_stall_local;
wire [31:0] local_bb4_var__u99;

assign local_bb4_var__u99 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i43_stall_local;
wire local_bb4_or_cond_not_i43;

assign local_bb4_or_cond_not_i43 = (local_bb4_cmp25_i32 & local_bb4_lnot30_not_i42);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i52_stall_local;
wire [31:0] local_bb4__27_i52;

assign local_bb4__27_i52 = (local_bb4_lnot_i30 ? 32'h0 : ((local_bb4_shl_i51 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i47_stall_local;
wire local_bb4_reduction_8_i47;

assign local_bb4_reduction_8_i47 = (rnode_395to397_bb4_cmp27_i33_1_NO_SHIFT_REG & local_bb4_or_cond_i39);

// This section implements an unregistered operation.
// 
wire local_bb4_sub239_i_stall_local;
wire [31:0] local_bb4_sub239_i;

assign local_bb4_sub239_i = (32'h0 - (local_bb4_and9_i_i & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl204_i_stall_local;
wire [31:0] local_bb4_shl204_i;

assign local_bb4_shl204_i = ((rnode_393to394_bb4_and193_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and203_i & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb4_and72_tr_i61_stall_local;
wire [7:0] local_bb4_and72_tr_i61;
wire [31:0] local_bb4_and72_tr_i61$ps;

assign local_bb4_and72_tr_i61$ps = (local_bb4_and72_i60 & 32'hFFFFFF);
assign local_bb4_and72_tr_i61 = local_bb4_and72_tr_i61$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp76_i64_stall_local;
wire local_bb4_cmp76_i64;

assign local_bb4_cmp76_i64 = ((local_bb4_and75_i63 & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp79_i66_stall_local;
wire local_bb4_cmp79_i66;

assign local_bb4_cmp79_i66 = ((local_bb4_and78_i65 & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and142_i95_stall_local;
wire [31:0] local_bb4_and142_i95;

assign local_bb4_and142_i95 = (local_bb4_shr94_i68 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr150_i97_stall_local;
wire [31:0] local_bb4_shr150_i97;

assign local_bb4_shr150_i97 = (local_bb4_shr94_i68 >> (local_bb4_and149_i96 & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u100_stall_local;
wire [31:0] local_bb4_var__u100;

assign local_bb4_var__u100 = (local_bb4_shr94_i68 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and146_i100_stall_local;
wire [31:0] local_bb4_and146_i100;

assign local_bb4_and146_i100 = (local_bb4_shr94_i68 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i74_stall_local;
wire local_bb4_cmp91_i74;

assign local_bb4_cmp91_i74 = ((local_bb4_and90_i71 & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp88_i75_stall_local;
wire local_bb4_cmp88_i75;

assign local_bb4_cmp88_i75 = ((local_bb4_and87_i72 & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp85_i76_stall_local;
wire local_bb4_cmp85_i76;

assign local_bb4_cmp85_i76 = ((local_bb4_and84_i73 & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u101_stall_local;
wire local_bb4_var__u101;

assign local_bb4_var__u101 = ((local_bb4_var__u99 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cond244_i_stall_local;
wire [31:0] local_bb4_cond244_i;

assign local_bb4_cond244_i = (rnode_392to394_bb4_cmp37_i_2_NO_SHIFT_REG ? local_bb4_sub239_i : (local_bb4__43_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and205_i_stall_local;
wire [31:0] local_bb4_and205_i;

assign local_bb4_and205_i = (local_bb4_shl204_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool74_i62_stall_local;
wire [7:0] local_bb4_frombool74_i62;

assign local_bb4_frombool74_i62 = (local_bb4_and72_tr_i61 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u102_stall_local;
wire [31:0] local_bb4_var__u102;

assign local_bb4_var__u102 = ((local_bb4_and146_i100 & 32'h3FFFFFFF) | local_bb4_shr94_i68);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i82_stall_local;
wire local_bb4__31_v_i82;

assign local_bb4__31_v_i82 = (local_bb4_cmp96_i70 ? local_bb4_cmp79_i66 : local_bb4_cmp91_i74);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i80_stall_local;
wire local_bb4__30_v_i80;

assign local_bb4__30_v_i80 = (local_bb4_cmp96_i70 ? local_bb4_cmp76_i64 : local_bb4_cmp88_i75);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool109_i78_stall_local;
wire [7:0] local_bb4_frombool109_i78;

assign local_bb4_frombool109_i78[7:1] = 7'h0;
assign local_bb4_frombool109_i78[0] = local_bb4_cmp85_i76;

// This section implements an unregistered operation.
// 
wire local_bb4_or107_i77_stall_local;
wire [31:0] local_bb4_or107_i77;

assign local_bb4_or107_i77[31:1] = 31'h0;
assign local_bb4_or107_i77[0] = local_bb4_var__u101;

// This section implements an unregistered operation.
// 
wire local_bb4_add245_i_stall_local;
wire [31:0] local_bb4_add245_i;

assign local_bb4_add245_i = (local_bb4_cond244_i + (rnode_392to394_bb4_and17_i_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i10_stall_local;
wire [31:0] local_bb4_fold_i10;

assign local_bb4_fold_i10 = (local_bb4_cond244_i + (rnode_392to394_bb4_shr16_i_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl207_i_stall_local;
wire [31:0] local_bb4_shl207_i;

assign local_bb4_shl207_i = ((local_bb4_and205_i & 32'h7FFFFFF) << (local_bb4_and206_i & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb4_or1596_i101_stall_local;
wire [31:0] local_bb4_or1596_i101;

assign local_bb4_or1596_i101 = (local_bb4_var__u102 | (local_bb4_and142_i95 & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i83_stall_local;
wire [7:0] local_bb4__31_i83;

assign local_bb4__31_i83[7:1] = 7'h0;
assign local_bb4__31_i83[0] = local_bb4__31_v_i82;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i81_stall_local;
wire [7:0] local_bb4__30_i81;

assign local_bb4__30_i81[7:1] = 7'h0;
assign local_bb4__30_i81[0] = local_bb4__30_v_i80;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i79_stall_local;
wire [7:0] local_bb4__29_i79;

assign local_bb4__29_i79 = (local_bb4_cmp96_i70 ? (local_bb4_frombool74_i62 & 8'h1) : (local_bb4_frombool109_i78 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i84_stall_local;
wire [31:0] local_bb4__32_i84;

assign local_bb4__32_i84 = (local_bb4_cmp96_i70 ? 32'h0 : (local_bb4_or107_i77 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i_stall_local;
wire [31:0] local_bb4_and250_i;

assign local_bb4_and250_i = (local_bb4_fold_i10 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and269_i_stall_local;
wire [31:0] local_bb4_and269_i;

assign local_bb4_and269_i = (local_bb4_fold_i10 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and208_i_stall_local;
wire [31:0] local_bb4_and208_i;

assign local_bb4_and208_i = (local_bb4_shl207_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_or162_i102_stall_local;
wire [31:0] local_bb4_or162_i102;

assign local_bb4_or162_i102 = (local_bb4_or1596_i101 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1237_i87_stall_local;
wire [7:0] local_bb4_or1237_i87;

assign local_bb4_or1237_i87 = ((local_bb4__30_i81 & 8'h1) | (local_bb4__29_i79 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i89_stall_local;
wire [7:0] local_bb4__33_i89;

assign local_bb4__33_i89 = (local_bb4_cmp116_i86 ? (local_bb4__29_i79 & 8'h1) : (local_bb4__31_i83 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__44_i_stall_local;
wire [31:0] local_bb4__44_i;

assign local_bb4__44_i = (local_bb4__40_demorgan_i ? (local_bb4_and208_i & 32'h7FFFFFF) : (local_bb4_or219_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i103_stall_local;
wire [31:0] local_bb4__37_v_i103;

assign local_bb4__37_v_i103 = (local_bb4_Pivot20_i98 ? 32'h0 : (local_bb4_or162_i102 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or123_i88_stall_local;
wire [31:0] local_bb4_or123_i88;

assign local_bb4_or123_i88[31:8] = 24'h0;
assign local_bb4_or123_i88[7:0] = (local_bb4_or1237_i87 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u103_stall_local;
wire [7:0] local_bb4_var__u103;

assign local_bb4_var__u103 = ((local_bb4__33_i89 & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i_valid_out;
wire local_bb4_and250_i_stall_in;
wire local_bb4_and269_i_valid_out;
wire local_bb4_and269_i_stall_in;
wire local_bb4_add245_i_valid_out;
wire local_bb4_add245_i_stall_in;
wire local_bb4__45_i_valid_out;
wire local_bb4__45_i_stall_in;
wire local_bb4_not_cmp37_i_valid_out_1;
wire local_bb4_not_cmp37_i_stall_in_1;
wire local_bb4__45_i_inputs_ready;
wire local_bb4__45_i_stall_local;
wire [31:0] local_bb4__45_i;

assign local_bb4__45_i_inputs_ready = (rnode_392to394_bb4_shr16_i_0_valid_out_NO_SHIFT_REG & rnode_392to394_bb4_and17_i_0_valid_out_NO_SHIFT_REG & rnode_392to394_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG & rnode_392to394_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG & rnode_393to394_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG & rnode_392to394_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG & rnode_393to394_bb4_and195_i_0_valid_out_NO_SHIFT_REG & rnode_393to394_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG & rnode_393to394_bb4_and198_i_0_valid_out_NO_SHIFT_REG & rnode_393to394_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG & rnode_393to394_bb4__and_i_i9_0_valid_out_1_NO_SHIFT_REG & rnode_393to394_bb4__and_i_i9_0_valid_out_2_NO_SHIFT_REG & rnode_393to394_bb4__and_i_i9_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i = (local_bb4__42_i ? (rnode_393to394_bb4_and193_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i & 32'h7FFFFFF));
assign local_bb4_and250_i_valid_out = 1'b1;
assign local_bb4_and269_i_valid_out = 1'b1;
assign local_bb4_add245_i_valid_out = 1'b1;
assign local_bb4__45_i_valid_out = 1'b1;
assign local_bb4_not_cmp37_i_valid_out_1 = 1'b1;
assign rnode_392to394_bb4_shr16_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_and17_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_cmp37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_392to394_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and195_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and198_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4_and193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4__and_i_i9_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4__and_i_i9_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_393to394_bb4__and_i_i9_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i104_stall_local;
wire [31:0] local_bb4__39_v_i104;

assign local_bb4__39_v_i104 = (local_bb4_SwitchLeaf_i99 ? (local_bb4_var__u100 & 32'h1) : (local_bb4__37_v_i103 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i90_stall_local;
wire [31:0] local_bb4_or124_i90;

assign local_bb4_or124_i90 = (local_bb4_cmp116_i86 ? 32'h0 : (local_bb4_or123_i88 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv135_i92_stall_local;
wire [31:0] local_bb4_conv135_i92;

assign local_bb4_conv135_i92[31:8] = 24'h0;
assign local_bb4_conv135_i92[7:0] = (local_bb4_var__u103 & 8'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_and250_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and250_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_and250_i_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and250_i_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_and250_i_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and250_i_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and250_i_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_and250_i_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_and250_i_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_and250_i_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_and250_i_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_and250_i_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_and250_i_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in((local_bb4_and250_i & 32'hFF)),
	.data_out(rnode_394to395_bb4_and250_i_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_and250_i_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_and250_i_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_394to395_bb4_and250_i_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_and250_i_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_and250_i_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and250_i_stall_in = 1'b0;
assign rnode_394to395_bb4_and250_i_0_NO_SHIFT_REG = rnode_394to395_bb4_and250_i_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_and250_i_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_and250_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_394to396_bb4_and269_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_394to396_bb4_and269_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_394to396_bb4_and269_i_0_NO_SHIFT_REG;
 logic rnode_394to396_bb4_and269_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to396_bb4_and269_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_394to396_bb4_and269_i_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_394to396_bb4_and269_i_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_394to396_bb4_and269_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_394to396_bb4_and269_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to396_bb4_and269_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to396_bb4_and269_i_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_394to396_bb4_and269_i_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_394to396_bb4_and269_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in((local_bb4_and269_i & 32'hFF800000)),
	.data_out(rnode_394to396_bb4_and269_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_394to396_bb4_and269_i_0_reg_396_fifo.DEPTH = 2;
defparam rnode_394to396_bb4_and269_i_0_reg_396_fifo.DATA_WIDTH = 32;
defparam rnode_394to396_bb4_and269_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to396_bb4_and269_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_394to396_bb4_and269_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and269_i_stall_in = 1'b0;
assign rnode_394to396_bb4_and269_i_0_NO_SHIFT_REG = rnode_394to396_bb4_and269_i_0_reg_396_NO_SHIFT_REG;
assign rnode_394to396_bb4_and269_i_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_394to396_bb4_and269_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_add245_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_add245_i_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4_add245_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_add245_i_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4_add245_i_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4_add245_i_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_add245_i_0_valid_out_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_add245_i_0_stall_in_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_add245_i_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_add245_i_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_add245_i_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_add245_i_0_stall_in_0_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_add245_i_0_valid_out_0_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_add245_i_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(local_bb4_add245_i),
	.data_out(rnode_394to395_bb4_add245_i_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_add245_i_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_add245_i_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_394to395_bb4_add245_i_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_add245_i_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_add245_i_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add245_i_stall_in = 1'b0;
assign rnode_394to395_bb4_add245_i_0_stall_in_0_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4_add245_i_0_NO_SHIFT_REG = rnode_394to395_bb4_add245_i_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4_add245_i_1_NO_SHIFT_REG = rnode_394to395_bb4_add245_i_0_reg_395_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4__45_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4__45_i_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4__45_i_1_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4__45_i_2_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_394to395_bb4__45_i_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_valid_out_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_stall_in_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4__45_i_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4__45_i_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4__45_i_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4__45_i_0_stall_in_0_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4__45_i_0_valid_out_0_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4__45_i_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in((local_bb4__45_i & 32'hFFFFFFF)),
	.data_out(rnode_394to395_bb4__45_i_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4__45_i_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4__45_i_0_reg_395_fifo.DATA_WIDTH = 32;
defparam rnode_394to395_bb4__45_i_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4__45_i_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4__45_i_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i_stall_in = 1'b0;
assign rnode_394to395_bb4__45_i_0_stall_in_0_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4__45_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4__45_i_0_NO_SHIFT_REG = rnode_394to395_bb4__45_i_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4__45_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4__45_i_1_NO_SHIFT_REG = rnode_394to395_bb4__45_i_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4__45_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_394to395_bb4__45_i_2_NO_SHIFT_REG = rnode_394to395_bb4__45_i_0_reg_395_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_394to395_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_394to395_bb4_not_cmp37_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_394to395_bb4_not_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_394to395_bb4_not_cmp37_i_0_reg_395_inputs_ready_NO_SHIFT_REG;
 logic rnode_394to395_bb4_not_cmp37_i_0_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_not_cmp37_i_0_valid_out_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_not_cmp37_i_0_stall_in_reg_395_NO_SHIFT_REG;
 logic rnode_394to395_bb4_not_cmp37_i_0_stall_out_reg_395_NO_SHIFT_REG;

acl_data_fifo rnode_394to395_bb4_not_cmp37_i_0_reg_395_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_394to395_bb4_not_cmp37_i_0_reg_395_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_394to395_bb4_not_cmp37_i_0_stall_in_reg_395_NO_SHIFT_REG),
	.valid_out(rnode_394to395_bb4_not_cmp37_i_0_valid_out_reg_395_NO_SHIFT_REG),
	.stall_out(rnode_394to395_bb4_not_cmp37_i_0_stall_out_reg_395_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp37_i),
	.data_out(rnode_394to395_bb4_not_cmp37_i_0_reg_395_NO_SHIFT_REG)
);

defparam rnode_394to395_bb4_not_cmp37_i_0_reg_395_fifo.DEPTH = 1;
defparam rnode_394to395_bb4_not_cmp37_i_0_reg_395_fifo.DATA_WIDTH = 1;
defparam rnode_394to395_bb4_not_cmp37_i_0_reg_395_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_394to395_bb4_not_cmp37_i_0_reg_395_fifo.IMPL = "shift_reg";

assign rnode_394to395_bb4_not_cmp37_i_0_reg_395_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp37_i_stall_in_1 = 1'b0;
assign rnode_394to395_bb4_not_cmp37_i_0_NO_SHIFT_REG = rnode_394to395_bb4_not_cmp37_i_0_reg_395_NO_SHIFT_REG;
assign rnode_394to395_bb4_not_cmp37_i_0_stall_in_reg_395_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i105_stall_local;
wire [31:0] local_bb4_reduction_3_i105;

assign local_bb4_reduction_3_i105 = ((local_bb4__32_i84 & 32'h1) | (local_bb4_or124_i90 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or136_i94_stall_local;
wire [31:0] local_bb4_or136_i94;

assign local_bb4_or136_i94 = (local_bb4_cmp131_not_i93 ? (local_bb4_conv135_i92 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i_stall_local;
wire local_bb4_notrhs_i;

assign local_bb4_notrhs_i = ((rnode_394to395_bb4_and250_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl273_i_stall_local;
wire [31:0] local_bb4_shl273_i;

assign local_bb4_shl273_i = ((rnode_394to396_bb4_and269_i_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and247_i_stall_local;
wire [31:0] local_bb4_and247_i;

assign local_bb4_and247_i = (rnode_394to395_bb4_add245_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp258_i_stall_local;
wire local_bb4_cmp258_i;

assign local_bb4_cmp258_i = ($signed(rnode_394to395_bb4_add245_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and225_i_stall_local;
wire [31:0] local_bb4_and225_i;

assign local_bb4_and225_i = ((rnode_394to395_bb4__45_i_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i_stall_local;
wire [31:0] local_bb4_and270_i;

assign local_bb4_and270_i = ((rnode_394to395_bb4__45_i_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr271_i_valid_out;
wire local_bb4_shr271_i_stall_in;
wire local_bb4_shr271_i_inputs_ready;
wire local_bb4_shr271_i_stall_local;
wire [31:0] local_bb4_shr271_i;

assign local_bb4_shr271_i_inputs_ready = rnode_394to395_bb4__45_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr271_i = ((rnode_394to395_bb4__45_i_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr271_i_valid_out = 1'b1;
assign rnode_394to395_bb4__45_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i107_stall_local;
wire [31:0] local_bb4_reduction_5_i107;

assign local_bb4_reduction_5_i107 = (local_bb4_shr150_i97 | (local_bb4_reduction_3_i105 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i106_stall_local;
wire [31:0] local_bb4_reduction_4_i106;

assign local_bb4_reduction_4_i106 = ((local_bb4_or136_i94 & 32'h1) | (local_bb4__39_v_i104 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i_stall_local;
wire local_bb4_notlhs_i;

assign local_bb4_notlhs_i = ((local_bb4_and247_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_i_stall_local;
wire local_bb4_cmp226_i;

assign local_bb4_cmp226_i = ((local_bb4_and225_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i_stall_local;
wire local_bb4_cmp296_i;

assign local_bb4_cmp296_i = ((local_bb4_and270_i & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i_valid_out;
wire local_bb4_cmp296_i_stall_in;
wire local_bb4_cmp299_i_valid_out;
wire local_bb4_cmp299_i_stall_in;
wire local_bb4_cmp299_i_inputs_ready;
wire local_bb4_cmp299_i_stall_local;
wire local_bb4_cmp299_i;

assign local_bb4_cmp299_i_inputs_ready = rnode_394to395_bb4__45_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp299_i = ((local_bb4_and270_i & 32'h7) == 32'h4);
assign local_bb4_cmp296_i_valid_out = 1'b1;
assign local_bb4_cmp299_i_valid_out = 1'b1;
assign rnode_394to395_bb4__45_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_shr271_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_395to396_bb4_shr271_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_shr271_i_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_shr271_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_shr271_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_shr271_i_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_shr271_i_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_shr271_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_shr271_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_shr271_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_shr271_i_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_shr271_i_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_shr271_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in((local_bb4_shr271_i & 32'h1FFFFFF)),
	.data_out(rnode_395to396_bb4_shr271_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_shr271_i_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_shr271_i_0_reg_396_fifo.DATA_WIDTH = 32;
defparam rnode_395to396_bb4_shr271_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_shr271_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_shr271_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr271_i_stall_in = 1'b0;
assign rnode_395to396_bb4_shr271_i_0_NO_SHIFT_REG = rnode_395to396_bb4_shr271_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_shr271_i_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_shr271_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i108_stall_local;
wire [31:0] local_bb4_reduction_6_i108;

assign local_bb4_reduction_6_i108 = ((local_bb4_reduction_4_i106 & 32'h1) | local_bb4_reduction_5_i107);

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i_stall_local;
wire local_bb4_not__46_i;

assign local_bb4_not__46_i = (local_bb4_notrhs_i | local_bb4_notlhs_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_not_i_stall_local;
wire local_bb4_cmp226_not_i;

assign local_bb4_cmp226_not_i = (local_bb4_cmp226_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp296_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp296_i_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp296_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp296_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp296_i_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp296_i_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp296_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_cmp296_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_cmp296_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_cmp296_i_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_cmp296_i_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_cmp296_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(local_bb4_cmp296_i),
	.data_out(rnode_395to396_bb4_cmp296_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_cmp296_i_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_cmp296_i_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_395to396_bb4_cmp296_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_cmp296_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_cmp296_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp296_i_stall_in = 1'b0;
assign rnode_395to396_bb4_cmp296_i_0_NO_SHIFT_REG = rnode_395to396_bb4_cmp296_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_cmp296_i_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp299_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp299_i_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp299_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp299_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp299_i_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp299_i_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_cmp299_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_cmp299_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_cmp299_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_cmp299_i_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_cmp299_i_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_cmp299_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(local_bb4_cmp299_i),
	.data_out(rnode_395to396_bb4_cmp299_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_cmp299_i_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_cmp299_i_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_395to396_bb4_cmp299_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_cmp299_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_cmp299_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp299_i_stall_in = 1'b0;
assign rnode_395to396_bb4_cmp299_i_0_NO_SHIFT_REG = rnode_395to396_bb4_cmp299_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_cmp299_i_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and272_i_stall_local;
wire [31:0] local_bb4_and272_i;

assign local_bb4_and272_i = ((rnode_395to396_bb4_shr271_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i40_valid_out;
wire local_bb4_lnot33_not_i40_stall_in;
wire local_bb4_cmp37_i36_valid_out;
wire local_bb4_cmp37_i36_stall_in;
wire local_bb4_and36_lobit_i111_valid_out;
wire local_bb4_and36_lobit_i111_stall_in;
wire local_bb4_xor188_i110_valid_out;
wire local_bb4_xor188_i110_stall_in;
wire local_bb4_xor188_i110_inputs_ready;
wire local_bb4_xor188_i110_stall_local;
wire [31:0] local_bb4_xor188_i110;

assign local_bb4_xor188_i110_inputs_ready = (rnode_395to396_bb4__22_i22_0_valid_out_0_NO_SHIFT_REG & rnode_395to396_bb4_lnot23_i31_0_valid_out_NO_SHIFT_REG & rnode_395to396_bb4_align_0_i59_0_valid_out_0_NO_SHIFT_REG & rnode_395to396_bb4_align_0_i59_0_valid_out_4_NO_SHIFT_REG & rnode_395to396_bb4_align_0_i59_0_valid_out_1_NO_SHIFT_REG & rnode_395to396_bb4_align_0_i59_0_valid_out_2_NO_SHIFT_REG & rnode_395to396_bb4_align_0_i59_0_valid_out_3_NO_SHIFT_REG & rnode_395to396_bb4__23_i23_0_valid_out_2_NO_SHIFT_REG & rnode_395to396_bb4__22_i22_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor188_i110 = (local_bb4_reduction_6_i108 ^ local_bb4_xor_lobit_i109);
assign local_bb4_lnot33_not_i40_valid_out = 1'b1;
assign local_bb4_cmp37_i36_valid_out = 1'b1;
assign local_bb4_and36_lobit_i111_valid_out = 1'b1;
assign local_bb4_xor188_i110_valid_out = 1'b1;
assign rnode_395to396_bb4__22_i22_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_lnot23_i31_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_align_0_i59_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_align_0_i59_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_align_0_i59_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_align_0_i59_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_align_0_i59_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__23_i23_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__22_i22_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__47_i_stall_local;
wire local_bb4__47_i;

assign local_bb4__47_i = (local_bb4_cmp226_i | local_bb4_not__46_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i_stall_local;
wire local_bb4_brmerge12_i;

assign local_bb4_brmerge12_i = (local_bb4_cmp226_not_i | rnode_394to395_bb4_not_cmp37_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot262__i_stall_local;
wire local_bb4_lnot262__i;

assign local_bb4_lnot262__i = (local_bb4_cmp258_i & local_bb4_cmp226_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29649_i_stall_local;
wire [31:0] local_bb4_cmp29649_i;

assign local_bb4_cmp29649_i[31:1] = 31'h0;
assign local_bb4_cmp29649_i[0] = rnode_395to396_bb4_cmp296_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv300_i_stall_local;
wire [31:0] local_bb4_conv300_i;

assign local_bb4_conv300_i[31:1] = 31'h0;
assign local_bb4_conv300_i[0] = rnode_395to396_bb4_cmp299_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or274_i_stall_local;
wire [31:0] local_bb4_or274_i;

assign local_bb4_or274_i = ((local_bb4_and272_i & 32'h7FFFFF) | (local_bb4_shl273_i & 32'h7F800000));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_lnot33_not_i40_0_valid_out_NO_SHIFT_REG;
 logic rnode_396to397_bb4_lnot33_not_i40_0_stall_in_NO_SHIFT_REG;
 logic rnode_396to397_bb4_lnot33_not_i40_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_lnot33_not_i40_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic rnode_396to397_bb4_lnot33_not_i40_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_lnot33_not_i40_0_valid_out_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_lnot33_not_i40_0_stall_in_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_lnot33_not_i40_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_lnot33_not_i40_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_lnot33_not_i40_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_lnot33_not_i40_0_stall_in_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_lnot33_not_i40_0_valid_out_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_lnot33_not_i40_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i40),
	.data_out(rnode_396to397_bb4_lnot33_not_i40_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_lnot33_not_i40_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_lnot33_not_i40_0_reg_397_fifo.DATA_WIDTH = 1;
defparam rnode_396to397_bb4_lnot33_not_i40_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_lnot33_not_i40_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_lnot33_not_i40_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i40_stall_in = 1'b0;
assign rnode_396to397_bb4_lnot33_not_i40_0_NO_SHIFT_REG = rnode_396to397_bb4_lnot33_not_i40_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_lnot33_not_i40_0_stall_in_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_lnot33_not_i40_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_valid_out_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_stall_in_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_cmp37_i36_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_cmp37_i36_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_cmp37_i36_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_cmp37_i36_0_stall_in_0_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_cmp37_i36_0_valid_out_0_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_cmp37_i36_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(local_bb4_cmp37_i36),
	.data_out(rnode_396to397_bb4_cmp37_i36_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_cmp37_i36_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_cmp37_i36_0_reg_397_fifo.DATA_WIDTH = 1;
defparam rnode_396to397_bb4_cmp37_i36_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_cmp37_i36_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_cmp37_i36_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp37_i36_stall_in = 1'b0;
assign rnode_396to397_bb4_cmp37_i36_0_stall_in_0_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_cmp37_i36_0_NO_SHIFT_REG = rnode_396to397_bb4_cmp37_i36_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_cmp37_i36_1_NO_SHIFT_REG = rnode_396to397_bb4_cmp37_i36_0_reg_397_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_and36_lobit_i111_0_valid_out_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and36_lobit_i111_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_and36_lobit_i111_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and36_lobit_i111_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_and36_lobit_i111_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and36_lobit_i111_0_valid_out_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and36_lobit_i111_0_stall_in_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_and36_lobit_i111_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_and36_lobit_i111_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_and36_lobit_i111_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_and36_lobit_i111_0_stall_in_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_and36_lobit_i111_0_valid_out_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_and36_lobit_i111_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in((local_bb4_and36_lobit_i111 & 32'h1)),
	.data_out(rnode_396to397_bb4_and36_lobit_i111_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_and36_lobit_i111_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_and36_lobit_i111_0_reg_397_fifo.DATA_WIDTH = 32;
defparam rnode_396to397_bb4_and36_lobit_i111_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_and36_lobit_i111_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_and36_lobit_i111_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and36_lobit_i111_stall_in = 1'b0;
assign rnode_396to397_bb4_and36_lobit_i111_0_NO_SHIFT_REG = rnode_396to397_bb4_and36_lobit_i111_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_and36_lobit_i111_0_stall_in_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_and36_lobit_i111_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4_xor188_i110_0_valid_out_NO_SHIFT_REG;
 logic rnode_396to397_bb4_xor188_i110_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_xor188_i110_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4_xor188_i110_0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4_xor188_i110_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_xor188_i110_0_valid_out_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_xor188_i110_0_stall_in_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4_xor188_i110_0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4_xor188_i110_0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4_xor188_i110_0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4_xor188_i110_0_stall_in_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4_xor188_i110_0_valid_out_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4_xor188_i110_0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(local_bb4_xor188_i110),
	.data_out(rnode_396to397_bb4_xor188_i110_0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4_xor188_i110_0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4_xor188_i110_0_reg_397_fifo.DATA_WIDTH = 32;
defparam rnode_396to397_bb4_xor188_i110_0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4_xor188_i110_0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4_xor188_i110_0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor188_i110_stall_in = 1'b0;
assign rnode_396to397_bb4_xor188_i110_0_NO_SHIFT_REG = rnode_396to397_bb4_xor188_i110_0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4_xor188_i110_0_stall_in_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_xor188_i110_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i_stall_local;
wire [31:0] local_bb4_resultSign_0_i;

assign local_bb4_resultSign_0_i = (local_bb4_brmerge12_i ? (rnode_394to395_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i_valid_out;
wire local_bb4_resultSign_0_i_stall_in;
wire local_bb4__47_i_valid_out;
wire local_bb4__47_i_stall_in;
wire local_bb4_or2662_i_valid_out;
wire local_bb4_or2662_i_stall_in;
wire local_bb4_or2662_i_inputs_ready;
wire local_bb4_or2662_i_stall_local;
wire local_bb4_or2662_i;

assign local_bb4_or2662_i_inputs_ready = (rnode_394to395_bb4_and35_i_0_valid_out_NO_SHIFT_REG & rnode_394to395_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG & rnode_394to395_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG & rnode_394to395_bb4_and250_i_0_valid_out_NO_SHIFT_REG & rnode_394to395_bb4__45_i_0_valid_out_0_NO_SHIFT_REG & rnode_394to395_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG & rnode_394to395_bb4_var__u88_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2662_i = (rnode_394to395_bb4_var__u88_0_NO_SHIFT_REG | local_bb4_lnot262__i);
assign local_bb4_resultSign_0_i_valid_out = 1'b1;
assign local_bb4__47_i_valid_out = 1'b1;
assign local_bb4_or2662_i_valid_out = 1'b1;
assign rnode_394to395_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_not_cmp37_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_add245_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_and250_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4__45_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_add245_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_394to395_bb4_var__u88_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i41_stall_local;
wire local_bb4_brmerge_not_i41;

assign local_bb4_brmerge_not_i41 = (rnode_395to397_bb4_cmp27_i33_0_NO_SHIFT_REG & rnode_396to397_bb4_lnot33_not_i40_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_397to399_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_1_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_2_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_valid_out_0_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_stall_in_0_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_cmp37_i36_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_397to399_bb4_cmp37_i36_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to399_bb4_cmp37_i36_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to399_bb4_cmp37_i36_0_stall_in_0_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_397to399_bb4_cmp37_i36_0_valid_out_0_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_397to399_bb4_cmp37_i36_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in(rnode_396to397_bb4_cmp37_i36_1_NO_SHIFT_REG),
	.data_out(rnode_397to399_bb4_cmp37_i36_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_397to399_bb4_cmp37_i36_0_reg_399_fifo.DEPTH = 2;
defparam rnode_397to399_bb4_cmp37_i36_0_reg_399_fifo.DATA_WIDTH = 1;
defparam rnode_397to399_bb4_cmp37_i36_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to399_bb4_cmp37_i36_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_397to399_bb4_cmp37_i36_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_cmp37_i36_0_stall_in_0_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_397to399_bb4_cmp37_i36_0_NO_SHIFT_REG = rnode_397to399_bb4_cmp37_i36_0_reg_399_NO_SHIFT_REG;
assign rnode_397to399_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_397to399_bb4_cmp37_i36_1_NO_SHIFT_REG = rnode_397to399_bb4_cmp37_i36_0_reg_399_NO_SHIFT_REG;
assign rnode_397to399_bb4_cmp37_i36_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_397to399_bb4_cmp37_i36_2_NO_SHIFT_REG = rnode_397to399_bb4_cmp37_i36_0_reg_399_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i112_stall_local;
wire [31:0] local_bb4_add_i112;

assign local_bb4_add_i112 = ((local_bb4__27_i52 & 32'h7FFFFF8) | (rnode_396to397_bb4_and36_lobit_i111_0_NO_SHIFT_REG & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_395to396_bb4_resultSign_0_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_resultSign_0_i_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_resultSign_0_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_395to396_bb4_resultSign_0_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_resultSign_0_i_0_valid_out_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_resultSign_0_i_0_stall_in_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_resultSign_0_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_resultSign_0_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_resultSign_0_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_resultSign_0_i_0_stall_in_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_resultSign_0_i_0_valid_out_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_resultSign_0_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i & 32'h80000000)),
	.data_out(rnode_395to396_bb4_resultSign_0_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_resultSign_0_i_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_resultSign_0_i_0_reg_396_fifo.DATA_WIDTH = 32;
defparam rnode_395to396_bb4_resultSign_0_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_resultSign_0_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_resultSign_0_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i_stall_in = 1'b0;
assign rnode_395to396_bb4_resultSign_0_i_0_NO_SHIFT_REG = rnode_395to396_bb4_resultSign_0_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_resultSign_0_i_0_stall_in_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4__47_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_valid_out_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_stall_in_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4__47_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4__47_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4__47_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4__47_i_0_stall_in_0_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4__47_i_0_valid_out_0_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4__47_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(local_bb4__47_i),
	.data_out(rnode_395to396_bb4__47_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4__47_i_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4__47_i_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_395to396_bb4__47_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4__47_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4__47_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i_stall_in = 1'b0;
assign rnode_395to396_bb4__47_i_0_stall_in_0_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__47_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__47_i_0_NO_SHIFT_REG = rnode_395to396_bb4__47_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4__47_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4__47_i_1_NO_SHIFT_REG = rnode_395to396_bb4__47_i_0_reg_396_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_395to396_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_1_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_2_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_reg_396_inputs_ready_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_valid_out_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_stall_in_0_reg_396_NO_SHIFT_REG;
 logic rnode_395to396_bb4_or2662_i_0_stall_out_reg_396_NO_SHIFT_REG;

acl_data_fifo rnode_395to396_bb4_or2662_i_0_reg_396_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_395to396_bb4_or2662_i_0_reg_396_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_395to396_bb4_or2662_i_0_stall_in_0_reg_396_NO_SHIFT_REG),
	.valid_out(rnode_395to396_bb4_or2662_i_0_valid_out_0_reg_396_NO_SHIFT_REG),
	.stall_out(rnode_395to396_bb4_or2662_i_0_stall_out_reg_396_NO_SHIFT_REG),
	.data_in(local_bb4_or2662_i),
	.data_out(rnode_395to396_bb4_or2662_i_0_reg_396_NO_SHIFT_REG)
);

defparam rnode_395to396_bb4_or2662_i_0_reg_396_fifo.DEPTH = 1;
defparam rnode_395to396_bb4_or2662_i_0_reg_396_fifo.DATA_WIDTH = 1;
defparam rnode_395to396_bb4_or2662_i_0_reg_396_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_395to396_bb4_or2662_i_0_reg_396_fifo.IMPL = "shift_reg";

assign rnode_395to396_bb4_or2662_i_0_reg_396_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2662_i_stall_in = 1'b0;
assign rnode_395to396_bb4_or2662_i_0_stall_in_0_reg_396_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_or2662_i_0_NO_SHIFT_REG = rnode_395to396_bb4_or2662_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_or2662_i_1_NO_SHIFT_REG = rnode_395to396_bb4_or2662_i_0_reg_396_NO_SHIFT_REG;
assign rnode_395to396_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_395to396_bb4_or2662_i_2_NO_SHIFT_REG = rnode_395to396_bb4_or2662_i_0_reg_396_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__24_i44_stall_local;
wire local_bb4__24_i44;

assign local_bb4__24_i44 = (local_bb4_or_cond_not_i43 | local_bb4_brmerge_not_i41);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i45_stall_local;
wire local_bb4_brmerge_not_not_i45;

assign local_bb4_brmerge_not_not_i45 = (local_bb4_brmerge_not_i41 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp37_i142_stall_local;
wire local_bb4_not_cmp37_i142;

assign local_bb4_not_cmp37_i142 = (rnode_397to399_bb4_cmp37_i36_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add192_i113_stall_local;
wire [31:0] local_bb4_add192_i113;

assign local_bb4_add192_i113 = ((local_bb4_add_i112 & 32'h7FFFFF9) + rnode_396to397_bb4_xor188_i110_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i_stall_local;
wire [31:0] local_bb4_or275_i;

assign local_bb4_or275_i = ((local_bb4_or274_i & 32'h7FFFFFFF) | (rnode_395to396_bb4_resultSign_0_i_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u104_stall_local;
wire [31:0] local_bb4_var__u104;

assign local_bb4_var__u104[31:1] = 31'h0;
assign local_bb4_var__u104[0] = rnode_395to396_bb4__47_i_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2804_i_stall_local;
wire local_bb4_or2804_i;

assign local_bb4_or2804_i = (rnode_395to396_bb4__47_i_0_NO_SHIFT_REG | rnode_395to396_bb4_or2662_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2875_i_stall_local;
wire local_bb4_or2875_i;

assign local_bb4_or2875_i = (rnode_395to396_bb4_or2662_i_1_NO_SHIFT_REG | rnode_395to396_bb4__26_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u105_stall_local;
wire [31:0] local_bb4_var__u105;

assign local_bb4_var__u105[31:1] = 31'h0;
assign local_bb4_var__u105[0] = rnode_395to396_bb4_or2662_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i46_stall_local;
wire local_bb4_reduction_7_i46;

assign local_bb4_reduction_7_i46 = (local_bb4_cmp25_i32 & local_bb4_brmerge_not_not_i45);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext314_i_stall_local;
wire [31:0] local_bb4_lnot_ext314_i;

assign local_bb4_lnot_ext314_i = ((local_bb4_var__u104 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond282_i_stall_local;
wire [31:0] local_bb4_cond282_i;

assign local_bb4_cond282_i = (local_bb4_or2804_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond289_i_stall_local;
wire [31:0] local_bb4_cond289_i;

assign local_bb4_cond289_i = (local_bb4_or2875_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext310_i_stall_local;
wire [31:0] local_bb4_lnot_ext310_i;

assign local_bb4_lnot_ext310_i = ((local_bb4_var__u105 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i48_stall_local;
wire local_bb4_reduction_9_i48;

assign local_bb4_reduction_9_i48 = (local_bb4_reduction_7_i46 & local_bb4_reduction_8_i47);

// This section implements an unregistered operation.
// 
wire local_bb4_and293_i_stall_local;
wire [31:0] local_bb4_and293_i;

assign local_bb4_and293_i = ((local_bb4_cond282_i | 32'h80000000) & local_bb4_or275_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or294_i_stall_local;
wire [31:0] local_bb4_or294_i;

assign local_bb4_or294_i = ((local_bb4_cond289_i & 32'h7F800000) | (local_bb4_cond292_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i_stall_local;
wire [31:0] local_bb4_reduction_0_i;

assign local_bb4_reduction_0_i = ((local_bb4_lnot_ext310_i & 32'h1) & (local_bb4_lnot_ext_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i25_valid_out_2;
wire local_bb4_and17_i25_stall_in_2;
wire local_bb4_var__u98_valid_out;
wire local_bb4_var__u98_stall_in;
wire local_bb4_add192_i113_valid_out;
wire local_bb4_add192_i113_stall_in;
wire local_bb4__26_i49_valid_out;
wire local_bb4__26_i49_stall_in;
wire local_bb4__26_i49_inputs_ready;
wire local_bb4__26_i49_stall_local;
wire local_bb4__26_i49;

assign local_bb4__26_i49_inputs_ready = (rnode_395to397_bb4_shr16_i24_0_valid_out_0_NO_SHIFT_REG & rnode_395to397_bb4_cmp27_i33_0_valid_out_2_NO_SHIFT_REG & rnode_396to397_bb4_and36_lobit_i111_0_valid_out_NO_SHIFT_REG & rnode_396to397_bb4_xor188_i110_0_valid_out_NO_SHIFT_REG & rnode_396to397_bb4_and20_i28_0_valid_out_0_NO_SHIFT_REG & rnode_395to397_bb4_cmp27_i33_0_valid_out_0_NO_SHIFT_REG & rnode_396to397_bb4_lnot33_not_i40_0_valid_out_NO_SHIFT_REG & rnode_395to397_bb4_cmp27_i33_0_valid_out_1_NO_SHIFT_REG & rnode_396to397_bb4_and20_i28_0_valid_out_1_NO_SHIFT_REG & rnode_396to397_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i49 = (local_bb4_reduction_9_i48 ? rnode_396to397_bb4_cmp37_i36_0_NO_SHIFT_REG : local_bb4__24_i44);
assign local_bb4_and17_i25_valid_out_2 = 1'b1;
assign local_bb4_var__u98_valid_out = 1'b1;
assign local_bb4_add192_i113_valid_out = 1'b1;
assign local_bb4__26_i49_valid_out = 1'b1;
assign rnode_395to397_bb4_shr16_i24_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to397_bb4_cmp27_i33_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_and36_lobit_i111_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_xor188_i110_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_and20_i28_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to397_bb4_cmp27_i33_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_lnot33_not_i40_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to397_bb4_cmp27_i33_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_and20_i28_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and302_i_stall_local;
wire [31:0] local_bb4_and302_i;

assign local_bb4_and302_i = ((local_bb4_conv300_i & 32'h1) & local_bb4_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i_stall_local;
wire [31:0] local_bb4_or295_i;

assign local_bb4_or295_i = ((local_bb4_or294_i & 32'h7FC00000) | local_bb4_and293_i);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_397to399_bb4_and17_i25_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and17_i25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_397to399_bb4_and17_i25_0_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and17_i25_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_397to399_bb4_and17_i25_0_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and17_i25_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and17_i25_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_397to399_bb4_and17_i25_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_397to399_bb4_and17_i25_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to399_bb4_and17_i25_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to399_bb4_and17_i25_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_397to399_bb4_and17_i25_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_397to399_bb4_and17_i25_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i25 & 32'hFF)),
	.data_out(rnode_397to399_bb4_and17_i25_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_397to399_bb4_and17_i25_0_reg_399_fifo.DEPTH = 2;
defparam rnode_397to399_bb4_and17_i25_0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_397to399_bb4_and17_i25_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to399_bb4_and17_i25_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_397to399_bb4_and17_i25_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i25_stall_in_2 = 1'b0;
assign rnode_397to399_bb4_and17_i25_0_NO_SHIFT_REG = rnode_397to399_bb4_and17_i25_0_reg_399_NO_SHIFT_REG;
assign rnode_397to399_bb4_and17_i25_0_stall_in_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_and17_i25_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_397to398_bb4_var__u98_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to398_bb4_var__u98_0_stall_in_NO_SHIFT_REG;
 logic rnode_397to398_bb4_var__u98_0_NO_SHIFT_REG;
 logic rnode_397to398_bb4_var__u98_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic rnode_397to398_bb4_var__u98_0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_var__u98_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_var__u98_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_var__u98_0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_397to398_bb4_var__u98_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to398_bb4_var__u98_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to398_bb4_var__u98_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_397to398_bb4_var__u98_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_397to398_bb4_var__u98_0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(local_bb4_var__u98),
	.data_out(rnode_397to398_bb4_var__u98_0_reg_398_NO_SHIFT_REG)
);

defparam rnode_397to398_bb4_var__u98_0_reg_398_fifo.DEPTH = 1;
defparam rnode_397to398_bb4_var__u98_0_reg_398_fifo.DATA_WIDTH = 1;
defparam rnode_397to398_bb4_var__u98_0_reg_398_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to398_bb4_var__u98_0_reg_398_fifo.IMPL = "shift_reg";

assign rnode_397to398_bb4_var__u98_0_reg_398_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u98_stall_in = 1'b0;
assign rnode_397to398_bb4_var__u98_0_NO_SHIFT_REG = rnode_397to398_bb4_var__u98_0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb4_var__u98_0_stall_in_reg_398_NO_SHIFT_REG = 1'b0;
assign rnode_397to398_bb4_var__u98_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_397to398_bb4_add192_i113_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb4_add192_i113_0_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb4_add192_i113_1_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb4_add192_i113_2_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb4_add192_i113_3_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb4_add192_i113_0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_valid_out_0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_stall_in_0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4_add192_i113_0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_397to398_bb4_add192_i113_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to398_bb4_add192_i113_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to398_bb4_add192_i113_0_stall_in_0_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_397to398_bb4_add192_i113_0_valid_out_0_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_397to398_bb4_add192_i113_0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(local_bb4_add192_i113),
	.data_out(rnode_397to398_bb4_add192_i113_0_reg_398_NO_SHIFT_REG)
);

defparam rnode_397to398_bb4_add192_i113_0_reg_398_fifo.DEPTH = 1;
defparam rnode_397to398_bb4_add192_i113_0_reg_398_fifo.DATA_WIDTH = 32;
defparam rnode_397to398_bb4_add192_i113_0_reg_398_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to398_bb4_add192_i113_0_reg_398_fifo.IMPL = "shift_reg";

assign rnode_397to398_bb4_add192_i113_0_reg_398_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add192_i113_stall_in = 1'b0;
assign rnode_397to398_bb4_add192_i113_0_stall_in_0_reg_398_NO_SHIFT_REG = 1'b0;
assign rnode_397to398_bb4_add192_i113_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4_add192_i113_0_NO_SHIFT_REG = rnode_397to398_bb4_add192_i113_0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb4_add192_i113_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4_add192_i113_1_NO_SHIFT_REG = rnode_397to398_bb4_add192_i113_0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb4_add192_i113_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4_add192_i113_2_NO_SHIFT_REG = rnode_397to398_bb4_add192_i113_0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb4_add192_i113_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4_add192_i113_3_NO_SHIFT_REG = rnode_397to398_bb4_add192_i113_0_reg_398_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_397to398_bb4__26_i49_0_valid_out_NO_SHIFT_REG;
 logic rnode_397to398_bb4__26_i49_0_stall_in_NO_SHIFT_REG;
 logic rnode_397to398_bb4__26_i49_0_NO_SHIFT_REG;
 logic rnode_397to398_bb4__26_i49_0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic rnode_397to398_bb4__26_i49_0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4__26_i49_0_valid_out_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4__26_i49_0_stall_in_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4__26_i49_0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_397to398_bb4__26_i49_0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to398_bb4__26_i49_0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to398_bb4__26_i49_0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_397to398_bb4__26_i49_0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_397to398_bb4__26_i49_0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(local_bb4__26_i49),
	.data_out(rnode_397to398_bb4__26_i49_0_reg_398_NO_SHIFT_REG)
);

defparam rnode_397to398_bb4__26_i49_0_reg_398_fifo.DEPTH = 1;
defparam rnode_397to398_bb4__26_i49_0_reg_398_fifo.DATA_WIDTH = 1;
defparam rnode_397to398_bb4__26_i49_0_reg_398_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to398_bb4__26_i49_0_reg_398_fifo.IMPL = "shift_reg";

assign rnode_397to398_bb4__26_i49_0_reg_398_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i49_stall_in = 1'b0;
assign rnode_397to398_bb4__26_i49_0_NO_SHIFT_REG = rnode_397to398_bb4__26_i49_0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb4__26_i49_0_stall_in_reg_398_NO_SHIFT_REG = 1'b0;
assign rnode_397to398_bb4__26_i49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i_stall_local;
wire [31:0] local_bb4_lor_ext_i;

assign local_bb4_lor_ext_i = ((local_bb4_cmp29649_i & 32'h1) | (local_bb4_and302_i & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_398to399_bb4_var__u98_0_valid_out_NO_SHIFT_REG;
 logic rnode_398to399_bb4_var__u98_0_stall_in_NO_SHIFT_REG;
 logic rnode_398to399_bb4_var__u98_0_NO_SHIFT_REG;
 logic rnode_398to399_bb4_var__u98_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic rnode_398to399_bb4_var__u98_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_var__u98_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_var__u98_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_var__u98_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_398to399_bb4_var__u98_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to399_bb4_var__u98_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to399_bb4_var__u98_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_398to399_bb4_var__u98_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_398to399_bb4_var__u98_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in(rnode_397to398_bb4_var__u98_0_NO_SHIFT_REG),
	.data_out(rnode_398to399_bb4_var__u98_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_398to399_bb4_var__u98_0_reg_399_fifo.DEPTH = 1;
defparam rnode_398to399_bb4_var__u98_0_reg_399_fifo.DATA_WIDTH = 1;
defparam rnode_398to399_bb4_var__u98_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to399_bb4_var__u98_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_398to399_bb4_var__u98_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4_var__u98_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_var__u98_0_NO_SHIFT_REG = rnode_398to399_bb4_var__u98_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4_var__u98_0_stall_in_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_var__u98_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and193_i114_valid_out;
wire local_bb4_and193_i114_stall_in;
wire local_bb4_and193_i114_inputs_ready;
wire local_bb4_and193_i114_stall_local;
wire [31:0] local_bb4_and193_i114;

assign local_bb4_and193_i114_inputs_ready = rnode_397to398_bb4_add192_i113_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and193_i114 = (rnode_397to398_bb4_add192_i113_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and193_i114_valid_out = 1'b1;
assign rnode_397to398_bb4_add192_i113_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and195_i115_valid_out;
wire local_bb4_and195_i115_stall_in;
wire local_bb4_and195_i115_inputs_ready;
wire local_bb4_and195_i115_stall_local;
wire [31:0] local_bb4_and195_i115;

assign local_bb4_and195_i115_inputs_ready = rnode_397to398_bb4_add192_i113_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and195_i115 = (rnode_397to398_bb4_add192_i113_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and195_i115_valid_out = 1'b1;
assign rnode_397to398_bb4_add192_i113_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and198_i116_valid_out;
wire local_bb4_and198_i116_stall_in;
wire local_bb4_and198_i116_inputs_ready;
wire local_bb4_and198_i116_stall_local;
wire [31:0] local_bb4_and198_i116;

assign local_bb4_and198_i116_inputs_ready = rnode_397to398_bb4_add192_i113_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and198_i116 = (rnode_397to398_bb4_add192_i113_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and198_i116_valid_out = 1'b1;
assign rnode_397to398_bb4_add192_i113_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and201_i117_stall_local;
wire [31:0] local_bb4_and201_i117;

assign local_bb4_and201_i117 = (rnode_397to398_bb4_add192_i113_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_398to400_bb4__26_i49_0_valid_out_NO_SHIFT_REG;
 logic rnode_398to400_bb4__26_i49_0_stall_in_NO_SHIFT_REG;
 logic rnode_398to400_bb4__26_i49_0_NO_SHIFT_REG;
 logic rnode_398to400_bb4__26_i49_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic rnode_398to400_bb4__26_i49_0_reg_400_NO_SHIFT_REG;
 logic rnode_398to400_bb4__26_i49_0_valid_out_reg_400_NO_SHIFT_REG;
 logic rnode_398to400_bb4__26_i49_0_stall_in_reg_400_NO_SHIFT_REG;
 logic rnode_398to400_bb4__26_i49_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_398to400_bb4__26_i49_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to400_bb4__26_i49_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to400_bb4__26_i49_0_stall_in_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_398to400_bb4__26_i49_0_valid_out_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_398to400_bb4__26_i49_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in(rnode_397to398_bb4__26_i49_0_NO_SHIFT_REG),
	.data_out(rnode_398to400_bb4__26_i49_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_398to400_bb4__26_i49_0_reg_400_fifo.DEPTH = 2;
defparam rnode_398to400_bb4__26_i49_0_reg_400_fifo.DATA_WIDTH = 1;
defparam rnode_398to400_bb4__26_i49_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to400_bb4__26_i49_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_398to400_bb4__26_i49_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4__26_i49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_398to400_bb4__26_i49_0_NO_SHIFT_REG = rnode_398to400_bb4__26_i49_0_reg_400_NO_SHIFT_REG;
assign rnode_398to400_bb4__26_i49_0_stall_in_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_398to400_bb4__26_i49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i_stall_local;
wire [31:0] local_bb4_reduction_1_i;

assign local_bb4_reduction_1_i = ((local_bb4_lnot_ext314_i & 32'h1) & (local_bb4_lor_ext_i & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_399to400_bb4_var__u98_0_valid_out_NO_SHIFT_REG;
 logic rnode_399to400_bb4_var__u98_0_stall_in_NO_SHIFT_REG;
 logic rnode_399to400_bb4_var__u98_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4_var__u98_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic rnode_399to400_bb4_var__u98_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_var__u98_0_valid_out_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_var__u98_0_stall_in_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_var__u98_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_399to400_bb4_var__u98_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to400_bb4_var__u98_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to400_bb4_var__u98_0_stall_in_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_399to400_bb4_var__u98_0_valid_out_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_399to400_bb4_var__u98_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in(rnode_398to399_bb4_var__u98_0_NO_SHIFT_REG),
	.data_out(rnode_399to400_bb4_var__u98_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_399to400_bb4_var__u98_0_reg_400_fifo.DEPTH = 1;
defparam rnode_399to400_bb4_var__u98_0_reg_400_fifo.DATA_WIDTH = 1;
defparam rnode_399to400_bb4_var__u98_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to400_bb4_var__u98_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_399to400_bb4_var__u98_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4_var__u98_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_var__u98_0_NO_SHIFT_REG = rnode_399to400_bb4_var__u98_0_reg_400_NO_SHIFT_REG;
assign rnode_399to400_bb4_var__u98_0_stall_in_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_var__u98_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_398to399_bb4_and193_i114_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and193_i114_0_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and193_i114_1_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and193_i114_2_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and193_i114_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_valid_out_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_stall_in_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and193_i114_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_398to399_bb4_and193_i114_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to399_bb4_and193_i114_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to399_bb4_and193_i114_0_stall_in_0_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_398to399_bb4_and193_i114_0_valid_out_0_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_398to399_bb4_and193_i114_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in((local_bb4_and193_i114 & 32'hFFFFFFF)),
	.data_out(rnode_398to399_bb4_and193_i114_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_398to399_bb4_and193_i114_0_reg_399_fifo.DEPTH = 1;
defparam rnode_398to399_bb4_and193_i114_0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_398to399_bb4_and193_i114_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to399_bb4_and193_i114_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_398to399_bb4_and193_i114_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and193_i114_stall_in = 1'b0;
assign rnode_398to399_bb4_and193_i114_0_stall_in_0_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and193_i114_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4_and193_i114_0_NO_SHIFT_REG = rnode_398to399_bb4_and193_i114_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4_and193_i114_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4_and193_i114_1_NO_SHIFT_REG = rnode_398to399_bb4_and193_i114_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4_and193_i114_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4_and193_i114_2_NO_SHIFT_REG = rnode_398to399_bb4_and193_i114_0_reg_399_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_398to399_bb4_and195_i115_0_valid_out_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and195_i115_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and195_i115_0_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and195_i115_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and195_i115_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and195_i115_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and195_i115_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and195_i115_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_398to399_bb4_and195_i115_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to399_bb4_and195_i115_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to399_bb4_and195_i115_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_398to399_bb4_and195_i115_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_398to399_bb4_and195_i115_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in((local_bb4_and195_i115 & 32'h1F)),
	.data_out(rnode_398to399_bb4_and195_i115_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_398to399_bb4_and195_i115_0_reg_399_fifo.DEPTH = 1;
defparam rnode_398to399_bb4_and195_i115_0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_398to399_bb4_and195_i115_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to399_bb4_and195_i115_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_398to399_bb4_and195_i115_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and195_i115_stall_in = 1'b0;
assign rnode_398to399_bb4_and195_i115_0_NO_SHIFT_REG = rnode_398to399_bb4_and195_i115_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4_and195_i115_0_stall_in_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and195_i115_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_398to399_bb4_and198_i116_0_valid_out_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and198_i116_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and198_i116_0_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and198_i116_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_and198_i116_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and198_i116_0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and198_i116_0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_and198_i116_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_398to399_bb4_and198_i116_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to399_bb4_and198_i116_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to399_bb4_and198_i116_0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_398to399_bb4_and198_i116_0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_398to399_bb4_and198_i116_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in((local_bb4_and198_i116 & 32'h1)),
	.data_out(rnode_398to399_bb4_and198_i116_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_398to399_bb4_and198_i116_0_reg_399_fifo.DEPTH = 1;
defparam rnode_398to399_bb4_and198_i116_0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_398to399_bb4_and198_i116_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to399_bb4_and198_i116_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_398to399_bb4_and198_i116_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and198_i116_stall_in = 1'b0;
assign rnode_398to399_bb4_and198_i116_0_NO_SHIFT_REG = rnode_398to399_bb4_and198_i116_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4_and198_i116_0_stall_in_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and198_i116_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i118_stall_local;
wire [31:0] local_bb4_shr_i_i118;

assign local_bb4_shr_i_i118 = ((local_bb4_and201_i117 & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4__26_i49_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_2_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_valid_out_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_stall_in_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4__26_i49_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4__26_i49_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4__26_i49_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4__26_i49_0_stall_in_0_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4__26_i49_0_valid_out_0_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4__26_i49_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(rnode_398to400_bb4__26_i49_0_NO_SHIFT_REG),
	.data_out(rnode_400to401_bb4__26_i49_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4__26_i49_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4__26_i49_0_reg_401_fifo.DATA_WIDTH = 1;
defparam rnode_400to401_bb4__26_i49_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4__26_i49_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4__26_i49_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_398to400_bb4__26_i49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__26_i49_0_stall_in_0_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__26_i49_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4__26_i49_0_NO_SHIFT_REG = rnode_400to401_bb4__26_i49_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4__26_i49_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4__26_i49_1_NO_SHIFT_REG = rnode_400to401_bb4__26_i49_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4__26_i49_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4__26_i49_2_NO_SHIFT_REG = rnode_400to401_bb4__26_i49_0_reg_401_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i_stall_local;
wire [31:0] local_bb4_reduction_2_i;

assign local_bb4_reduction_2_i = ((local_bb4_reduction_0_i & 32'h1) & (local_bb4_reduction_1_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr216_i139_stall_local;
wire [31:0] local_bb4_shr216_i139;

assign local_bb4_shr216_i139 = ((rnode_398to399_bb4_and193_i114_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i137_stall_local;
wire [31:0] local_bb4__pre_i137;

assign local_bb4__pre_i137 = ((rnode_398to399_bb4_and195_i115_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i119_stall_local;
wire [31:0] local_bb4_or_i_i119;

assign local_bb4_or_i_i119 = ((local_bb4_shr_i_i118 & 32'h3FFFFFF) | (local_bb4_and201_i117 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond292_i176_stall_local;
wire [31:0] local_bb4_cond292_i176;

assign local_bb4_cond292_i176 = (rnode_400to401_bb4__26_i49_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u106_stall_local;
wire [31:0] local_bb4_var__u106;

assign local_bb4_var__u106[31:1] = 31'h0;
assign local_bb4_var__u106[0] = rnode_400to401_bb4__26_i49_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add320_i_stall_local;
wire [31:0] local_bb4_add320_i;

assign local_bb4_add320_i = ((local_bb4_reduction_2_i & 32'h1) + local_bb4_or295_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or219_i140_stall_local;
wire [31:0] local_bb4_or219_i140;

assign local_bb4_or219_i140 = ((local_bb4_shr216_i139 & 32'h7FFFFFF) | (rnode_398to399_bb4_and198_i116_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool213_i138_stall_local;
wire local_bb4_tobool213_i138;

assign local_bb4_tobool213_i138 = ((local_bb4__pre_i137 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i120_stall_local;
wire [31:0] local_bb4_shr1_i_i120;

assign local_bb4_shr1_i_i120 = ((local_bb4_or_i_i119 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i186_stall_local;
wire [31:0] local_bb4_lnot_ext_i186;

assign local_bb4_lnot_ext_i186 = ((local_bb4_var__u106 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u107_stall_local;
wire [31:0] local_bb4_var__u107;

assign local_bb4_var__u107 = local_bb4_add320_i;

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i141_stall_local;
wire local_bb4__40_demorgan_i141;

assign local_bb4__40_demorgan_i141 = (rnode_397to399_bb4_cmp37_i36_0_NO_SHIFT_REG | local_bb4_tobool213_i138);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i143_stall_local;
wire local_bb4__42_i143;

assign local_bb4__42_i143 = (local_bb4_tobool213_i138 & local_bb4_not_cmp37_i142);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i121_stall_local;
wire [31:0] local_bb4_or2_i_i121;

assign local_bb4_or2_i_i121 = ((local_bb4_shr1_i_i120 & 32'h1FFFFFF) | (local_bb4_or_i_i119 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4___valid_out;
wire local_bb4___stall_in;
wire local_bb4___inputs_ready;
wire local_bb4___stall_local;
wire [31:0] local_bb4__;

assign local_bb4___inputs_ready = (rnode_395to396_bb4_c1_ene7_0_valid_out_0_NO_SHIFT_REG & rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_valid_out_NO_SHIFT_REG & rnode_394to396_bb4_and269_i_0_valid_out_NO_SHIFT_REG & rnode_395to396_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG & rnode_395to396_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG & rnode_395to396_bb4__26_i_0_valid_out_0_NO_SHIFT_REG & rnode_395to396_bb4__26_i_0_valid_out_1_NO_SHIFT_REG & rnode_395to396_bb4__47_i_0_valid_out_0_NO_SHIFT_REG & rnode_395to396_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG & rnode_395to396_bb4__26_i_0_valid_out_2_NO_SHIFT_REG & rnode_395to396_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG & rnode_395to396_bb4_shr271_i_0_valid_out_NO_SHIFT_REG & rnode_395to396_bb4__47_i_0_valid_out_1_NO_SHIFT_REG & rnode_395to396_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG & rnode_395to396_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4__ = (rnode_395to396_bb4_c1_ene7_0_NO_SHIFT_REG ? local_bb4_var__u107 : rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_NO_SHIFT_REG);
assign local_bb4___valid_out = 1'b1;
assign rnode_395to396_bb4_c1_ene7_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_sum_312_pop9_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_394to396_bb4_and269_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_resultSign_0_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_or2662_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__26_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__26_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__47_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_or2662_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__26_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_or2662_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_shr271_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4__47_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_cmp296_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_395to396_bb4_cmp299_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__43_i144_stall_local;
wire [31:0] local_bb4__43_i144;

assign local_bb4__43_i144 = (local_bb4__42_i143 ? 32'h0 : (local_bb4__pre_i137 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i122_stall_local;
wire [31:0] local_bb4_shr3_i_i122;

assign local_bb4_shr3_i_i122 = ((local_bb4_or2_i_i121 & 32'h7FFFFFF) >> 32'h4);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_396to397_bb4___0_valid_out_0_NO_SHIFT_REG;
 logic rnode_396to397_bb4___0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4___0_NO_SHIFT_REG;
 logic rnode_396to397_bb4___0_valid_out_1_NO_SHIFT_REG;
 logic rnode_396to397_bb4___0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4___1_NO_SHIFT_REG;
 logic rnode_396to397_bb4___0_reg_397_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_396to397_bb4___0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4___0_valid_out_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4___0_stall_in_0_reg_397_NO_SHIFT_REG;
 logic rnode_396to397_bb4___0_stall_out_reg_397_NO_SHIFT_REG;

acl_data_fifo rnode_396to397_bb4___0_reg_397_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_396to397_bb4___0_reg_397_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_396to397_bb4___0_stall_in_0_reg_397_NO_SHIFT_REG),
	.valid_out(rnode_396to397_bb4___0_valid_out_0_reg_397_NO_SHIFT_REG),
	.stall_out(rnode_396to397_bb4___0_stall_out_reg_397_NO_SHIFT_REG),
	.data_in(local_bb4__),
	.data_out(rnode_396to397_bb4___0_reg_397_NO_SHIFT_REG)
);

defparam rnode_396to397_bb4___0_reg_397_fifo.DEPTH = 1;
defparam rnode_396to397_bb4___0_reg_397_fifo.DATA_WIDTH = 32;
defparam rnode_396to397_bb4___0_reg_397_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_396to397_bb4___0_reg_397_fifo.IMPL = "shift_reg";

assign rnode_396to397_bb4___0_reg_397_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4___stall_in = 1'b0;
assign rnode_396to397_bb4___0_stall_in_0_reg_397_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4___0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4___0_NO_SHIFT_REG = rnode_396to397_bb4___0_reg_397_NO_SHIFT_REG;
assign rnode_396to397_bb4___0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4___1_NO_SHIFT_REG = rnode_396to397_bb4___0_reg_397_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i123_stall_local;
wire [31:0] local_bb4_or4_i_i123;

assign local_bb4_or4_i_i123 = ((local_bb4_shr3_i_i122 & 32'h7FFFFF) | (local_bb4_or2_i_i121 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire local_bb4_sum_312_push9___inputs_ready;
 reg local_bb4_sum_312_push9___valid_out_NO_SHIFT_REG;
wire local_bb4_sum_312_push9___stall_in;
wire local_bb4_sum_312_push9___output_regs_ready;
wire [31:0] local_bb4_sum_312_push9___result;
wire local_bb4_sum_312_push9___fu_valid_out;
wire local_bb4_sum_312_push9___fu_stall_out;
 reg [31:0] local_bb4_sum_312_push9___NO_SHIFT_REG;
wire local_bb4_sum_312_push9___causedstall;

acl_push local_bb4_sum_312_push9___feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_396to397_bb4_c1_ene8_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_396to397_bb4___0_NO_SHIFT_REG),
	.stall_out(local_bb4_sum_312_push9___fu_stall_out),
	.valid_in(SFC_3_VALID_396_397_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sum_312_push9___fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_sum_312_push9___result),
	.feedback_out(feedback_data_out_9),
	.feedback_valid_out(feedback_valid_out_9),
	.feedback_stall_in(feedback_stall_in_9)
);

defparam local_bb4_sum_312_push9___feedback.STALLFREE = 1;
defparam local_bb4_sum_312_push9___feedback.DATA_WIDTH = 32;
defparam local_bb4_sum_312_push9___feedback.FIFO_DEPTH = 9;
defparam local_bb4_sum_312_push9___feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_sum_312_push9___feedback.STYLE = "REGULAR";

assign local_bb4_sum_312_push9___inputs_ready = 1'b1;
assign local_bb4_sum_312_push9___output_regs_ready = 1'b1;
assign SFC_3_VALID_396_397_0_stall_in_1 = 1'b0;
assign rnode_396to397_bb4___0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_396to397_bb4_c1_ene8_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb4_sum_312_push9___causedstall = (SFC_3_VALID_396_397_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_sum_312_push9___NO_SHIFT_REG <= 'x;
		local_bb4_sum_312_push9___valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_sum_312_push9___output_regs_ready)
		begin
			local_bb4_sum_312_push9___NO_SHIFT_REG <= local_bb4_sum_312_push9___result;
			local_bb4_sum_312_push9___valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_sum_312_push9___stall_in))
			begin
				local_bb4_sum_312_push9___valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_397to398_bb4___0_valid_out_NO_SHIFT_REG;
 logic rnode_397to398_bb4___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb4___0_NO_SHIFT_REG;
 logic rnode_397to398_bb4___0_reg_398_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_397to398_bb4___0_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4___0_valid_out_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4___0_stall_in_reg_398_NO_SHIFT_REG;
 logic rnode_397to398_bb4___0_stall_out_reg_398_NO_SHIFT_REG;

acl_data_fifo rnode_397to398_bb4___0_reg_398_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_397to398_bb4___0_reg_398_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_397to398_bb4___0_stall_in_reg_398_NO_SHIFT_REG),
	.valid_out(rnode_397to398_bb4___0_valid_out_reg_398_NO_SHIFT_REG),
	.stall_out(rnode_397to398_bb4___0_stall_out_reg_398_NO_SHIFT_REG),
	.data_in(rnode_396to397_bb4___1_NO_SHIFT_REG),
	.data_out(rnode_397to398_bb4___0_reg_398_NO_SHIFT_REG)
);

defparam rnode_397to398_bb4___0_reg_398_fifo.DEPTH = 1;
defparam rnode_397to398_bb4___0_reg_398_fifo.DATA_WIDTH = 32;
defparam rnode_397to398_bb4___0_reg_398_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_397to398_bb4___0_reg_398_fifo.IMPL = "shift_reg";

assign rnode_397to398_bb4___0_reg_398_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_396to397_bb4___0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_397to398_bb4___0_NO_SHIFT_REG = rnode_397to398_bb4___0_reg_398_NO_SHIFT_REG;
assign rnode_397to398_bb4___0_stall_in_reg_398_NO_SHIFT_REG = 1'b0;
assign rnode_397to398_bb4___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i124_stall_local;
wire [31:0] local_bb4_shr5_i_i124;

assign local_bb4_shr5_i_i124 = ((local_bb4_or4_i_i123 & 32'h7FFFFFF) >> 32'h8);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_398to399_bb4_sum_312_push9___0_valid_out_NO_SHIFT_REG;
 logic rnode_398to399_bb4_sum_312_push9___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_sum_312_push9___0_NO_SHIFT_REG;
 logic rnode_398to399_bb4_sum_312_push9___0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4_sum_312_push9___0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_sum_312_push9___0_valid_out_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_sum_312_push9___0_stall_in_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4_sum_312_push9___0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_398to399_bb4_sum_312_push9___0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to399_bb4_sum_312_push9___0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to399_bb4_sum_312_push9___0_stall_in_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_398to399_bb4_sum_312_push9___0_valid_out_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_398to399_bb4_sum_312_push9___0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in(local_bb4_sum_312_push9___NO_SHIFT_REG),
	.data_out(rnode_398to399_bb4_sum_312_push9___0_reg_399_NO_SHIFT_REG)
);

defparam rnode_398to399_bb4_sum_312_push9___0_reg_399_fifo.DEPTH = 1;
defparam rnode_398to399_bb4_sum_312_push9___0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_398to399_bb4_sum_312_push9___0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to399_bb4_sum_312_push9___0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_398to399_bb4_sum_312_push9___0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_sum_312_push9___stall_in = 1'b0;
assign rnode_398to399_bb4_sum_312_push9___0_NO_SHIFT_REG = rnode_398to399_bb4_sum_312_push9___0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4_sum_312_push9___0_stall_in_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_sum_312_push9___0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_398to402_bb4___0_valid_out_NO_SHIFT_REG;
 logic rnode_398to402_bb4___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_398to402_bb4___0_NO_SHIFT_REG;
 logic rnode_398to402_bb4___0_reg_402_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_398to402_bb4___0_reg_402_NO_SHIFT_REG;
 logic rnode_398to402_bb4___0_valid_out_reg_402_NO_SHIFT_REG;
 logic rnode_398to402_bb4___0_stall_in_reg_402_NO_SHIFT_REG;
 logic rnode_398to402_bb4___0_stall_out_reg_402_NO_SHIFT_REG;

acl_data_fifo rnode_398to402_bb4___0_reg_402_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to402_bb4___0_reg_402_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to402_bb4___0_stall_in_reg_402_NO_SHIFT_REG),
	.valid_out(rnode_398to402_bb4___0_valid_out_reg_402_NO_SHIFT_REG),
	.stall_out(rnode_398to402_bb4___0_stall_out_reg_402_NO_SHIFT_REG),
	.data_in(rnode_397to398_bb4___0_NO_SHIFT_REG),
	.data_out(rnode_398to402_bb4___0_reg_402_NO_SHIFT_REG)
);

defparam rnode_398to402_bb4___0_reg_402_fifo.DEPTH = 4;
defparam rnode_398to402_bb4___0_reg_402_fifo.DATA_WIDTH = 32;
defparam rnode_398to402_bb4___0_reg_402_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to402_bb4___0_reg_402_fifo.IMPL = "shift_reg";

assign rnode_398to402_bb4___0_reg_402_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_397to398_bb4___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_398to402_bb4___0_NO_SHIFT_REG = rnode_398to402_bb4___0_reg_402_NO_SHIFT_REG;
assign rnode_398to402_bb4___0_stall_in_reg_402_NO_SHIFT_REG = 1'b0;
assign rnode_398to402_bb4___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i125_stall_local;
wire [31:0] local_bb4_or6_i_i125;

assign local_bb4_or6_i_i125 = ((local_bb4_shr5_i_i124 & 32'h7FFFF) | (local_bb4_or4_i_i123 & 32'h7FFFFFF));

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_399to402_bb4_sum_312_push9___0_valid_out_NO_SHIFT_REG;
 logic rnode_399to402_bb4_sum_312_push9___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_399to402_bb4_sum_312_push9___0_NO_SHIFT_REG;
 logic rnode_399to402_bb4_sum_312_push9___0_reg_402_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_399to402_bb4_sum_312_push9___0_reg_402_NO_SHIFT_REG;
 logic rnode_399to402_bb4_sum_312_push9___0_valid_out_reg_402_NO_SHIFT_REG;
 logic rnode_399to402_bb4_sum_312_push9___0_stall_in_reg_402_NO_SHIFT_REG;
 logic rnode_399to402_bb4_sum_312_push9___0_stall_out_reg_402_NO_SHIFT_REG;

acl_data_fifo rnode_399to402_bb4_sum_312_push9___0_reg_402_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to402_bb4_sum_312_push9___0_reg_402_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to402_bb4_sum_312_push9___0_stall_in_reg_402_NO_SHIFT_REG),
	.valid_out(rnode_399to402_bb4_sum_312_push9___0_valid_out_reg_402_NO_SHIFT_REG),
	.stall_out(rnode_399to402_bb4_sum_312_push9___0_stall_out_reg_402_NO_SHIFT_REG),
	.data_in(rnode_398to399_bb4_sum_312_push9___0_NO_SHIFT_REG),
	.data_out(rnode_399to402_bb4_sum_312_push9___0_reg_402_NO_SHIFT_REG)
);

defparam rnode_399to402_bb4_sum_312_push9___0_reg_402_fifo.DEPTH = 3;
defparam rnode_399to402_bb4_sum_312_push9___0_reg_402_fifo.DATA_WIDTH = 32;
defparam rnode_399to402_bb4_sum_312_push9___0_reg_402_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to402_bb4_sum_312_push9___0_reg_402_fifo.IMPL = "shift_reg";

assign rnode_399to402_bb4_sum_312_push9___0_reg_402_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4_sum_312_push9___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_399to402_bb4_sum_312_push9___0_NO_SHIFT_REG = rnode_399to402_bb4_sum_312_push9___0_reg_402_NO_SHIFT_REG;
assign rnode_399to402_bb4_sum_312_push9___0_stall_in_reg_402_NO_SHIFT_REG = 1'b0;
assign rnode_399to402_bb4_sum_312_push9___0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_402to403_bb4___0_valid_out_0_NO_SHIFT_REG;
 logic rnode_402to403_bb4___0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4___0_NO_SHIFT_REG;
 logic rnode_402to403_bb4___0_valid_out_1_NO_SHIFT_REG;
 logic rnode_402to403_bb4___0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4___1_NO_SHIFT_REG;
 logic rnode_402to403_bb4___0_reg_403_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4___0_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4___0_valid_out_0_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4___0_stall_in_0_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4___0_stall_out_reg_403_NO_SHIFT_REG;

acl_data_fifo rnode_402to403_bb4___0_reg_403_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_402to403_bb4___0_reg_403_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_402to403_bb4___0_stall_in_0_reg_403_NO_SHIFT_REG),
	.valid_out(rnode_402to403_bb4___0_valid_out_0_reg_403_NO_SHIFT_REG),
	.stall_out(rnode_402to403_bb4___0_stall_out_reg_403_NO_SHIFT_REG),
	.data_in(rnode_398to402_bb4___0_NO_SHIFT_REG),
	.data_out(rnode_402to403_bb4___0_reg_403_NO_SHIFT_REG)
);

defparam rnode_402to403_bb4___0_reg_403_fifo.DEPTH = 1;
defparam rnode_402to403_bb4___0_reg_403_fifo.DATA_WIDTH = 32;
defparam rnode_402to403_bb4___0_reg_403_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_402to403_bb4___0_reg_403_fifo.IMPL = "shift_reg";

assign rnode_402to403_bb4___0_reg_403_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_398to402_bb4___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_402to403_bb4___0_stall_in_0_reg_403_NO_SHIFT_REG = 1'b0;
assign rnode_402to403_bb4___0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_402to403_bb4___0_NO_SHIFT_REG = rnode_402to403_bb4___0_reg_403_NO_SHIFT_REG;
assign rnode_402to403_bb4___0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_402to403_bb4___1_NO_SHIFT_REG = rnode_402to403_bb4___0_reg_403_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i126_stall_local;
wire [31:0] local_bb4_shr7_i_i126;

assign local_bb4_shr7_i_i126 = ((local_bb4_or6_i_i125 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i127_stall_local;
wire [31:0] local_bb4_or6_masked_i_i127;

assign local_bb4_or6_masked_i_i127 = ((local_bb4_or6_i_i125 & 32'h7FFFFFF) & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_402to403_bb4_sum_312_push9___0_valid_out_NO_SHIFT_REG;
 logic rnode_402to403_bb4_sum_312_push9___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4_sum_312_push9___0_NO_SHIFT_REG;
 logic rnode_402to403_bb4_sum_312_push9___0_reg_403_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4_sum_312_push9___0_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4_sum_312_push9___0_valid_out_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4_sum_312_push9___0_stall_in_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4_sum_312_push9___0_stall_out_reg_403_NO_SHIFT_REG;

acl_data_fifo rnode_402to403_bb4_sum_312_push9___0_reg_403_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_402to403_bb4_sum_312_push9___0_reg_403_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_402to403_bb4_sum_312_push9___0_stall_in_reg_403_NO_SHIFT_REG),
	.valid_out(rnode_402to403_bb4_sum_312_push9___0_valid_out_reg_403_NO_SHIFT_REG),
	.stall_out(rnode_402to403_bb4_sum_312_push9___0_stall_out_reg_403_NO_SHIFT_REG),
	.data_in(rnode_399to402_bb4_sum_312_push9___0_NO_SHIFT_REG),
	.data_out(rnode_402to403_bb4_sum_312_push9___0_reg_403_NO_SHIFT_REG)
);

defparam rnode_402to403_bb4_sum_312_push9___0_reg_403_fifo.DEPTH = 1;
defparam rnode_402to403_bb4_sum_312_push9___0_reg_403_fifo.DATA_WIDTH = 32;
defparam rnode_402to403_bb4_sum_312_push9___0_reg_403_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_402to403_bb4_sum_312_push9___0_reg_403_fifo.IMPL = "shift_reg";

assign rnode_402to403_bb4_sum_312_push9___0_reg_403_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_399to402_bb4_sum_312_push9___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_402to403_bb4_sum_312_push9___0_NO_SHIFT_REG = rnode_402to403_bb4_sum_312_push9___0_reg_403_NO_SHIFT_REG;
assign rnode_402to403_bb4_sum_312_push9___0_stall_in_reg_403_NO_SHIFT_REG = 1'b0;
assign rnode_402to403_bb4_sum_312_push9___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4____valid_out;
wire local_bb4____stall_in;
wire local_bb4____inputs_ready;
wire local_bb4____stall_local;
 reg [31:0] ffwd_11_0_reg_NO_SHIFT_REG;

assign local_bb4____inputs_ready = (SFC_3_VALID_402_403_0_valid_out_1_NO_SHIFT_REG & rnode_402to403_bb4___0_valid_out_0_NO_SHIFT_REG);
assign ffwd_11_0 = ffwd_11_0_reg_NO_SHIFT_REG;
assign local_bb4____valid_out = 1'b1;
assign SFC_3_VALID_402_403_0_stall_in_1 = 1'b0;
assign rnode_402to403_bb4___0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock)
begin
	if ((1'b1 & SFC_3_VALID_402_403_0_NO_SHIFT_REG))
	begin
		ffwd_11_0_reg_NO_SHIFT_REG <= rnode_402to403_bb4___0_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_exi1_stall_local;
wire [95:0] local_bb4_c1_exi1;

assign local_bb4_c1_exi1[31:0] = 32'bx;
assign local_bb4_c1_exi1[63:32] = rnode_402to403_bb4___1_NO_SHIFT_REG;
assign local_bb4_c1_exi1[95:64] = 32'bx;

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i128_stall_local;
wire [31:0] local_bb4_neg_i_i128;

assign local_bb4_neg_i_i128 = ((local_bb4_or6_masked_i_i127 & 32'h7FFFFFF) | (local_bb4_shr7_i_i126 & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i129_stall_local;
wire [31:0] local_bb4_and_i_i129;

assign local_bb4_and_i_i129 = ((local_bb4_neg_i_i128 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i129_valid_out;
wire local_bb4__and_i_i129_stall_in;
wire local_bb4__and_i_i129_inputs_ready;
wire local_bb4__and_i_i129_stall_local;
wire [31:0] local_bb4__and_i_i129;

thirtysix_six_comp local_bb4__and_i_i129_popcnt_instance (
	.data((local_bb4_and_i_i129 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i129)
);


assign local_bb4__and_i_i129_inputs_ready = rnode_397to398_bb4_add192_i113_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i129_valid_out = 1'b1;
assign rnode_397to398_bb4_add192_i113_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_398to399_bb4__and_i_i129_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4__and_i_i129_0_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4__and_i_i129_1_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4__and_i_i129_2_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_reg_399_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_398to399_bb4__and_i_i129_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_valid_out_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_stall_in_0_reg_399_NO_SHIFT_REG;
 logic rnode_398to399_bb4__and_i_i129_0_stall_out_reg_399_NO_SHIFT_REG;

acl_data_fifo rnode_398to399_bb4__and_i_i129_0_reg_399_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_398to399_bb4__and_i_i129_0_reg_399_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_398to399_bb4__and_i_i129_0_stall_in_0_reg_399_NO_SHIFT_REG),
	.valid_out(rnode_398to399_bb4__and_i_i129_0_valid_out_0_reg_399_NO_SHIFT_REG),
	.stall_out(rnode_398to399_bb4__and_i_i129_0_stall_out_reg_399_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i129 & 32'h3F)),
	.data_out(rnode_398to399_bb4__and_i_i129_0_reg_399_NO_SHIFT_REG)
);

defparam rnode_398to399_bb4__and_i_i129_0_reg_399_fifo.DEPTH = 1;
defparam rnode_398to399_bb4__and_i_i129_0_reg_399_fifo.DATA_WIDTH = 32;
defparam rnode_398to399_bb4__and_i_i129_0_reg_399_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_398to399_bb4__and_i_i129_0_reg_399_fifo.IMPL = "shift_reg";

assign rnode_398to399_bb4__and_i_i129_0_reg_399_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i129_stall_in = 1'b0;
assign rnode_398to399_bb4__and_i_i129_0_stall_in_0_reg_399_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4__and_i_i129_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4__and_i_i129_0_NO_SHIFT_REG = rnode_398to399_bb4__and_i_i129_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4__and_i_i129_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4__and_i_i129_1_NO_SHIFT_REG = rnode_398to399_bb4__and_i_i129_0_reg_399_NO_SHIFT_REG;
assign rnode_398to399_bb4__and_i_i129_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_398to399_bb4__and_i_i129_2_NO_SHIFT_REG = rnode_398to399_bb4__and_i_i129_0_reg_399_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i130_stall_local;
wire [31:0] local_bb4_and9_i_i130;

assign local_bb4_and9_i_i130 = ((rnode_398to399_bb4__and_i_i129_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and203_i131_stall_local;
wire [31:0] local_bb4_and203_i131;

assign local_bb4_and203_i131 = ((rnode_398to399_bb4__and_i_i129_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i133_stall_local;
wire [31:0] local_bb4_and206_i133;

assign local_bb4_and206_i133 = ((rnode_398to399_bb4__and_i_i129_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_sub239_i152_stall_local;
wire [31:0] local_bb4_sub239_i152;

assign local_bb4_sub239_i152 = (32'h0 - (local_bb4_and9_i_i130 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl204_i132_stall_local;
wire [31:0] local_bb4_shl204_i132;

assign local_bb4_shl204_i132 = ((rnode_398to399_bb4_and193_i114_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and203_i131 & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb4_cond244_i153_stall_local;
wire [31:0] local_bb4_cond244_i153;

assign local_bb4_cond244_i153 = (rnode_397to399_bb4_cmp37_i36_2_NO_SHIFT_REG ? local_bb4_sub239_i152 : (local_bb4__43_i144 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and205_i134_stall_local;
wire [31:0] local_bb4_and205_i134;

assign local_bb4_and205_i134 = (local_bb4_shl204_i132 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_add245_i154_stall_local;
wire [31:0] local_bb4_add245_i154;

assign local_bb4_add245_i154 = (local_bb4_cond244_i153 + (rnode_397to399_bb4_and17_i25_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i156_stall_local;
wire [31:0] local_bb4_fold_i156;

assign local_bb4_fold_i156 = (local_bb4_cond244_i153 + (rnode_397to399_bb4_shr16_i24_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl207_i135_stall_local;
wire [31:0] local_bb4_shl207_i135;

assign local_bb4_shl207_i135 = ((local_bb4_and205_i134 & 32'h7FFFFFF) << (local_bb4_and206_i133 & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i157_stall_local;
wire [31:0] local_bb4_and250_i157;

assign local_bb4_and250_i157 = (local_bb4_fold_i156 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and269_i168_stall_local;
wire [31:0] local_bb4_and269_i168;

assign local_bb4_and269_i168 = (local_bb4_fold_i156 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and208_i136_stall_local;
wire [31:0] local_bb4_and208_i136;

assign local_bb4_and208_i136 = (local_bb4_shl207_i135 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__44_i145_stall_local;
wire [31:0] local_bb4__44_i145;

assign local_bb4__44_i145 = (local_bb4__40_demorgan_i141 ? (local_bb4_and208_i136 & 32'h7FFFFFF) : (local_bb4_or219_i140 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i157_valid_out;
wire local_bb4_and250_i157_stall_in;
wire local_bb4_and269_i168_valid_out;
wire local_bb4_and269_i168_stall_in;
wire local_bb4_add245_i154_valid_out;
wire local_bb4_add245_i154_stall_in;
wire local_bb4__45_i146_valid_out;
wire local_bb4__45_i146_stall_in;
wire local_bb4_not_cmp37_i142_valid_out_1;
wire local_bb4_not_cmp37_i142_stall_in_1;
wire local_bb4__45_i146_inputs_ready;
wire local_bb4__45_i146_stall_local;
wire [31:0] local_bb4__45_i146;

assign local_bb4__45_i146_inputs_ready = (rnode_397to399_bb4_shr16_i24_0_valid_out_NO_SHIFT_REG & rnode_397to399_bb4_and17_i25_0_valid_out_NO_SHIFT_REG & rnode_397to399_bb4_cmp37_i36_0_valid_out_2_NO_SHIFT_REG & rnode_397to399_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG & rnode_398to399_bb4_and193_i114_0_valid_out_2_NO_SHIFT_REG & rnode_397to399_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG & rnode_398to399_bb4_and195_i115_0_valid_out_NO_SHIFT_REG & rnode_398to399_bb4_and193_i114_0_valid_out_1_NO_SHIFT_REG & rnode_398to399_bb4_and198_i116_0_valid_out_NO_SHIFT_REG & rnode_398to399_bb4_and193_i114_0_valid_out_0_NO_SHIFT_REG & rnode_398to399_bb4__and_i_i129_0_valid_out_1_NO_SHIFT_REG & rnode_398to399_bb4__and_i_i129_0_valid_out_2_NO_SHIFT_REG & rnode_398to399_bb4__and_i_i129_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i146 = (local_bb4__42_i143 ? (rnode_398to399_bb4_and193_i114_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i145 & 32'h7FFFFFF));
assign local_bb4_and250_i157_valid_out = 1'b1;
assign local_bb4_and269_i168_valid_out = 1'b1;
assign local_bb4_add245_i154_valid_out = 1'b1;
assign local_bb4__45_i146_valid_out = 1'b1;
assign local_bb4_not_cmp37_i142_valid_out_1 = 1'b1;
assign rnode_397to399_bb4_shr16_i24_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_and17_i25_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_cmp37_i36_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and193_i114_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_397to399_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and195_i115_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and193_i114_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and198_i116_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4_and193_i114_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4__and_i_i129_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4__and_i_i129_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_398to399_bb4__and_i_i129_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_399to400_bb4_and250_i157_0_valid_out_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and250_i157_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4_and250_i157_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and250_i157_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4_and250_i157_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and250_i157_0_valid_out_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and250_i157_0_stall_in_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_and250_i157_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_399to400_bb4_and250_i157_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to400_bb4_and250_i157_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to400_bb4_and250_i157_0_stall_in_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_399to400_bb4_and250_i157_0_valid_out_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_399to400_bb4_and250_i157_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in((local_bb4_and250_i157 & 32'hFF)),
	.data_out(rnode_399to400_bb4_and250_i157_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_399to400_bb4_and250_i157_0_reg_400_fifo.DEPTH = 1;
defparam rnode_399to400_bb4_and250_i157_0_reg_400_fifo.DATA_WIDTH = 32;
defparam rnode_399to400_bb4_and250_i157_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to400_bb4_and250_i157_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_399to400_bb4_and250_i157_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and250_i157_stall_in = 1'b0;
assign rnode_399to400_bb4_and250_i157_0_NO_SHIFT_REG = rnode_399to400_bb4_and250_i157_0_reg_400_NO_SHIFT_REG;
assign rnode_399to400_bb4_and250_i157_0_stall_in_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_and250_i157_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_399to401_bb4_and269_i168_0_valid_out_NO_SHIFT_REG;
 logic rnode_399to401_bb4_and269_i168_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_399to401_bb4_and269_i168_0_NO_SHIFT_REG;
 logic rnode_399to401_bb4_and269_i168_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_399to401_bb4_and269_i168_0_reg_401_NO_SHIFT_REG;
 logic rnode_399to401_bb4_and269_i168_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_399to401_bb4_and269_i168_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_399to401_bb4_and269_i168_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_399to401_bb4_and269_i168_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to401_bb4_and269_i168_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to401_bb4_and269_i168_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_399to401_bb4_and269_i168_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_399to401_bb4_and269_i168_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in((local_bb4_and269_i168 & 32'hFF800000)),
	.data_out(rnode_399to401_bb4_and269_i168_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_399to401_bb4_and269_i168_0_reg_401_fifo.DEPTH = 2;
defparam rnode_399to401_bb4_and269_i168_0_reg_401_fifo.DATA_WIDTH = 32;
defparam rnode_399to401_bb4_and269_i168_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to401_bb4_and269_i168_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_399to401_bb4_and269_i168_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and269_i168_stall_in = 1'b0;
assign rnode_399to401_bb4_and269_i168_0_NO_SHIFT_REG = rnode_399to401_bb4_and269_i168_0_reg_401_NO_SHIFT_REG;
assign rnode_399to401_bb4_and269_i168_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_399to401_bb4_and269_i168_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_399to400_bb4_add245_i154_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4_add245_i154_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4_add245_i154_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4_add245_i154_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_399to400_bb4_add245_i154_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4_add245_i154_1_NO_SHIFT_REG;
 logic rnode_399to400_bb4_add245_i154_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4_add245_i154_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_add245_i154_0_valid_out_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_add245_i154_0_stall_in_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_add245_i154_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_399to400_bb4_add245_i154_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to400_bb4_add245_i154_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to400_bb4_add245_i154_0_stall_in_0_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_399to400_bb4_add245_i154_0_valid_out_0_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_399to400_bb4_add245_i154_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in(local_bb4_add245_i154),
	.data_out(rnode_399to400_bb4_add245_i154_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_399to400_bb4_add245_i154_0_reg_400_fifo.DEPTH = 1;
defparam rnode_399to400_bb4_add245_i154_0_reg_400_fifo.DATA_WIDTH = 32;
defparam rnode_399to400_bb4_add245_i154_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to400_bb4_add245_i154_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_399to400_bb4_add245_i154_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add245_i154_stall_in = 1'b0;
assign rnode_399to400_bb4_add245_i154_0_stall_in_0_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_add245_i154_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_399to400_bb4_add245_i154_0_NO_SHIFT_REG = rnode_399to400_bb4_add245_i154_0_reg_400_NO_SHIFT_REG;
assign rnode_399to400_bb4_add245_i154_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_399to400_bb4_add245_i154_1_NO_SHIFT_REG = rnode_399to400_bb4_add245_i154_0_reg_400_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_399to400_bb4__45_i146_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4__45_i146_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4__45_i146_1_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4__45_i146_2_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_399to400_bb4__45_i146_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_valid_out_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_stall_in_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4__45_i146_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_399to400_bb4__45_i146_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to400_bb4__45_i146_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to400_bb4__45_i146_0_stall_in_0_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_399to400_bb4__45_i146_0_valid_out_0_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_399to400_bb4__45_i146_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in((local_bb4__45_i146 & 32'hFFFFFFF)),
	.data_out(rnode_399to400_bb4__45_i146_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_399to400_bb4__45_i146_0_reg_400_fifo.DEPTH = 1;
defparam rnode_399to400_bb4__45_i146_0_reg_400_fifo.DATA_WIDTH = 32;
defparam rnode_399to400_bb4__45_i146_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to400_bb4__45_i146_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_399to400_bb4__45_i146_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i146_stall_in = 1'b0;
assign rnode_399to400_bb4__45_i146_0_stall_in_0_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4__45_i146_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_399to400_bb4__45_i146_0_NO_SHIFT_REG = rnode_399to400_bb4__45_i146_0_reg_400_NO_SHIFT_REG;
assign rnode_399to400_bb4__45_i146_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_399to400_bb4__45_i146_1_NO_SHIFT_REG = rnode_399to400_bb4__45_i146_0_reg_400_NO_SHIFT_REG;
assign rnode_399to400_bb4__45_i146_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_399to400_bb4__45_i146_2_NO_SHIFT_REG = rnode_399to400_bb4__45_i146_0_reg_400_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_399to400_bb4_not_cmp37_i142_0_valid_out_NO_SHIFT_REG;
 logic rnode_399to400_bb4_not_cmp37_i142_0_stall_in_NO_SHIFT_REG;
 logic rnode_399to400_bb4_not_cmp37_i142_0_NO_SHIFT_REG;
 logic rnode_399to400_bb4_not_cmp37_i142_0_reg_400_inputs_ready_NO_SHIFT_REG;
 logic rnode_399to400_bb4_not_cmp37_i142_0_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_not_cmp37_i142_0_valid_out_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_not_cmp37_i142_0_stall_in_reg_400_NO_SHIFT_REG;
 logic rnode_399to400_bb4_not_cmp37_i142_0_stall_out_reg_400_NO_SHIFT_REG;

acl_data_fifo rnode_399to400_bb4_not_cmp37_i142_0_reg_400_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_399to400_bb4_not_cmp37_i142_0_reg_400_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_399to400_bb4_not_cmp37_i142_0_stall_in_reg_400_NO_SHIFT_REG),
	.valid_out(rnode_399to400_bb4_not_cmp37_i142_0_valid_out_reg_400_NO_SHIFT_REG),
	.stall_out(rnode_399to400_bb4_not_cmp37_i142_0_stall_out_reg_400_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp37_i142),
	.data_out(rnode_399to400_bb4_not_cmp37_i142_0_reg_400_NO_SHIFT_REG)
);

defparam rnode_399to400_bb4_not_cmp37_i142_0_reg_400_fifo.DEPTH = 1;
defparam rnode_399to400_bb4_not_cmp37_i142_0_reg_400_fifo.DATA_WIDTH = 1;
defparam rnode_399to400_bb4_not_cmp37_i142_0_reg_400_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_399to400_bb4_not_cmp37_i142_0_reg_400_fifo.IMPL = "shift_reg";

assign rnode_399to400_bb4_not_cmp37_i142_0_reg_400_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp37_i142_stall_in_1 = 1'b0;
assign rnode_399to400_bb4_not_cmp37_i142_0_NO_SHIFT_REG = rnode_399to400_bb4_not_cmp37_i142_0_reg_400_NO_SHIFT_REG;
assign rnode_399to400_bb4_not_cmp37_i142_0_stall_in_reg_400_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_not_cmp37_i142_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i159_stall_local;
wire local_bb4_notrhs_i159;

assign local_bb4_notrhs_i159 = ((rnode_399to400_bb4_and250_i157_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl273_i169_stall_local;
wire [31:0] local_bb4_shl273_i169;

assign local_bb4_shl273_i169 = ((rnode_399to401_bb4_and269_i168_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and247_i155_stall_local;
wire [31:0] local_bb4_and247_i155;

assign local_bb4_and247_i155 = (rnode_399to400_bb4_add245_i154_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp258_i162_stall_local;
wire local_bb4_cmp258_i162;

assign local_bb4_cmp258_i162 = ($signed(rnode_399to400_bb4_add245_i154_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and225_i147_stall_local;
wire [31:0] local_bb4_and225_i147;

assign local_bb4_and225_i147 = ((rnode_399to400_bb4__45_i146_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i165_stall_local;
wire [31:0] local_bb4_and270_i165;

assign local_bb4_and270_i165 = ((rnode_399to400_bb4__45_i146_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr271_i166_valid_out;
wire local_bb4_shr271_i166_stall_in;
wire local_bb4_shr271_i166_inputs_ready;
wire local_bb4_shr271_i166_stall_local;
wire [31:0] local_bb4_shr271_i166;

assign local_bb4_shr271_i166_inputs_ready = rnode_399to400_bb4__45_i146_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr271_i166 = ((rnode_399to400_bb4__45_i146_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr271_i166_valid_out = 1'b1;
assign rnode_399to400_bb4__45_i146_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i158_stall_local;
wire local_bb4_notlhs_i158;

assign local_bb4_notlhs_i158 = ((local_bb4_and247_i155 & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_i148_stall_local;
wire local_bb4_cmp226_i148;

assign local_bb4_cmp226_i148 = ((local_bb4_and225_i147 & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i180_stall_local;
wire local_bb4_cmp296_i180;

assign local_bb4_cmp296_i180 = ((local_bb4_and270_i165 & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i180_valid_out;
wire local_bb4_cmp296_i180_stall_in;
wire local_bb4_cmp299_i181_valid_out;
wire local_bb4_cmp299_i181_stall_in;
wire local_bb4_cmp299_i181_inputs_ready;
wire local_bb4_cmp299_i181_stall_local;
wire local_bb4_cmp299_i181;

assign local_bb4_cmp299_i181_inputs_ready = rnode_399to400_bb4__45_i146_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp299_i181 = ((local_bb4_and270_i165 & 32'h7) == 32'h4);
assign local_bb4_cmp296_i180_valid_out = 1'b1;
assign local_bb4_cmp299_i181_valid_out = 1'b1;
assign rnode_399to400_bb4__45_i146_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4_shr271_i166_0_valid_out_NO_SHIFT_REG;
 logic rnode_400to401_bb4_shr271_i166_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_400to401_bb4_shr271_i166_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_shr271_i166_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_400to401_bb4_shr271_i166_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_shr271_i166_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_shr271_i166_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_shr271_i166_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4_shr271_i166_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4_shr271_i166_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4_shr271_i166_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4_shr271_i166_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4_shr271_i166_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in((local_bb4_shr271_i166 & 32'h1FFFFFF)),
	.data_out(rnode_400to401_bb4_shr271_i166_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4_shr271_i166_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4_shr271_i166_0_reg_401_fifo.DATA_WIDTH = 32;
defparam rnode_400to401_bb4_shr271_i166_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4_shr271_i166_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4_shr271_i166_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr271_i166_stall_in = 1'b0;
assign rnode_400to401_bb4_shr271_i166_0_NO_SHIFT_REG = rnode_400to401_bb4_shr271_i166_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_shr271_i166_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_shr271_i166_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i160_stall_local;
wire local_bb4_not__46_i160;

assign local_bb4_not__46_i160 = (local_bb4_notrhs_i159 | local_bb4_notlhs_i158);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_not_i149_stall_local;
wire local_bb4_cmp226_not_i149;

assign local_bb4_cmp226_not_i149 = (local_bb4_cmp226_i148 ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4_cmp296_i180_0_valid_out_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp296_i180_0_stall_in_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp296_i180_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp296_i180_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp296_i180_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp296_i180_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp296_i180_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp296_i180_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4_cmp296_i180_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4_cmp296_i180_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4_cmp296_i180_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4_cmp296_i180_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4_cmp296_i180_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(local_bb4_cmp296_i180),
	.data_out(rnode_400to401_bb4_cmp296_i180_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4_cmp296_i180_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4_cmp296_i180_0_reg_401_fifo.DATA_WIDTH = 1;
defparam rnode_400to401_bb4_cmp296_i180_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4_cmp296_i180_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4_cmp296_i180_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp296_i180_stall_in = 1'b0;
assign rnode_400to401_bb4_cmp296_i180_0_NO_SHIFT_REG = rnode_400to401_bb4_cmp296_i180_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_cmp296_i180_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_cmp296_i180_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4_cmp299_i181_0_valid_out_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp299_i181_0_stall_in_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp299_i181_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp299_i181_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp299_i181_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp299_i181_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp299_i181_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_cmp299_i181_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4_cmp299_i181_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4_cmp299_i181_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4_cmp299_i181_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4_cmp299_i181_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4_cmp299_i181_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(local_bb4_cmp299_i181),
	.data_out(rnode_400to401_bb4_cmp299_i181_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4_cmp299_i181_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4_cmp299_i181_0_reg_401_fifo.DATA_WIDTH = 1;
defparam rnode_400to401_bb4_cmp299_i181_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4_cmp299_i181_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4_cmp299_i181_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp299_i181_stall_in = 1'b0;
assign rnode_400to401_bb4_cmp299_i181_0_NO_SHIFT_REG = rnode_400to401_bb4_cmp299_i181_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_cmp299_i181_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_cmp299_i181_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and272_i167_stall_local;
wire [31:0] local_bb4_and272_i167;

assign local_bb4_and272_i167 = ((rnode_400to401_bb4_shr271_i166_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__47_i161_stall_local;
wire local_bb4__47_i161;

assign local_bb4__47_i161 = (local_bb4_cmp226_i148 | local_bb4_not__46_i160);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i150_stall_local;
wire local_bb4_brmerge12_i150;

assign local_bb4_brmerge12_i150 = (local_bb4_cmp226_not_i149 | rnode_399to400_bb4_not_cmp37_i142_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot262__i163_stall_local;
wire local_bb4_lnot262__i163;

assign local_bb4_lnot262__i163 = (local_bb4_cmp258_i162 & local_bb4_cmp226_not_i149);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29649_i184_stall_local;
wire [31:0] local_bb4_cmp29649_i184;

assign local_bb4_cmp29649_i184[31:1] = 31'h0;
assign local_bb4_cmp29649_i184[0] = rnode_400to401_bb4_cmp296_i180_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv300_i182_stall_local;
wire [31:0] local_bb4_conv300_i182;

assign local_bb4_conv300_i182[31:1] = 31'h0;
assign local_bb4_conv300_i182[0] = rnode_400to401_bb4_cmp299_i181_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or274_i170_stall_local;
wire [31:0] local_bb4_or274_i170;

assign local_bb4_or274_i170 = ((local_bb4_and272_i167 & 32'h7FFFFF) | (local_bb4_shl273_i169 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i151_stall_local;
wire [31:0] local_bb4_resultSign_0_i151;

assign local_bb4_resultSign_0_i151 = (local_bb4_brmerge12_i150 ? (rnode_399to400_bb4_and35_i34_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i151_valid_out;
wire local_bb4_resultSign_0_i151_stall_in;
wire local_bb4__47_i161_valid_out;
wire local_bb4__47_i161_stall_in;
wire local_bb4_or2662_i164_valid_out;
wire local_bb4_or2662_i164_stall_in;
wire local_bb4_or2662_i164_inputs_ready;
wire local_bb4_or2662_i164_stall_local;
wire local_bb4_or2662_i164;

assign local_bb4_or2662_i164_inputs_ready = (rnode_399to400_bb4_and35_i34_0_valid_out_NO_SHIFT_REG & rnode_399to400_bb4_not_cmp37_i142_0_valid_out_NO_SHIFT_REG & rnode_399to400_bb4_add245_i154_0_valid_out_0_NO_SHIFT_REG & rnode_399to400_bb4_and250_i157_0_valid_out_NO_SHIFT_REG & rnode_399to400_bb4__45_i146_0_valid_out_0_NO_SHIFT_REG & rnode_399to400_bb4_add245_i154_0_valid_out_1_NO_SHIFT_REG & rnode_399to400_bb4_var__u98_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2662_i164 = (rnode_399to400_bb4_var__u98_0_NO_SHIFT_REG | local_bb4_lnot262__i163);
assign local_bb4_resultSign_0_i151_valid_out = 1'b1;
assign local_bb4__47_i161_valid_out = 1'b1;
assign local_bb4_or2662_i164_valid_out = 1'b1;
assign rnode_399to400_bb4_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_not_cmp37_i142_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_add245_i154_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_and250_i157_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4__45_i146_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_add245_i154_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_399to400_bb4_var__u98_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4_resultSign_0_i151_0_valid_out_NO_SHIFT_REG;
 logic rnode_400to401_bb4_resultSign_0_i151_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_400to401_bb4_resultSign_0_i151_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_resultSign_0_i151_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_400to401_bb4_resultSign_0_i151_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_resultSign_0_i151_0_valid_out_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_resultSign_0_i151_0_stall_in_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_resultSign_0_i151_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4_resultSign_0_i151_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4_resultSign_0_i151_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4_resultSign_0_i151_0_stall_in_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4_resultSign_0_i151_0_valid_out_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4_resultSign_0_i151_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i151 & 32'h80000000)),
	.data_out(rnode_400to401_bb4_resultSign_0_i151_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4_resultSign_0_i151_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4_resultSign_0_i151_0_reg_401_fifo.DATA_WIDTH = 32;
defparam rnode_400to401_bb4_resultSign_0_i151_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4_resultSign_0_i151_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4_resultSign_0_i151_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i151_stall_in = 1'b0;
assign rnode_400to401_bb4_resultSign_0_i151_0_NO_SHIFT_REG = rnode_400to401_bb4_resultSign_0_i151_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_resultSign_0_i151_0_stall_in_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_resultSign_0_i151_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4__47_i161_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_valid_out_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_stall_in_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4__47_i161_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4__47_i161_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4__47_i161_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4__47_i161_0_stall_in_0_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4__47_i161_0_valid_out_0_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4__47_i161_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(local_bb4__47_i161),
	.data_out(rnode_400to401_bb4__47_i161_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4__47_i161_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4__47_i161_0_reg_401_fifo.DATA_WIDTH = 1;
defparam rnode_400to401_bb4__47_i161_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4__47_i161_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4__47_i161_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i161_stall_in = 1'b0;
assign rnode_400to401_bb4__47_i161_0_stall_in_0_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__47_i161_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4__47_i161_0_NO_SHIFT_REG = rnode_400to401_bb4__47_i161_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4__47_i161_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4__47_i161_1_NO_SHIFT_REG = rnode_400to401_bb4__47_i161_0_reg_401_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_400to401_bb4_or2662_i164_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_1_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_2_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_reg_401_inputs_ready_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_valid_out_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_stall_in_0_reg_401_NO_SHIFT_REG;
 logic rnode_400to401_bb4_or2662_i164_0_stall_out_reg_401_NO_SHIFT_REG;

acl_data_fifo rnode_400to401_bb4_or2662_i164_0_reg_401_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_400to401_bb4_or2662_i164_0_reg_401_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_400to401_bb4_or2662_i164_0_stall_in_0_reg_401_NO_SHIFT_REG),
	.valid_out(rnode_400to401_bb4_or2662_i164_0_valid_out_0_reg_401_NO_SHIFT_REG),
	.stall_out(rnode_400to401_bb4_or2662_i164_0_stall_out_reg_401_NO_SHIFT_REG),
	.data_in(local_bb4_or2662_i164),
	.data_out(rnode_400to401_bb4_or2662_i164_0_reg_401_NO_SHIFT_REG)
);

defparam rnode_400to401_bb4_or2662_i164_0_reg_401_fifo.DEPTH = 1;
defparam rnode_400to401_bb4_or2662_i164_0_reg_401_fifo.DATA_WIDTH = 1;
defparam rnode_400to401_bb4_or2662_i164_0_reg_401_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_400to401_bb4_or2662_i164_0_reg_401_fifo.IMPL = "shift_reg";

assign rnode_400to401_bb4_or2662_i164_0_reg_401_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2662_i164_stall_in = 1'b0;
assign rnode_400to401_bb4_or2662_i164_0_stall_in_0_reg_401_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_or2662_i164_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4_or2662_i164_0_NO_SHIFT_REG = rnode_400to401_bb4_or2662_i164_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_or2662_i164_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4_or2662_i164_1_NO_SHIFT_REG = rnode_400to401_bb4_or2662_i164_0_reg_401_NO_SHIFT_REG;
assign rnode_400to401_bb4_or2662_i164_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_400to401_bb4_or2662_i164_2_NO_SHIFT_REG = rnode_400to401_bb4_or2662_i164_0_reg_401_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i171_stall_local;
wire [31:0] local_bb4_or275_i171;

assign local_bb4_or275_i171 = ((local_bb4_or274_i170 & 32'h7FFFFFFF) | (rnode_400to401_bb4_resultSign_0_i151_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u108_stall_local;
wire [31:0] local_bb4_var__u108;

assign local_bb4_var__u108[31:1] = 31'h0;
assign local_bb4_var__u108[0] = rnode_400to401_bb4__47_i161_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2804_i172_stall_local;
wire local_bb4_or2804_i172;

assign local_bb4_or2804_i172 = (rnode_400to401_bb4__47_i161_0_NO_SHIFT_REG | rnode_400to401_bb4_or2662_i164_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2875_i174_stall_local;
wire local_bb4_or2875_i174;

assign local_bb4_or2875_i174 = (rnode_400to401_bb4_or2662_i164_1_NO_SHIFT_REG | rnode_400to401_bb4__26_i49_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u109_stall_local;
wire [31:0] local_bb4_var__u109;

assign local_bb4_var__u109[31:1] = 31'h0;
assign local_bb4_var__u109[0] = rnode_400to401_bb4_or2662_i164_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext314_i188_stall_local;
wire [31:0] local_bb4_lnot_ext314_i188;

assign local_bb4_lnot_ext314_i188 = ((local_bb4_var__u108 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond282_i173_stall_local;
wire [31:0] local_bb4_cond282_i173;

assign local_bb4_cond282_i173 = (local_bb4_or2804_i172 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond289_i175_stall_local;
wire [31:0] local_bb4_cond289_i175;

assign local_bb4_cond289_i175 = (local_bb4_or2875_i174 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext310_i187_stall_local;
wire [31:0] local_bb4_lnot_ext310_i187;

assign local_bb4_lnot_ext310_i187 = ((local_bb4_var__u109 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and293_i177_stall_local;
wire [31:0] local_bb4_and293_i177;

assign local_bb4_and293_i177 = ((local_bb4_cond282_i173 | 32'h80000000) & local_bb4_or275_i171);

// This section implements an unregistered operation.
// 
wire local_bb4_or294_i178_stall_local;
wire [31:0] local_bb4_or294_i178;

assign local_bb4_or294_i178 = ((local_bb4_cond289_i175 & 32'h7F800000) | (local_bb4_cond292_i176 & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i189_stall_local;
wire [31:0] local_bb4_reduction_0_i189;

assign local_bb4_reduction_0_i189 = ((local_bb4_lnot_ext310_i187 & 32'h1) & (local_bb4_lnot_ext_i186 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and302_i183_stall_local;
wire [31:0] local_bb4_and302_i183;

assign local_bb4_and302_i183 = ((local_bb4_conv300_i182 & 32'h1) & local_bb4_and293_i177);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i179_stall_local;
wire [31:0] local_bb4_or295_i179;

assign local_bb4_or295_i179 = ((local_bb4_or294_i178 & 32'h7FC00000) | local_bb4_and293_i177);

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i185_stall_local;
wire [31:0] local_bb4_lor_ext_i185;

assign local_bb4_lor_ext_i185 = ((local_bb4_cmp29649_i184 & 32'h1) | (local_bb4_and302_i183 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i190_stall_local;
wire [31:0] local_bb4_reduction_1_i190;

assign local_bb4_reduction_1_i190 = ((local_bb4_lnot_ext314_i188 & 32'h1) & (local_bb4_lor_ext_i185 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i191_stall_local;
wire [31:0] local_bb4_reduction_2_i191;

assign local_bb4_reduction_2_i191 = ((local_bb4_reduction_0_i189 & 32'h1) & (local_bb4_reduction_1_i190 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_add320_i192_stall_local;
wire [31:0] local_bb4_add320_i192;

assign local_bb4_add320_i192 = ((local_bb4_reduction_2_i191 & 32'h1) + local_bb4_or295_i179);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u110_stall_local;
wire [31:0] local_bb4_var__u110;

assign local_bb4_var__u110 = local_bb4_add320_i192;

// This section implements an unregistered operation.
// 
wire local_bb4__40_valid_out;
wire local_bb4__40_stall_in;
wire local_bb4__40_inputs_ready;
wire local_bb4__40_stall_local;
wire [31:0] local_bb4__40;

assign local_bb4__40_inputs_ready = (rnode_400to401_bb4_c1_ene7_0_valid_out_NO_SHIFT_REG & rnode_400to401_bb4_t_313_pop8_c1_ene4_0_valid_out_NO_SHIFT_REG & rnode_399to401_bb4_and269_i168_0_valid_out_NO_SHIFT_REG & rnode_400to401_bb4_resultSign_0_i151_0_valid_out_NO_SHIFT_REG & rnode_400to401_bb4_or2662_i164_0_valid_out_1_NO_SHIFT_REG & rnode_400to401_bb4__26_i49_0_valid_out_0_NO_SHIFT_REG & rnode_400to401_bb4__26_i49_0_valid_out_1_NO_SHIFT_REG & rnode_400to401_bb4__47_i161_0_valid_out_0_NO_SHIFT_REG & rnode_400to401_bb4_or2662_i164_0_valid_out_0_NO_SHIFT_REG & rnode_400to401_bb4__26_i49_0_valid_out_2_NO_SHIFT_REG & rnode_400to401_bb4_or2662_i164_0_valid_out_2_NO_SHIFT_REG & rnode_400to401_bb4_shr271_i166_0_valid_out_NO_SHIFT_REG & rnode_400to401_bb4__47_i161_0_valid_out_1_NO_SHIFT_REG & rnode_400to401_bb4_cmp296_i180_0_valid_out_NO_SHIFT_REG & rnode_400to401_bb4_cmp299_i181_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40 = (rnode_400to401_bb4_c1_ene7_0_NO_SHIFT_REG ? local_bb4_var__u110 : rnode_400to401_bb4_t_313_pop8_c1_ene4_0_NO_SHIFT_REG);
assign local_bb4__40_valid_out = 1'b1;
assign rnode_400to401_bb4_c1_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_t_313_pop8_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_399to401_bb4_and269_i168_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_resultSign_0_i151_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_or2662_i164_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__26_i49_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__26_i49_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__47_i161_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_or2662_i164_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__26_i49_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_or2662_i164_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_shr271_i166_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4__47_i161_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_cmp296_i180_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_400to401_bb4_cmp299_i181_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_401to402_bb4__40_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_401to402_bb4__40_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_401to402_bb4__40_0_NO_SHIFT_REG;
 logic rnode_401to402_bb4__40_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_401to402_bb4__40_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_401to402_bb4__40_1_NO_SHIFT_REG;
 logic rnode_401to402_bb4__40_0_reg_402_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_401to402_bb4__40_0_reg_402_NO_SHIFT_REG;
 logic rnode_401to402_bb4__40_0_valid_out_0_reg_402_NO_SHIFT_REG;
 logic rnode_401to402_bb4__40_0_stall_in_0_reg_402_NO_SHIFT_REG;
 logic rnode_401to402_bb4__40_0_stall_out_reg_402_NO_SHIFT_REG;

acl_data_fifo rnode_401to402_bb4__40_0_reg_402_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_401to402_bb4__40_0_reg_402_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_401to402_bb4__40_0_stall_in_0_reg_402_NO_SHIFT_REG),
	.valid_out(rnode_401to402_bb4__40_0_valid_out_0_reg_402_NO_SHIFT_REG),
	.stall_out(rnode_401to402_bb4__40_0_stall_out_reg_402_NO_SHIFT_REG),
	.data_in(local_bb4__40),
	.data_out(rnode_401to402_bb4__40_0_reg_402_NO_SHIFT_REG)
);

defparam rnode_401to402_bb4__40_0_reg_402_fifo.DEPTH = 1;
defparam rnode_401to402_bb4__40_0_reg_402_fifo.DATA_WIDTH = 32;
defparam rnode_401to402_bb4__40_0_reg_402_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_401to402_bb4__40_0_reg_402_fifo.IMPL = "shift_reg";

assign rnode_401to402_bb4__40_0_reg_402_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_stall_in = 1'b0;
assign rnode_401to402_bb4__40_0_stall_in_0_reg_402_NO_SHIFT_REG = 1'b0;
assign rnode_401to402_bb4__40_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_401to402_bb4__40_0_NO_SHIFT_REG = rnode_401to402_bb4__40_0_reg_402_NO_SHIFT_REG;
assign rnode_401to402_bb4__40_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_401to402_bb4__40_1_NO_SHIFT_REG = rnode_401to402_bb4__40_0_reg_402_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_t_313_push8__40_inputs_ready;
 reg local_bb4_t_313_push8__40_valid_out_NO_SHIFT_REG;
wire local_bb4_t_313_push8__40_stall_in;
wire local_bb4_t_313_push8__40_output_regs_ready;
wire [31:0] local_bb4_t_313_push8__40_result;
wire local_bb4_t_313_push8__40_fu_valid_out;
wire local_bb4_t_313_push8__40_fu_stall_out;
 reg [31:0] local_bb4_t_313_push8__40_NO_SHIFT_REG;
wire local_bb4_t_313_push8__40_causedstall;

acl_push local_bb4_t_313_push8__40_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_401to402_bb4_c1_ene8_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_401to402_bb4__40_0_NO_SHIFT_REG),
	.stall_out(local_bb4_t_313_push8__40_fu_stall_out),
	.valid_in(SFC_3_VALID_401_402_0_NO_SHIFT_REG),
	.valid_out(local_bb4_t_313_push8__40_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_t_313_push8__40_result),
	.feedback_out(feedback_data_out_8),
	.feedback_valid_out(feedback_valid_out_8),
	.feedback_stall_in(feedback_stall_in_8)
);

defparam local_bb4_t_313_push8__40_feedback.STALLFREE = 1;
defparam local_bb4_t_313_push8__40_feedback.DATA_WIDTH = 32;
defparam local_bb4_t_313_push8__40_feedback.FIFO_DEPTH = 9;
defparam local_bb4_t_313_push8__40_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_t_313_push8__40_feedback.STYLE = "REGULAR";

assign local_bb4_t_313_push8__40_inputs_ready = 1'b1;
assign local_bb4_t_313_push8__40_output_regs_ready = 1'b1;
assign SFC_3_VALID_401_402_0_stall_in_1 = 1'b0;
assign rnode_401to402_bb4__40_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_401to402_bb4_c1_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_t_313_push8__40_causedstall = (SFC_3_VALID_401_402_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_t_313_push8__40_NO_SHIFT_REG <= 'x;
		local_bb4_t_313_push8__40_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_t_313_push8__40_output_regs_ready)
		begin
			local_bb4_t_313_push8__40_NO_SHIFT_REG <= local_bb4_t_313_push8__40_result;
			local_bb4_t_313_push8__40_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_t_313_push8__40_stall_in))
			begin
				local_bb4_t_313_push8__40_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_402to403_bb4__40_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_402to403_bb4__40_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4__40_0_NO_SHIFT_REG;
 logic rnode_402to403_bb4__40_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_402to403_bb4__40_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4__40_1_NO_SHIFT_REG;
 logic rnode_402to403_bb4__40_0_reg_403_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_402to403_bb4__40_0_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4__40_0_valid_out_0_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4__40_0_stall_in_0_reg_403_NO_SHIFT_REG;
 logic rnode_402to403_bb4__40_0_stall_out_reg_403_NO_SHIFT_REG;

acl_data_fifo rnode_402to403_bb4__40_0_reg_403_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_402to403_bb4__40_0_reg_403_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_402to403_bb4__40_0_stall_in_0_reg_403_NO_SHIFT_REG),
	.valid_out(rnode_402to403_bb4__40_0_valid_out_0_reg_403_NO_SHIFT_REG),
	.stall_out(rnode_402to403_bb4__40_0_stall_out_reg_403_NO_SHIFT_REG),
	.data_in(rnode_401to402_bb4__40_1_NO_SHIFT_REG),
	.data_out(rnode_402to403_bb4__40_0_reg_403_NO_SHIFT_REG)
);

defparam rnode_402to403_bb4__40_0_reg_403_fifo.DEPTH = 1;
defparam rnode_402to403_bb4__40_0_reg_403_fifo.DATA_WIDTH = 32;
defparam rnode_402to403_bb4__40_0_reg_403_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_402to403_bb4__40_0_reg_403_fifo.IMPL = "shift_reg";

assign rnode_402to403_bb4__40_0_reg_403_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_401to402_bb4__40_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_402to403_bb4__40_0_stall_in_0_reg_403_NO_SHIFT_REG = 1'b0;
assign rnode_402to403_bb4__40_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_402to403_bb4__40_0_NO_SHIFT_REG = rnode_402to403_bb4__40_0_reg_403_NO_SHIFT_REG;
assign rnode_402to403_bb4__40_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_402to403_bb4__40_1_NO_SHIFT_REG = rnode_402to403_bb4__40_0_reg_403_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4___40_valid_out;
wire local_bb4___40_stall_in;
wire local_bb4___40_inputs_ready;
wire local_bb4___40_stall_local;
 reg [31:0] ffwd_12_0_reg_NO_SHIFT_REG;

assign local_bb4___40_inputs_ready = (SFC_3_VALID_402_403_0_valid_out_2_NO_SHIFT_REG & rnode_402to403_bb4__40_0_valid_out_0_NO_SHIFT_REG);
assign ffwd_12_0 = ffwd_12_0_reg_NO_SHIFT_REG;
assign local_bb4___40_valid_out = 1'b1;
assign SFC_3_VALID_402_403_0_stall_in_2 = 1'b0;
assign rnode_402to403_bb4__40_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock)
begin
	if ((1'b1 & SFC_3_VALID_402_403_0_NO_SHIFT_REG))
	begin
		ffwd_12_0_reg_NO_SHIFT_REG <= rnode_402to403_bb4__40_0_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_exi2_valid_out;
wire local_bb4_c1_exi2_stall_in;
wire local_bb4_c1_exi2_inputs_ready;
wire local_bb4_c1_exi2_stall_local;
wire [95:0] local_bb4_c1_exi2;

assign local_bb4_c1_exi2_inputs_ready = (rnode_402to403_bb4___0_valid_out_1_NO_SHIFT_REG & rnode_402to403_bb4__40_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_c1_exi2[63:0] = local_bb4_c1_exi1[63:0];
assign local_bb4_c1_exi2[95:64] = rnode_402to403_bb4__40_1_NO_SHIFT_REG;
assign local_bb4_c1_exi2_valid_out = 1'b1;
assign rnode_402to403_bb4___0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_402to403_bb4__40_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_c1_exit_c1_exi2_inputs_ready;
 reg local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG;
wire local_bb4_c1_exit_c1_exi2_stall_in;
 reg [95:0] local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG;
wire [95:0] local_bb4_c1_exit_c1_exi2_in;
wire local_bb4_c1_exit_c1_exi2_valid;
wire local_bb4_c1_exit_c1_exi2_causedstall;

acl_stall_free_sink local_bb4_c1_exit_c1_exi2_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb4_c1_exi2),
	.data_out(local_bb4_c1_exit_c1_exi2_in),
	.input_accepted(local_bb4_c1_enter_c1_eni8_input_accepted),
	.valid_out(local_bb4_c1_exit_c1_exi2_valid),
	.stall_in(~(local_bb4_c1_exit_c1_exi2_output_regs_ready)),
	.stall_entry(local_bb4_c1_exit_c1_exi2_entry_stall),
	.valid_in(local_bb4_c1_exit_c1_exi2_valid_in),
	.IIphases(local_bb4_c1_exit_c1_exi2_phases),
	.inc_pipelined_thread(local_bb4_c1_enter_c1_eni8_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb4_c1_enter_c1_eni8_dec_pipelined_thread)
);

defparam local_bb4_c1_exit_c1_exi2_instance.DATA_WIDTH = 96;
defparam local_bb4_c1_exit_c1_exi2_instance.PIPELINE_DEPTH = 69;
defparam local_bb4_c1_exit_c1_exi2_instance.SHARINGII = 1;
defparam local_bb4_c1_exit_c1_exi2_instance.SCHEDULEII = 9;
defparam local_bb4_c1_exit_c1_exi2_instance.ALWAYS_THROTTLE = 0;

assign local_bb4_c1_exit_c1_exi2_inputs_ready = 1'b1;
assign local_bb4_c1_exit_c1_exi2_output_regs_ready = (&(~(local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG) | ~(local_bb4_c1_exit_c1_exi2_stall_in)));
assign local_bb4_c1_exit_c1_exi2_valid_in = SFC_3_VALID_402_403_0_NO_SHIFT_REG;
assign local_bb4_c1_exi2_stall_in = 1'b0;
assign local_bb4_t_313_push8__40_stall_in = 1'b0;
assign local_bb4____stall_in = 1'b0;
assign local_bb4___40_stall_in = 1'b0;
assign SFC_3_VALID_402_403_0_stall_in_0 = 1'b0;
assign rnode_402to403_bb4_sum_312_push9___0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_c1_exit_c1_exi2_causedstall = (1'b1 && (1'b0 && !(~(local_bb4_c1_exit_c1_exi2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG <= 'x;
		local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c1_exit_c1_exi2_output_regs_ready)
		begin
			local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_in;
			local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_valid;
		end
		else
		begin
			if (~(local_bb4_c1_exit_c1_exi2_stall_in))
			begin
				local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [319:0] lvb_bb4_c0_exit214_c0_exi7_0_reg_NO_SHIFT_REG;
 reg lvb_bb4_c0_exe7_0_reg_NO_SHIFT_REG;
 reg [95:0] lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG & local_bb4_c0_exe7_valid_out & local_bb4_c0_exe4218_valid_out & rnode_407to408_bb4_c0_exit214_c0_exi7_0_valid_out_2_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb4_c1_exit_c1_exi2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe7_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe4218_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_407to408_bb4_c0_exit214_c0_exi7_0_stall_in_2_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb4_c0_exit214_c0_exi7_0 = lvb_bb4_c0_exit214_c0_exi7_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exit214_c0_exi7_1 = lvb_bb4_c0_exit214_c0_exi7_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe7_0 = lvb_bb4_c0_exe7_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe7_1 = lvb_bb4_c0_exe7_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exit_c1_exi2_0 = lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exit_c1_exi2_1 = lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_bb4_c0_exit214_c0_exi7_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe7_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb4_c0_exit214_c0_exi7_0_reg_NO_SHIFT_REG <= rnode_407to408_bb4_c0_exit214_c0_exi7_2_NO_SHIFT_REG;
			lvb_bb4_c0_exe7_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe7;
			lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG;
			branch_compare_result_NO_SHIFT_REG <= local_bb4_c0_exe4218;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_5
	(
		input 		clock,
		input 		resetn,
		input 		input_wii_cmp1017,
		input [31:0] 		input_wii_mul39,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u111,
		input 		valid_in,
		output 		stall_out,
		input [319:0] 		input_c0_exit214_c0_exi7,
		input 		input_c0_exe7,
		input [95:0] 		input_c1_exit_c1_exi2,
		output 		valid_out_0,
		input 		stall_in_0,
		output 		valid_out_1,
		input 		stall_in_1,
		input [31:0] 		workgroup_size,
		input 		start,
		output 		feedback_valid_out_5,
		input 		feedback_stall_in_5,
		output [31:0] 		feedback_data_out_5,
		output 		feedback_valid_out_6,
		input 		feedback_stall_in_6,
		output [31:0] 		feedback_data_out_6
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [319:0] input_c0_exit214_c0_exi7_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe7_staging_reg_NO_SHIFT_REG;
 reg [95:0] input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG;
 reg [319:0] local_lvm_c0_exit214_c0_exi7_NO_SHIFT_REG;
 reg local_lvm_c0_exe7_NO_SHIFT_REG;
 reg [95:0] local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_c0_exit214_c0_exi7_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe7_staging_reg_NO_SHIFT_REG <= 'x;
		input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_c0_exit214_c0_exi7_staging_reg_NO_SHIFT_REG <= input_c0_exit214_c0_exi7;
				input_c0_exe7_staging_reg_NO_SHIFT_REG <= input_c0_exe7;
				input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG <= input_c1_exit_c1_exi2;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_c0_exit214_c0_exi7_NO_SHIFT_REG <= input_c0_exit214_c0_exi7_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe7_NO_SHIFT_REG <= input_c0_exe7_staging_reg_NO_SHIFT_REG;
					local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG <= input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_c0_exit214_c0_exi7_NO_SHIFT_REG <= input_c0_exit214_c0_exi7;
					local_lvm_c0_exe7_NO_SHIFT_REG <= input_c0_exe7;
					local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG <= input_c1_exit_c1_exi2;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5_c1_exe2_valid_out;
wire local_bb5_c1_exe2_stall_in;
wire local_bb5_c1_exe2_inputs_ready;
wire local_bb5_c1_exe2_stall_local;
wire [31:0] local_bb5_c1_exe2;

assign local_bb5_c1_exe2_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb5_c1_exe2 = local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG[95:64];
assign local_bb5_c1_exe2_valid_out = local_bb5_c1_exe2_inputs_ready;
assign local_bb5_c1_exe2_stall_local = local_bb5_c1_exe2_stall_in;
assign merge_node_stall_in_0 = (|local_bb5_c1_exe2_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb5_c1_exe1_valid_out;
wire local_bb5_c1_exe1_stall_in;
wire local_bb5_c1_exe1_inputs_ready;
wire local_bb5_c1_exe1_stall_local;
wire [31:0] local_bb5_c1_exe1;

assign local_bb5_c1_exe1_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb5_c1_exe1 = local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG[63:32];
assign local_bb5_c1_exe1_valid_out = local_bb5_c1_exe1_inputs_ready;
assign local_bb5_c1_exe1_stall_local = local_bb5_c1_exe1_stall_in;
assign merge_node_stall_in_1 = (|local_bb5_c1_exe1_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb5_c0_exe6_valid_out;
wire local_bb5_c0_exe6_stall_in;
wire local_bb5_c0_exe6_inputs_ready;
wire local_bb5_c0_exe6_stall_local;
wire local_bb5_c0_exe6;

assign local_bb5_c0_exe6_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign local_bb5_c0_exe6 = local_lvm_c0_exit214_c0_exi7_NO_SHIFT_REG[272];
assign local_bb5_c0_exe6_valid_out = local_bb5_c0_exe6_inputs_ready;
assign local_bb5_c0_exe6_stall_local = local_bb5_c0_exe6_stall_in;
assign merge_node_stall_in_2 = (|local_bb5_c0_exe6_stall_local);

// This section implements a registered operation.
// 
wire local_bb5_t_219_push5_c1_exe2_inputs_ready;
 reg local_bb5_t_219_push5_c1_exe2_valid_out_NO_SHIFT_REG;
wire local_bb5_t_219_push5_c1_exe2_stall_in;
wire local_bb5_t_219_push5_c1_exe2_output_regs_ready;
wire [31:0] local_bb5_t_219_push5_c1_exe2_result;
wire local_bb5_t_219_push5_c1_exe2_fu_valid_out;
wire local_bb5_t_219_push5_c1_exe2_fu_stall_out;
 reg [31:0] local_bb5_t_219_push5_c1_exe2_NO_SHIFT_REG;
wire local_bb5_t_219_push5_c1_exe2_causedstall;

acl_push local_bb5_t_219_push5_c1_exe2_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_c0_exe7_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb5_c1_exe2),
	.stall_out(local_bb5_t_219_push5_c1_exe2_fu_stall_out),
	.valid_in(local_bb5_t_219_push5_c1_exe2_inputs_ready),
	.valid_out(local_bb5_t_219_push5_c1_exe2_fu_valid_out),
	.stall_in(~(local_bb5_t_219_push5_c1_exe2_output_regs_ready)),
	.data_out(local_bb5_t_219_push5_c1_exe2_result),
	.feedback_out(feedback_data_out_5),
	.feedback_valid_out(feedback_valid_out_5),
	.feedback_stall_in(feedback_stall_in_5)
);

defparam local_bb5_t_219_push5_c1_exe2_feedback.STALLFREE = 0;
defparam local_bb5_t_219_push5_c1_exe2_feedback.DATA_WIDTH = 32;
defparam local_bb5_t_219_push5_c1_exe2_feedback.FIFO_DEPTH = 3;
defparam local_bb5_t_219_push5_c1_exe2_feedback.MIN_FIFO_LATENCY = 3;
defparam local_bb5_t_219_push5_c1_exe2_feedback.STYLE = "REGULAR";

assign local_bb5_t_219_push5_c1_exe2_inputs_ready = (local_bb5_c1_exe2_valid_out & merge_node_valid_out_4_NO_SHIFT_REG);
assign local_bb5_t_219_push5_c1_exe2_output_regs_ready = (&(~(local_bb5_t_219_push5_c1_exe2_valid_out_NO_SHIFT_REG) | ~(local_bb5_t_219_push5_c1_exe2_stall_in)));
assign local_bb5_c1_exe2_stall_in = (local_bb5_t_219_push5_c1_exe2_fu_stall_out | ~(local_bb5_t_219_push5_c1_exe2_inputs_ready));
assign merge_node_stall_in_4 = (local_bb5_t_219_push5_c1_exe2_fu_stall_out | ~(local_bb5_t_219_push5_c1_exe2_inputs_ready));
assign local_bb5_t_219_push5_c1_exe2_causedstall = (local_bb5_t_219_push5_c1_exe2_inputs_ready && (local_bb5_t_219_push5_c1_exe2_fu_stall_out && !(~(local_bb5_t_219_push5_c1_exe2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_t_219_push5_c1_exe2_NO_SHIFT_REG <= 'x;
		local_bb5_t_219_push5_c1_exe2_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_t_219_push5_c1_exe2_output_regs_ready)
		begin
			local_bb5_t_219_push5_c1_exe2_NO_SHIFT_REG <= local_bb5_t_219_push5_c1_exe2_result;
			local_bb5_t_219_push5_c1_exe2_valid_out_NO_SHIFT_REG <= local_bb5_t_219_push5_c1_exe2_fu_valid_out;
		end
		else
		begin
			if (~(local_bb5_t_219_push5_c1_exe2_stall_in))
			begin
				local_bb5_t_219_push5_c1_exe2_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb5_sum_218_push6_c1_exe1_inputs_ready;
 reg local_bb5_sum_218_push6_c1_exe1_valid_out_NO_SHIFT_REG;
wire local_bb5_sum_218_push6_c1_exe1_stall_in;
wire local_bb5_sum_218_push6_c1_exe1_output_regs_ready;
wire [31:0] local_bb5_sum_218_push6_c1_exe1_result;
wire local_bb5_sum_218_push6_c1_exe1_fu_valid_out;
wire local_bb5_sum_218_push6_c1_exe1_fu_stall_out;
 reg [31:0] local_bb5_sum_218_push6_c1_exe1_NO_SHIFT_REG;
wire local_bb5_sum_218_push6_c1_exe1_causedstall;

acl_push local_bb5_sum_218_push6_c1_exe1_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_c0_exe7_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb5_c1_exe1),
	.stall_out(local_bb5_sum_218_push6_c1_exe1_fu_stall_out),
	.valid_in(local_bb5_sum_218_push6_c1_exe1_inputs_ready),
	.valid_out(local_bb5_sum_218_push6_c1_exe1_fu_valid_out),
	.stall_in(~(local_bb5_sum_218_push6_c1_exe1_output_regs_ready)),
	.data_out(local_bb5_sum_218_push6_c1_exe1_result),
	.feedback_out(feedback_data_out_6),
	.feedback_valid_out(feedback_valid_out_6),
	.feedback_stall_in(feedback_stall_in_6)
);

defparam local_bb5_sum_218_push6_c1_exe1_feedback.STALLFREE = 0;
defparam local_bb5_sum_218_push6_c1_exe1_feedback.DATA_WIDTH = 32;
defparam local_bb5_sum_218_push6_c1_exe1_feedback.FIFO_DEPTH = 3;
defparam local_bb5_sum_218_push6_c1_exe1_feedback.MIN_FIFO_LATENCY = 3;
defparam local_bb5_sum_218_push6_c1_exe1_feedback.STYLE = "REGULAR";

assign local_bb5_sum_218_push6_c1_exe1_inputs_ready = (local_bb5_c1_exe1_valid_out & merge_node_valid_out_3_NO_SHIFT_REG);
assign local_bb5_sum_218_push6_c1_exe1_output_regs_ready = (&(~(local_bb5_sum_218_push6_c1_exe1_valid_out_NO_SHIFT_REG) | ~(local_bb5_sum_218_push6_c1_exe1_stall_in)));
assign local_bb5_c1_exe1_stall_in = (local_bb5_sum_218_push6_c1_exe1_fu_stall_out | ~(local_bb5_sum_218_push6_c1_exe1_inputs_ready));
assign merge_node_stall_in_3 = (local_bb5_sum_218_push6_c1_exe1_fu_stall_out | ~(local_bb5_sum_218_push6_c1_exe1_inputs_ready));
assign local_bb5_sum_218_push6_c1_exe1_causedstall = (local_bb5_sum_218_push6_c1_exe1_inputs_ready && (local_bb5_sum_218_push6_c1_exe1_fu_stall_out && !(~(local_bb5_sum_218_push6_c1_exe1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_sum_218_push6_c1_exe1_NO_SHIFT_REG <= 'x;
		local_bb5_sum_218_push6_c1_exe1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_sum_218_push6_c1_exe1_output_regs_ready)
		begin
			local_bb5_sum_218_push6_c1_exe1_NO_SHIFT_REG <= local_bb5_sum_218_push6_c1_exe1_result;
			local_bb5_sum_218_push6_c1_exe1_valid_out_NO_SHIFT_REG <= local_bb5_sum_218_push6_c1_exe1_fu_valid_out;
		end
		else
		begin
			if (~(local_bb5_sum_218_push6_c1_exe1_stall_in))
			begin
				local_bb5_sum_218_push6_c1_exe1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb5_c0_exe6_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe6_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe6_0_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe6_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe6_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe6_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe6_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe6_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb5_c0_exe6_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb5_c0_exe6_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb5_c0_exe6_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb5_c0_exe6_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb5_c0_exe6_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb5_c0_exe6),
	.data_out(rnode_1to2_bb5_c0_exe6_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb5_c0_exe6_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb5_c0_exe6_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb5_c0_exe6_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb5_c0_exe6_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb5_c0_exe6_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb5_c0_exe6_valid_out;
assign local_bb5_c0_exe6_stall_in = rnode_1to2_bb5_c0_exe6_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb5_c0_exe6_0_NO_SHIFT_REG = rnode_1to2_bb5_c0_exe6_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb5_c0_exe6_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb5_c0_exe6_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb5_c0_exe6_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb5_c0_exe6_0_valid_out_reg_2_NO_SHIFT_REG;

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;

assign branch_var__inputs_ready = (local_bb5_t_219_push5_c1_exe2_valid_out_NO_SHIFT_REG & local_bb5_sum_218_push6_c1_exe1_valid_out_NO_SHIFT_REG & rnode_1to2_bb5_c0_exe6_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb5_t_219_push5_c1_exe2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb5_sum_218_push6_c1_exe1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to2_bb5_c0_exe6_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			branch_compare_result_NO_SHIFT_REG <= rnode_1to2_bb5_c0_exe6_0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_6
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_out,
		input 		input_wii_cmp1017,
		input [31:0] 		input_wii_mul39,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u112,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out_0,
		input 		stall_in_0,
		output [63:0] 		lvb_bb6_indvars_iv_next31_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [63:0] 		lvb_bb6_indvars_iv_next31_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		ffwd_10_0,
		input 		ffwd_6_0,
		input [31:0] 		ffwd_12_0,
		input [31:0] 		ffwd_11_0,
		input [63:0] 		ffwd_7_0,
		input [63:0] 		ffwd_4_0,
		input 		ffwd_9_0,
		output [63:0] 		ffwd_13_0,
		input [511:0] 		avm_local_bb6_st_c0_exe2225_readdata,
		input 		avm_local_bb6_st_c0_exe2225_readdatavalid,
		input 		avm_local_bb6_st_c0_exe2225_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe2225_address,
		output 		avm_local_bb6_st_c0_exe2225_read,
		output 		avm_local_bb6_st_c0_exe2225_write,
		input 		avm_local_bb6_st_c0_exe2225_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe2225_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe2225_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe2225_burstcount,
		output 		local_bb6_st_c0_exe2225_active,
		input 		clock2x
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb6_c0_enter219__inputs_ready;
 reg local_bb6_c0_enter219__valid_out_0_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_0;
 reg local_bb6_c0_enter219__valid_out_1_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_1;
 reg local_bb6_c0_enter219__valid_out_2_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_2;
 reg local_bb6_c0_enter219__valid_out_3_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_3;
 reg local_bb6_c0_enter219__valid_out_4_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_4;
 reg local_bb6_c0_enter219__valid_out_5_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_5;
 reg local_bb6_c0_enter219__valid_out_6_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_6;
 reg local_bb6_c0_enter219__valid_out_7_NO_SHIFT_REG;
wire local_bb6_c0_enter219__stall_in_7;
wire local_bb6_c0_enter219__output_regs_ready;
 reg [7:0] local_bb6_c0_enter219__NO_SHIFT_REG;
wire local_bb6_c0_enter219__input_accepted;
 reg local_bb6_c0_enter219__valid_bit_NO_SHIFT_REG;
wire local_bb6_c0_exit223_c0_exi3222_entry_stall;
wire local_bb6_c0_exit223_c0_exi3222_output_regs_ready;
wire [15:0] local_bb6_c0_exit223_c0_exi3222_valid_bits;
wire local_bb6_c0_exit223_c0_exi3222_valid_in;
wire local_bb6_c0_exit223_c0_exi3222_phases;
wire local_bb6_c0_enter219__inc_pipelined_thread;
wire local_bb6_c0_enter219__dec_pipelined_thread;
wire local_bb6_c0_enter219__causedstall;

assign local_bb6_c0_enter219__inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb6_c0_enter219__output_regs_ready = 1'b1;
assign local_bb6_c0_enter219__input_accepted = (local_bb6_c0_enter219__inputs_ready && !(local_bb6_c0_exit223_c0_exi3222_entry_stall));
assign local_bb6_c0_enter219__inc_pipelined_thread = 1'b1;
assign local_bb6_c0_enter219__dec_pipelined_thread = ~(1'b0);
assign merge_node_stall_in_0 = ((~(local_bb6_c0_enter219__inputs_ready) | local_bb6_c0_exit223_c0_exi3222_entry_stall) | ~(1'b1));
assign local_bb6_c0_enter219__causedstall = (1'b1 && ((~(local_bb6_c0_enter219__inputs_ready) | local_bb6_c0_exit223_c0_exi3222_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_enter219__valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb6_c0_enter219__valid_bit_NO_SHIFT_REG <= local_bb6_c0_enter219__input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_enter219__NO_SHIFT_REG <= 'x;
		local_bb6_c0_enter219__valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter219__valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter219__valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter219__valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter219__valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter219__valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter219__valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter219__valid_out_7_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_c0_enter219__output_regs_ready)
		begin
			local_bb6_c0_enter219__NO_SHIFT_REG <= 'x;
			local_bb6_c0_enter219__valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter219__valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter219__valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter219__valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter219__valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter219__valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter219__valid_out_6_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter219__valid_out_7_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb6_c0_enter219__stall_in_0))
			begin
				local_bb6_c0_enter219__valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter219__stall_in_1))
			begin
				local_bb6_c0_enter219__valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter219__stall_in_2))
			begin
				local_bb6_c0_enter219__valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter219__stall_in_3))
			begin
				local_bb6_c0_enter219__valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter219__stall_in_4))
			begin
				local_bb6_c0_enter219__valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter219__stall_in_5))
			begin
				local_bb6_c0_enter219__valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter219__stall_in_6))
			begin
				local_bb6_c0_enter219__valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter219__stall_in_7))
			begin
				local_bb6_c0_enter219__valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 18
//  * capacity = 18
 logic rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_valid_out_reg_19_NO_SHIFT_REG;
 logic rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_in_reg_19_NO_SHIFT_REG;
 logic rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_out_reg_19_NO_SHIFT_REG;

acl_data_fifo rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_in_reg_19_NO_SHIFT_REG),
	.valid_out(rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_valid_out_reg_19_NO_SHIFT_REG),
	.stall_out(rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_out_reg_19_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_fifo.DEPTH = 19;
defparam rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_fifo.DATA_WIDTH = 0;
defparam rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_fifo.IMPL = "ram";

assign rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_reg_19_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign merge_node_stall_in_1 = rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_out_reg_19_NO_SHIFT_REG;
assign rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_in_reg_19_NO_SHIFT_REG = rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_in_NO_SHIFT_REG;
assign rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_valid_out_NO_SHIFT_REG = rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_valid_out_reg_19_NO_SHIFT_REG;

// Register node:
//  * latency = 179
//  * capacity = 179
 logic rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_fifo.DEPTH = 180;
defparam rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_fifo.DATA_WIDTH = 0;
defparam rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_fifo.IMPL = "ram";

assign rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_180_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign merge_node_stall_in_2 = rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_out_reg_180_NO_SHIFT_REG;
assign rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_reg_180_NO_SHIFT_REG = rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_NO_SHIFT_REG;
assign rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_NO_SHIFT_REG = rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_10_stall_local;
wire local_bb6__acl_ffwd_dest_i1_10;

assign local_bb6__acl_ffwd_dest_i1_10 = ffwd_10_0;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_6_stall_local;
wire local_bb6__acl_ffwd_dest_i1_6;

assign local_bb6__acl_ffwd_dest_i1_6 = ffwd_6_0;

// This section implements an unregistered operation.
// 
wire local_bb6__40196_acl_ffwd_dest_f_12_stall_local;
wire [31:0] local_bb6__40196_acl_ffwd_dest_f_12;

assign local_bb6__40196_acl_ffwd_dest_f_12 = ffwd_12_0;

// This section implements an unregistered operation.
// 
wire local_bb6__195_acl_ffwd_dest_f_11_stall_local;
wire [31:0] local_bb6__195_acl_ffwd_dest_f_11;

assign local_bb6__195_acl_ffwd_dest_f_11 = ffwd_11_0;

// This section implements an unregistered operation.
// 
wire SFC_4_VALID_2_2_0_valid_out;
wire SFC_4_VALID_2_2_0_stall_in;
wire SFC_4_VALID_2_2_0_inputs_ready;
wire SFC_4_VALID_2_2_0_stall_local;
wire SFC_4_VALID_2_2_0;

assign SFC_4_VALID_2_2_0_inputs_ready = local_bb6_c0_enter219__valid_out_4_NO_SHIFT_REG;
assign SFC_4_VALID_2_2_0 = local_bb6_c0_enter219__valid_bit_NO_SHIFT_REG;
assign SFC_4_VALID_2_2_0_valid_out = 1'b1;
assign local_bb6_c0_enter219__stall_in_4 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_c0_enter219__stall_in_5 = 1'b0;
assign rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_c0_enter219__stall_in_6 = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_c0_enter219__stall_in_7 = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_valid_out_NO_SHIFT_REG;
 logic rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_in_NO_SHIFT_REG;
 logic rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_inputs_ready_NO_SHIFT_REG;
 logic rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_valid_out_reg_20_NO_SHIFT_REG;
 logic rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_in_reg_20_NO_SHIFT_REG;
 logic rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_out_reg_20_NO_SHIFT_REG;

acl_data_fifo rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_in_reg_20_NO_SHIFT_REG),
	.valid_out(rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_valid_out_reg_20_NO_SHIFT_REG),
	.stall_out(rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_out_reg_20_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_fifo.DEPTH = 1;
defparam rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_fifo.DATA_WIDTH = 0;
defparam rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_fifo.IMPL = "ll_reg";

assign rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_reg_20_inputs_ready_NO_SHIFT_REG = rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_valid_out_NO_SHIFT_REG;
assign rnode_1to19_bb6__acl_ffwd_dest_i64_7_0_stall_in_NO_SHIFT_REG = rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_out_reg_20_NO_SHIFT_REG;
assign rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_in_reg_20_NO_SHIFT_REG = rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_in_NO_SHIFT_REG;
assign rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_valid_out_NO_SHIFT_REG = rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_valid_out_reg_20_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_fifo.DATA_WIDTH = 0;
defparam rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_fifo.IMPL = "ll_reg";

assign rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_reg_181_inputs_ready_NO_SHIFT_REG = rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_NO_SHIFT_REG;
assign rnode_1to180_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_NO_SHIFT_REG = rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_out_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_reg_181_NO_SHIFT_REG = rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_NO_SHIFT_REG;
assign rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_NO_SHIFT_REG = rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_reg_181_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end48_loopexit_select92_stall_local;
wire local_bb6_do_directly_for_end48_loopexit_select92;

assign local_bb6_do_directly_for_end48_loopexit_select92 = (local_bb6__acl_ffwd_dest_i1_10 ^ 1'b1);

// This section implements a registered operation.
// 
wire SFC_4_VALID_2_3_0_inputs_ready;
 reg SFC_4_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_2_3_0_stall_in;
wire SFC_4_VALID_2_3_0_output_regs_ready;
 reg SFC_4_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_2_3_0_causedstall;

assign SFC_4_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_4_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_2_2_0_stall_in = 1'b0;
assign SFC_4_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_2_3_0_output_regs_ready)
		begin
			SFC_4_VALID_2_3_0_NO_SHIFT_REG <= SFC_4_VALID_2_2_0;
		end
	end
end


// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i64_7_stall_local;
wire [63:0] local_bb6__acl_ffwd_dest_i64_7;

assign local_bb6__acl_ffwd_dest_i64_7 = ffwd_7_0;

// This section implements an unregistered operation.
// 
wire local_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_stall_local;
wire [63:0] local_bb6_indvars_iv30193_acl_ffwd_dest_i64_4;

assign local_bb6_indvars_iv30193_acl_ffwd_dest_i64_4 = ffwd_4_0;

// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end48_loopexit_select_stall_local;
wire local_bb6_do_directly_for_end48_loopexit_select;

assign local_bb6_do_directly_for_end48_loopexit_select = (local_bb6__acl_ffwd_dest_i1_6 & local_bb6_do_directly_for_end48_loopexit_select92);

// This section implements a registered operation.
// 
wire SFC_4_VALID_3_4_0_inputs_ready;
 reg SFC_4_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_3_4_0_stall_in;
wire SFC_4_VALID_3_4_0_output_regs_ready;
 reg SFC_4_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_3_4_0_causedstall;

assign SFC_4_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_4_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_2_3_0_stall_in = 1'b0;
assign SFC_4_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_3_4_0_output_regs_ready)
		begin
			SFC_4_VALID_3_4_0_NO_SHIFT_REG <= SFC_4_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb6_arrayidx53_valid_out;
wire local_bb6_arrayidx53_stall_in;
wire local_bb6_arrayidx53_inputs_ready;
wire local_bb6_arrayidx53_stall_local;
wire [63:0] local_bb6_arrayidx53;

assign local_bb6_arrayidx53_inputs_ready = rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_valid_out_NO_SHIFT_REG;
assign local_bb6_arrayidx53 = ((input_out & 64'hFFFFFFFFFFFFFC00) + (local_bb6__acl_ffwd_dest_i64_7 << 6'h2));
assign local_bb6_arrayidx53_valid_out = local_bb6_arrayidx53_inputs_ready;
assign local_bb6_arrayidx53_stall_local = local_bb6_arrayidx53_stall_in;
assign rnode_19to20_bb6__acl_ffwd_dest_i64_7_0_stall_in_NO_SHIFT_REG = (|local_bb6_arrayidx53_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_indvars_iv_next31_valid_out;
wire local_bb6_indvars_iv_next31_stall_in;
wire local_bb6_indvars_iv_next31_inputs_ready;
wire local_bb6_indvars_iv_next31_stall_local;
wire [63:0] local_bb6_indvars_iv_next31;

assign local_bb6_indvars_iv_next31_inputs_ready = rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_valid_out_NO_SHIFT_REG;
assign local_bb6_indvars_iv_next31 = (local_bb6_indvars_iv30193_acl_ffwd_dest_i64_4 + 64'h1);
assign local_bb6_indvars_iv_next31_valid_out = local_bb6_indvars_iv_next31_inputs_ready;
assign local_bb6_indvars_iv_next31_stall_local = local_bb6_indvars_iv_next31_stall_in;
assign rnode_180to181_bb6_indvars_iv30193_acl_ffwd_dest_i64_4_0_stall_in_NO_SHIFT_REG = (|local_bb6_indvars_iv_next31_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_select73_stall_local;
wire [31:0] local_bb6_select73;

assign local_bb6_select73 = (local_bb6_do_directly_for_end48_loopexit_select ? local_bb6__40196_acl_ffwd_dest_f_12 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end48_loopexit_select_valid_out_2;
wire local_bb6_do_directly_for_end48_loopexit_select_stall_in_2;
wire local_bb6_select73_valid_out;
wire local_bb6_select73_stall_in;
wire local_bb6_select76_valid_out;
wire local_bb6_select76_stall_in;
wire local_bb6_select76_inputs_ready;
wire local_bb6_select76_stall_local;
wire [31:0] local_bb6_select76;

assign local_bb6_select76_inputs_ready = (local_bb6_c0_enter219__valid_out_0_NO_SHIFT_REG & local_bb6_c0_enter219__valid_out_1_NO_SHIFT_REG & local_bb6_c0_enter219__valid_out_2_NO_SHIFT_REG & local_bb6_c0_enter219__valid_out_3_NO_SHIFT_REG);
assign local_bb6_select76 = (local_bb6_do_directly_for_end48_loopexit_select ? local_bb6__195_acl_ffwd_dest_f_11 : 32'h0);
assign local_bb6_do_directly_for_end48_loopexit_select_valid_out_2 = 1'b1;
assign local_bb6_select73_valid_out = 1'b1;
assign local_bb6_select76_valid_out = 1'b1;
assign local_bb6_c0_enter219__stall_in_0 = 1'b0;
assign local_bb6_c0_enter219__stall_in_1 = 1'b0;
assign local_bb6_c0_enter219__stall_in_2 = 1'b0;
assign local_bb6_c0_enter219__stall_in_3 = 1'b0;

// This section implements a registered operation.
// 
wire SFC_4_VALID_4_5_0_inputs_ready;
 reg SFC_4_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_4_5_0_stall_in;
wire SFC_4_VALID_4_5_0_output_regs_ready;
 reg SFC_4_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_4_5_0_causedstall;

assign SFC_4_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_4_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_3_4_0_stall_in = 1'b0;
assign SFC_4_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_4_5_0_output_regs_ready)
		begin
			SFC_4_VALID_4_5_0_NO_SHIFT_REG <= SFC_4_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_cmp4194_acl_ffwd_dest_i1_9_stall_local;
wire local_bb6_cmp4194_acl_ffwd_dest_i1_9;

assign local_bb6_cmp4194_acl_ffwd_dest_i1_9 = ffwd_9_0;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_6_u113_stall_local;
wire local_bb6__acl_ffwd_dest_i1_6_u113;

assign local_bb6__acl_ffwd_dest_i1_6_u113 = ffwd_6_0;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_10_u114_stall_local;
wire local_bb6__acl_ffwd_dest_i1_10_u114;

assign local_bb6__acl_ffwd_dest_i1_10_u114 = ffwd_10_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_20to21_bb6_arrayidx53_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx53_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx53_0_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx53_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx53_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx53_1_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx53_0_reg_21_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx53_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx53_0_valid_out_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx53_0_stall_in_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx53_0_stall_out_reg_21_NO_SHIFT_REG;
 reg rnode_20to21_bb6_arrayidx53_0_consumed_0_NO_SHIFT_REG;
 reg rnode_20to21_bb6_arrayidx53_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_20to21_bb6_arrayidx53_0_reg_21_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_20to21_bb6_arrayidx53_0_reg_21_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_20to21_bb6_arrayidx53_0_stall_in_0_reg_21_NO_SHIFT_REG),
	.valid_out(rnode_20to21_bb6_arrayidx53_0_valid_out_0_reg_21_NO_SHIFT_REG),
	.stall_out(rnode_20to21_bb6_arrayidx53_0_stall_out_reg_21_NO_SHIFT_REG),
	.data_in((local_bb6_arrayidx53 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_20to21_bb6_arrayidx53_0_reg_21_NO_SHIFT_REG)
);

defparam rnode_20to21_bb6_arrayidx53_0_reg_21_fifo.DEPTH = 2;
defparam rnode_20to21_bb6_arrayidx53_0_reg_21_fifo.DATA_WIDTH = 64;
defparam rnode_20to21_bb6_arrayidx53_0_reg_21_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_20to21_bb6_arrayidx53_0_reg_21_fifo.IMPL = "ll_reg";

assign rnode_20to21_bb6_arrayidx53_0_reg_21_inputs_ready_NO_SHIFT_REG = local_bb6_arrayidx53_valid_out;
assign local_bb6_arrayidx53_stall_in = rnode_20to21_bb6_arrayidx53_0_stall_out_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb6_arrayidx53_0_stall_in_0_reg_21_NO_SHIFT_REG = ((rnode_20to21_bb6_arrayidx53_0_stall_in_0_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx53_0_consumed_0_NO_SHIFT_REG)) | (rnode_20to21_bb6_arrayidx53_0_stall_in_1_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx53_0_consumed_1_NO_SHIFT_REG)));
assign rnode_20to21_bb6_arrayidx53_0_valid_out_0_NO_SHIFT_REG = (rnode_20to21_bb6_arrayidx53_0_valid_out_0_reg_21_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx53_0_consumed_0_NO_SHIFT_REG));
assign rnode_20to21_bb6_arrayidx53_0_valid_out_1_NO_SHIFT_REG = (rnode_20to21_bb6_arrayidx53_0_valid_out_0_reg_21_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx53_0_consumed_1_NO_SHIFT_REG));
assign rnode_20to21_bb6_arrayidx53_0_NO_SHIFT_REG = rnode_20to21_bb6_arrayidx53_0_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb6_arrayidx53_1_NO_SHIFT_REG = rnode_20to21_bb6_arrayidx53_0_reg_21_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_20to21_bb6_arrayidx53_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_20to21_bb6_arrayidx53_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_20to21_bb6_arrayidx53_0_consumed_0_NO_SHIFT_REG <= (rnode_20to21_bb6_arrayidx53_0_valid_out_0_reg_21_NO_SHIFT_REG & (rnode_20to21_bb6_arrayidx53_0_consumed_0_NO_SHIFT_REG | ~(rnode_20to21_bb6_arrayidx53_0_stall_in_0_NO_SHIFT_REG)) & rnode_20to21_bb6_arrayidx53_0_stall_in_0_reg_21_NO_SHIFT_REG);
		rnode_20to21_bb6_arrayidx53_0_consumed_1_NO_SHIFT_REG <= (rnode_20to21_bb6_arrayidx53_0_valid_out_0_reg_21_NO_SHIFT_REG & (rnode_20to21_bb6_arrayidx53_0_consumed_1_NO_SHIFT_REG | ~(rnode_20to21_bb6_arrayidx53_0_stall_in_1_NO_SHIFT_REG)) & rnode_20to21_bb6_arrayidx53_0_stall_in_0_reg_21_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb6_do_directly_for_end48_loopexit_select),
	.data_out(rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_do_directly_for_end48_loopexit_select_stall_in_2 = 1'b0;
assign rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG = rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb6_div49_inputs_ready;
 reg local_bb6_div49_valid_out_NO_SHIFT_REG;
wire local_bb6_div49_stall_in;
wire local_bb6_div49_output_regs_ready;
wire [31:0] local_bb6_div49;
 reg local_bb6_div49_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb6_div49_valid_pipe_12_NO_SHIFT_REG;
wire local_bb6_div49_causedstall;

acl_fp_div_s5 fp_module_local_bb6_div49 (
	.clock(clock),
	.dataa(local_bb6_select73),
	.datab(local_bb6_select76),
	.enable(local_bb6_div49_output_regs_ready),
	.result(local_bb6_div49)
);


assign local_bb6_div49_inputs_ready = 1'b1;
assign local_bb6_div49_output_regs_ready = 1'b1;
assign local_bb6_select73_stall_in = 1'b0;
assign local_bb6_select76_stall_in = 1'b0;
assign local_bb6_div49_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_div49_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb6_div49_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_div49_output_regs_ready)
		begin
			local_bb6_div49_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb6_div49_valid_pipe_1_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_0_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_2_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_1_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_3_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_2_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_4_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_3_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_5_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_4_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_6_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_5_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_7_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_6_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_8_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_7_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_9_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_8_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_10_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_9_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_11_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_10_NO_SHIFT_REG;
			local_bb6_div49_valid_pipe_12_NO_SHIFT_REG <= local_bb6_div49_valid_pipe_11_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_div49_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_div49_output_regs_ready)
		begin
			local_bb6_div49_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb6_div49_stall_in))
			begin
				local_bb6_div49_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_5_6_0_inputs_ready;
 reg SFC_4_VALID_5_6_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_5_6_0_stall_in;
wire SFC_4_VALID_5_6_0_output_regs_ready;
 reg SFC_4_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_5_6_0_causedstall;

assign SFC_4_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_4_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_4_5_0_stall_in = 1'b0;
assign SFC_4_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_5_6_0_output_regs_ready)
		begin
			SFC_4_VALID_5_6_0_NO_SHIFT_REG <= SFC_4_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_cmp4_not_stall_local;
wire local_bb6_cmp4_not;

assign local_bb6_cmp4_not = (local_bb6_cmp4194_acl_ffwd_dest_i1_9 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb6__arrayidx53_valid_out;
wire local_bb6__arrayidx53_stall_in;
wire local_bb6__arrayidx53_inputs_ready;
wire local_bb6__arrayidx53_stall_local;
 reg [63:0] ffwd_13_0_reg_NO_SHIFT_REG;

assign local_bb6__arrayidx53_inputs_ready = rnode_20to21_bb6_arrayidx53_0_valid_out_1_NO_SHIFT_REG;
assign ffwd_13_0 = ffwd_13_0_reg_NO_SHIFT_REG;
assign local_bb6__arrayidx53_valid_out = local_bb6__arrayidx53_inputs_ready;
assign local_bb6__arrayidx53_stall_local = local_bb6__arrayidx53_stall_in;
assign rnode_20to21_bb6_arrayidx53_0_stall_in_1_NO_SHIFT_REG = (|local_bb6__arrayidx53_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb6__arrayidx53_inputs_ready))
	begin
		ffwd_13_0_reg_NO_SHIFT_REG <= (rnode_20to21_bb6_arrayidx53_1_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
	end
end


// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG),
	.data_out(rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_NO_SHIFT_REG)
);

defparam rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_fifo.DATA_WIDTH = 1;
defparam rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6_do_directly_for_end48_loopexit_select_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG = rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_reg_15_NO_SHIFT_REG;
assign rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_4_VALID_6_7_0_inputs_ready;
 reg SFC_4_VALID_6_7_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_6_7_0_stall_in;
wire SFC_4_VALID_6_7_0_output_regs_ready;
 reg SFC_4_VALID_6_7_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_6_7_0_causedstall;

assign SFC_4_VALID_6_7_0_inputs_ready = 1'b1;
assign SFC_4_VALID_6_7_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_5_6_0_stall_in = 1'b0;
assign SFC_4_VALID_6_7_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_6_7_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_6_7_0_output_regs_ready)
		begin
			SFC_4_VALID_6_7_0_NO_SHIFT_REG <= SFC_4_VALID_5_6_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_not__phi_decision86_select_stall_local;
wire local_bb6_not__phi_decision86_select;

assign local_bb6_not__phi_decision86_select = (local_bb6__acl_ffwd_dest_i1_6_u113 & local_bb6_cmp4_not);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG),
	.data_out(rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_NO_SHIFT_REG)
);

defparam rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_fifo.DATA_WIDTH = 1;
defparam rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6_do_directly_for_end48_loopexit_select_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG = rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_reg_16_NO_SHIFT_REG;
assign rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_4_VALID_7_8_0_inputs_ready;
 reg SFC_4_VALID_7_8_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_7_8_0_stall_in;
wire SFC_4_VALID_7_8_0_output_regs_ready;
 reg SFC_4_VALID_7_8_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_7_8_0_causedstall;

assign SFC_4_VALID_7_8_0_inputs_ready = 1'b1;
assign SFC_4_VALID_7_8_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_6_7_0_stall_in = 1'b0;
assign SFC_4_VALID_7_8_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_7_8_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_7_8_0_output_regs_ready)
		begin
			SFC_4_VALID_7_8_0_NO_SHIFT_REG <= SFC_4_VALID_6_7_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end48_select_stall_local;
wire local_bb6_do_directly_for_end48_select;

assign local_bb6_do_directly_for_end48_select = (local_bb6__acl_ffwd_dest_i1_10_u114 & local_bb6_not__phi_decision86_select);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exi1220_stall_local;
wire [95:0] local_bb6_c0_exi1220;

assign local_bb6_c0_exi1220[7:0] = 8'bx;
assign local_bb6_c0_exi1220[8] = local_bb6_not__phi_decision86_select;
assign local_bb6_c0_exi1220[95:9] = 87'bx;

// This section implements a registered operation.
// 
wire SFC_4_VALID_8_9_0_inputs_ready;
 reg SFC_4_VALID_8_9_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_8_9_0_stall_in;
wire SFC_4_VALID_8_9_0_output_regs_ready;
 reg SFC_4_VALID_8_9_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_8_9_0_causedstall;

assign SFC_4_VALID_8_9_0_inputs_ready = 1'b1;
assign SFC_4_VALID_8_9_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_7_8_0_stall_in = 1'b0;
assign SFC_4_VALID_8_9_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_8_9_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_8_9_0_output_regs_ready)
		begin
			SFC_4_VALID_8_9_0_NO_SHIFT_REG <= SFC_4_VALID_7_8_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_or_stall_local;
wire local_bb6_or;

assign local_bb6_or = (local_bb6_do_directly_for_end48_select | rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exi2221_stall_local;
wire [95:0] local_bb6_c0_exi2221;

assign local_bb6_c0_exi2221[31:0] = local_bb6_c0_exi1220[31:0];
assign local_bb6_c0_exi2221[63:32] = local_bb6_div49;
assign local_bb6_c0_exi2221[95:64] = local_bb6_c0_exi1220[95:64];

// This section implements a registered operation.
// 
wire SFC_4_VALID_9_10_0_inputs_ready;
 reg SFC_4_VALID_9_10_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_9_10_0_stall_in;
wire SFC_4_VALID_9_10_0_output_regs_ready;
 reg SFC_4_VALID_9_10_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_9_10_0_causedstall;

assign SFC_4_VALID_9_10_0_inputs_ready = 1'b1;
assign SFC_4_VALID_9_10_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_8_9_0_stall_in = 1'b0;
assign SFC_4_VALID_9_10_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_9_10_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_9_10_0_output_regs_ready)
		begin
			SFC_4_VALID_9_10_0_NO_SHIFT_REG <= SFC_4_VALID_8_9_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_cmp_phi_decision80_xor_or_stall_local;
wire local_bb6_cmp_phi_decision80_xor_or;

assign local_bb6_cmp_phi_decision80_xor_or = (local_bb6_or ^ 1'b1);

// This section implements a registered operation.
// 
wire SFC_4_VALID_10_11_0_inputs_ready;
 reg SFC_4_VALID_10_11_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_10_11_0_stall_in;
wire SFC_4_VALID_10_11_0_output_regs_ready;
 reg SFC_4_VALID_10_11_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_10_11_0_causedstall;

assign SFC_4_VALID_10_11_0_inputs_ready = 1'b1;
assign SFC_4_VALID_10_11_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_9_10_0_stall_in = 1'b0;
assign SFC_4_VALID_10_11_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_10_11_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_10_11_0_output_regs_ready)
		begin
			SFC_4_VALID_10_11_0_NO_SHIFT_REG <= SFC_4_VALID_9_10_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_c0_exi3222_valid_out;
wire local_bb6_c0_exi3222_stall_in;
wire local_bb6_c0_exi3222_inputs_ready;
wire local_bb6_c0_exi3222_stall_local;
wire [95:0] local_bb6_c0_exi3222;

assign local_bb6_c0_exi3222_inputs_ready = (local_bb6_div49_valid_out_NO_SHIFT_REG & rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG & rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_valid_out_NO_SHIFT_REG & rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_valid_out_NO_SHIFT_REG & rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_valid_out_NO_SHIFT_REG);
assign local_bb6_c0_exi3222[63:0] = local_bb6_c0_exi2221[63:0];
assign local_bb6_c0_exi3222[64] = local_bb6_cmp_phi_decision80_xor_or;
assign local_bb6_c0_exi3222[95:65] = local_bb6_c0_exi2221[95:65];
assign local_bb6_c0_exi3222_valid_out = 1'b1;
assign local_bb6_div49_stall_in = 1'b0;
assign rnode_15to16_bb6_cmp4194_acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_6_u113_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_10_u114_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_do_directly_for_end48_loopexit_select_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_4_VALID_11_12_0_inputs_ready;
 reg SFC_4_VALID_11_12_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_11_12_0_stall_in;
wire SFC_4_VALID_11_12_0_output_regs_ready;
 reg SFC_4_VALID_11_12_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_11_12_0_causedstall;

assign SFC_4_VALID_11_12_0_inputs_ready = 1'b1;
assign SFC_4_VALID_11_12_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_10_11_0_stall_in = 1'b0;
assign SFC_4_VALID_11_12_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_11_12_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_11_12_0_output_regs_ready)
		begin
			SFC_4_VALID_11_12_0_NO_SHIFT_REG <= SFC_4_VALID_10_11_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_12_13_0_inputs_ready;
 reg SFC_4_VALID_12_13_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_12_13_0_stall_in;
wire SFC_4_VALID_12_13_0_output_regs_ready;
 reg SFC_4_VALID_12_13_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_12_13_0_causedstall;

assign SFC_4_VALID_12_13_0_inputs_ready = 1'b1;
assign SFC_4_VALID_12_13_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_11_12_0_stall_in = 1'b0;
assign SFC_4_VALID_12_13_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_12_13_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_12_13_0_output_regs_ready)
		begin
			SFC_4_VALID_12_13_0_NO_SHIFT_REG <= SFC_4_VALID_11_12_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_13_14_0_inputs_ready;
 reg SFC_4_VALID_13_14_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_13_14_0_stall_in;
wire SFC_4_VALID_13_14_0_output_regs_ready;
 reg SFC_4_VALID_13_14_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_13_14_0_causedstall;

assign SFC_4_VALID_13_14_0_inputs_ready = 1'b1;
assign SFC_4_VALID_13_14_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_12_13_0_stall_in = 1'b0;
assign SFC_4_VALID_13_14_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_13_14_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_13_14_0_output_regs_ready)
		begin
			SFC_4_VALID_13_14_0_NO_SHIFT_REG <= SFC_4_VALID_12_13_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_14_15_0_inputs_ready;
 reg SFC_4_VALID_14_15_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_14_15_0_stall_in;
wire SFC_4_VALID_14_15_0_output_regs_ready;
 reg SFC_4_VALID_14_15_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_14_15_0_causedstall;

assign SFC_4_VALID_14_15_0_inputs_ready = 1'b1;
assign SFC_4_VALID_14_15_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_13_14_0_stall_in = 1'b0;
assign SFC_4_VALID_14_15_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_14_15_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_14_15_0_output_regs_ready)
		begin
			SFC_4_VALID_14_15_0_NO_SHIFT_REG <= SFC_4_VALID_13_14_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_15_16_0_inputs_ready;
 reg SFC_4_VALID_15_16_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_15_16_0_stall_in;
wire SFC_4_VALID_15_16_0_output_regs_ready;
 reg SFC_4_VALID_15_16_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_15_16_0_causedstall;

assign SFC_4_VALID_15_16_0_inputs_ready = 1'b1;
assign SFC_4_VALID_15_16_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_14_15_0_stall_in = 1'b0;
assign SFC_4_VALID_15_16_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_15_16_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_15_16_0_output_regs_ready)
		begin
			SFC_4_VALID_15_16_0_NO_SHIFT_REG <= SFC_4_VALID_14_15_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb6_c0_exit223_c0_exi3222_inputs_ready;
 reg local_bb6_c0_exit223_c0_exi3222_valid_out_0_NO_SHIFT_REG;
wire local_bb6_c0_exit223_c0_exi3222_stall_in_0;
 reg local_bb6_c0_exit223_c0_exi3222_valid_out_1_NO_SHIFT_REG;
wire local_bb6_c0_exit223_c0_exi3222_stall_in_1;
 reg local_bb6_c0_exit223_c0_exi3222_valid_out_2_NO_SHIFT_REG;
wire local_bb6_c0_exit223_c0_exi3222_stall_in_2;
 reg [95:0] local_bb6_c0_exit223_c0_exi3222_NO_SHIFT_REG;
wire [95:0] local_bb6_c0_exit223_c0_exi3222_in;
wire local_bb6_c0_exit223_c0_exi3222_valid;
wire local_bb6_c0_exit223_c0_exi3222_causedstall;

acl_stall_free_sink local_bb6_c0_exit223_c0_exi3222_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb6_c0_exi3222),
	.data_out(local_bb6_c0_exit223_c0_exi3222_in),
	.input_accepted(local_bb6_c0_enter219__input_accepted),
	.valid_out(local_bb6_c0_exit223_c0_exi3222_valid),
	.stall_in(~(local_bb6_c0_exit223_c0_exi3222_output_regs_ready)),
	.stall_entry(local_bb6_c0_exit223_c0_exi3222_entry_stall),
	.valid_in(local_bb6_c0_exit223_c0_exi3222_valid_in),
	.IIphases(local_bb6_c0_exit223_c0_exi3222_phases),
	.inc_pipelined_thread(local_bb6_c0_enter219__inc_pipelined_thread),
	.dec_pipelined_thread(local_bb6_c0_enter219__dec_pipelined_thread)
);

defparam local_bb6_c0_exit223_c0_exi3222_instance.DATA_WIDTH = 96;
defparam local_bb6_c0_exit223_c0_exi3222_instance.PIPELINE_DEPTH = 20;
defparam local_bb6_c0_exit223_c0_exi3222_instance.SHARINGII = 1;
defparam local_bb6_c0_exit223_c0_exi3222_instance.SCHEDULEII = 1;
defparam local_bb6_c0_exit223_c0_exi3222_instance.ALWAYS_THROTTLE = 0;

assign local_bb6_c0_exit223_c0_exi3222_inputs_ready = 1'b1;
assign local_bb6_c0_exit223_c0_exi3222_output_regs_ready = ((~(local_bb6_c0_exit223_c0_exi3222_valid_out_0_NO_SHIFT_REG) | ~(local_bb6_c0_exit223_c0_exi3222_stall_in_0)) & (~(local_bb6_c0_exit223_c0_exi3222_valid_out_1_NO_SHIFT_REG) | ~(local_bb6_c0_exit223_c0_exi3222_stall_in_1)) & (~(local_bb6_c0_exit223_c0_exi3222_valid_out_2_NO_SHIFT_REG) | ~(local_bb6_c0_exit223_c0_exi3222_stall_in_2)));
assign local_bb6_c0_exit223_c0_exi3222_valid_in = SFC_4_VALID_15_16_0_NO_SHIFT_REG;
assign local_bb6_c0_exi3222_stall_in = 1'b0;
assign SFC_4_VALID_15_16_0_stall_in = 1'b0;
assign local_bb6_c0_exit223_c0_exi3222_causedstall = (1'b1 && (1'b0 && !(~(local_bb6_c0_exit223_c0_exi3222_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_exit223_c0_exi3222_NO_SHIFT_REG <= 'x;
		local_bb6_c0_exit223_c0_exi3222_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_exit223_c0_exi3222_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_exit223_c0_exi3222_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_c0_exit223_c0_exi3222_output_regs_ready)
		begin
			local_bb6_c0_exit223_c0_exi3222_NO_SHIFT_REG <= local_bb6_c0_exit223_c0_exi3222_in;
			local_bb6_c0_exit223_c0_exi3222_valid_out_0_NO_SHIFT_REG <= local_bb6_c0_exit223_c0_exi3222_valid;
			local_bb6_c0_exit223_c0_exi3222_valid_out_1_NO_SHIFT_REG <= local_bb6_c0_exit223_c0_exi3222_valid;
			local_bb6_c0_exit223_c0_exi3222_valid_out_2_NO_SHIFT_REG <= local_bb6_c0_exit223_c0_exi3222_valid;
		end
		else
		begin
			if (~(local_bb6_c0_exit223_c0_exi3222_stall_in_0))
			begin
				local_bb6_c0_exit223_c0_exi3222_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_exit223_c0_exi3222_stall_in_1))
			begin
				local_bb6_c0_exit223_c0_exi3222_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_exit223_c0_exi3222_stall_in_2))
			begin
				local_bb6_c0_exit223_c0_exi3222_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_c0_exe1224_valid_out;
wire local_bb6_c0_exe1224_stall_in;
wire local_bb6_c0_exe1224_inputs_ready;
wire local_bb6_c0_exe1224_stall_local;
wire local_bb6_c0_exe1224;

assign local_bb6_c0_exe1224_inputs_ready = local_bb6_c0_exit223_c0_exi3222_valid_out_0_NO_SHIFT_REG;
assign local_bb6_c0_exe1224 = local_bb6_c0_exit223_c0_exi3222_NO_SHIFT_REG[8];
assign local_bb6_c0_exe1224_valid_out = local_bb6_c0_exe1224_inputs_ready;
assign local_bb6_c0_exe1224_stall_local = local_bb6_c0_exe1224_stall_in;
assign local_bb6_c0_exit223_c0_exi3222_stall_in_0 = (|local_bb6_c0_exe1224_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exe2225_valid_out;
wire local_bb6_c0_exe2225_stall_in;
wire local_bb6_c0_exe2225_inputs_ready;
wire local_bb6_c0_exe2225_stall_local;
wire [31:0] local_bb6_c0_exe2225;

assign local_bb6_c0_exe2225_inputs_ready = local_bb6_c0_exit223_c0_exi3222_valid_out_1_NO_SHIFT_REG;
assign local_bb6_c0_exe2225 = local_bb6_c0_exit223_c0_exi3222_NO_SHIFT_REG[63:32];
assign local_bb6_c0_exe2225_valid_out = local_bb6_c0_exe2225_inputs_ready;
assign local_bb6_c0_exe2225_stall_local = local_bb6_c0_exe2225_stall_in;
assign local_bb6_c0_exit223_c0_exi3222_stall_in_1 = (|local_bb6_c0_exe2225_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exe3226_valid_out;
wire local_bb6_c0_exe3226_stall_in;
wire local_bb6_c0_exe3226_inputs_ready;
wire local_bb6_c0_exe3226_stall_local;
wire local_bb6_c0_exe3226;
wire rci_rcnode_21to180_rc0_bb6__arrayidx53_0_reg_21;

assign local_bb6_c0_exe3226_inputs_ready = local_bb6_c0_exit223_c0_exi3222_valid_out_2_NO_SHIFT_REG;
assign local_bb6_c0_exe3226 = local_bb6_c0_exit223_c0_exi3222_NO_SHIFT_REG[64];
assign local_bb6_c0_exe3226_valid_out = local_bb6_c0_exe3226_inputs_ready;
assign local_bb6_c0_exe3226_stall_local = local_bb6_c0_exe3226_stall_in;
assign local_bb6_c0_exit223_c0_exi3222_stall_in_2 = (|local_bb6_c0_exe3226_stall_local);
assign rci_rcnode_21to180_rc0_bb6__arrayidx53_0_reg_21 = local_bb6_c0_exe1224;

// Register node:
//  * latency = 159
//  * capacity = 159
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_valid_out_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_stall_in_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_stall_out_0_reg_180_IP_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx53_0_stall_out_0_reg_180_NO_SHIFT_REG;

acl_data_fifo rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_21to180_rc0_bb6__arrayidx53_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rcnode_21to180_rc0_bb6__arrayidx53_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rcnode_21to180_rc0_bb6__arrayidx53_0_stall_out_0_reg_180_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_21to180_rc0_bb6__arrayidx53_0_reg_21),
	.data_out(rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_NO_SHIFT_REG)
);

defparam rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_fifo.DEPTH = 160;
defparam rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_fifo.IMPL = "ram";

assign rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_inputs_ready_NO_SHIFT_REG = (local_bb6__arrayidx53_valid_out & local_bb6_c0_exe1224_valid_out);
assign rcnode_21to180_rc0_bb6__arrayidx53_0_stall_out_0_reg_180_NO_SHIFT_REG = (~(rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_inputs_ready_NO_SHIFT_REG) | rcnode_21to180_rc0_bb6__arrayidx53_0_stall_out_0_reg_180_IP_NO_SHIFT_REG);
assign local_bb6__arrayidx53_stall_in = rcnode_21to180_rc0_bb6__arrayidx53_0_stall_out_0_reg_180_NO_SHIFT_REG;
assign local_bb6_c0_exe1224_stall_in = rcnode_21to180_rc0_bb6__arrayidx53_0_stall_out_0_reg_180_NO_SHIFT_REG;
assign rcnode_21to180_rc0_bb6__arrayidx53_0_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx53_0_reg_180_NO_SHIFT_REG;
assign rcnode_21to180_rc0_bb6__arrayidx53_0_stall_in_reg_180_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx53_0_stall_in_NO_SHIFT_REG;
assign rcnode_21to180_rc0_bb6__arrayidx53_0_valid_out_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx53_0_valid_out_reg_180_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb6_st_c0_exe2225_inputs_ready;
 reg local_bb6_st_c0_exe2225_valid_out_NO_SHIFT_REG;
wire local_bb6_st_c0_exe2225_stall_in;
wire local_bb6_st_c0_exe2225_output_regs_ready;
wire local_bb6_st_c0_exe2225_fu_stall_out;
wire local_bb6_st_c0_exe2225_fu_valid_out;
wire [31:0] local_bb6_st_c0_exe2225_lsu_wackout;
 reg local_bb6_st_c0_exe2225_NO_SHIFT_REG;
wire local_bb6_st_c0_exe2225_causedstall;
wire rci_rcnode_180to181_rc0_bb6__arrayidx53_0_reg_180;

lsu_top lsu_local_bb6_st_c0_exe2225 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb6_st_c0_exe2225_fu_stall_out),
	.i_valid(local_bb6_st_c0_exe2225_inputs_ready),
	.i_address((rnode_20to21_bb6_arrayidx53_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(local_bb6_c0_exe2225),
	.i_cmpdata(),
	.i_predicate(local_bb6_c0_exe3226),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb6_st_c0_exe2225_output_regs_ready)),
	.o_valid(local_bb6_st_c0_exe2225_fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(local_bb6_st_c0_exe2225_lsu_wackout),
	.i_atomic_op(3'h0),
	.o_active(local_bb6_st_c0_exe2225_active),
	.avm_address(avm_local_bb6_st_c0_exe2225_address),
	.avm_read(avm_local_bb6_st_c0_exe2225_read),
	.avm_readdata(avm_local_bb6_st_c0_exe2225_readdata),
	.avm_write(avm_local_bb6_st_c0_exe2225_write),
	.avm_writeack(avm_local_bb6_st_c0_exe2225_writeack),
	.avm_burstcount(avm_local_bb6_st_c0_exe2225_burstcount),
	.avm_writedata(avm_local_bb6_st_c0_exe2225_writedata),
	.avm_byteenable(avm_local_bb6_st_c0_exe2225_byteenable),
	.avm_waitrequest(avm_local_bb6_st_c0_exe2225_waitrequest),
	.avm_readdatavalid(avm_local_bb6_st_c0_exe2225_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb6_st_c0_exe2225.AWIDTH = 33;
defparam lsu_local_bb6_st_c0_exe2225.WIDTH_BYTES = 4;
defparam lsu_local_bb6_st_c0_exe2225.MWIDTH_BYTES = 64;
defparam lsu_local_bb6_st_c0_exe2225.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb6_st_c0_exe2225.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb6_st_c0_exe2225.READ = 0;
defparam lsu_local_bb6_st_c0_exe2225.ATOMIC = 0;
defparam lsu_local_bb6_st_c0_exe2225.WIDTH = 32;
defparam lsu_local_bb6_st_c0_exe2225.MWIDTH = 512;
defparam lsu_local_bb6_st_c0_exe2225.ATOMIC_WIDTH = 3;
defparam lsu_local_bb6_st_c0_exe2225.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb6_st_c0_exe2225.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb6_st_c0_exe2225.MEMORY_SIDE_MEM_LATENCY = 10;
defparam lsu_local_bb6_st_c0_exe2225.USE_WRITE_ACK = 1;
defparam lsu_local_bb6_st_c0_exe2225.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb6_st_c0_exe2225.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb6_st_c0_exe2225.NUMBER_BANKS = 1;
defparam lsu_local_bb6_st_c0_exe2225.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb6_st_c0_exe2225.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb6_st_c0_exe2225.USEINPUTFIFO = 0;
defparam lsu_local_bb6_st_c0_exe2225.USECACHING = 0;
defparam lsu_local_bb6_st_c0_exe2225.USEOUTPUTFIFO = 1;
defparam lsu_local_bb6_st_c0_exe2225.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb6_st_c0_exe2225.HIGH_FMAX = 1;
defparam lsu_local_bb6_st_c0_exe2225.ADDRSPACE = 1;
defparam lsu_local_bb6_st_c0_exe2225.STYLE = "BURST-COALESCED";
defparam lsu_local_bb6_st_c0_exe2225.USE_BYTE_EN = 0;

assign local_bb6_st_c0_exe2225_inputs_ready = (local_bb6_c0_exe2225_valid_out & local_bb6_c0_exe3226_valid_out & rnode_20to21_bb6_arrayidx53_0_valid_out_0_NO_SHIFT_REG);
assign local_bb6_st_c0_exe2225_output_regs_ready = (&(~(local_bb6_st_c0_exe2225_valid_out_NO_SHIFT_REG) | ~(local_bb6_st_c0_exe2225_stall_in)));
assign local_bb6_c0_exe2225_stall_in = (local_bb6_st_c0_exe2225_fu_stall_out | ~(local_bb6_st_c0_exe2225_inputs_ready));
assign local_bb6_c0_exe3226_stall_in = (local_bb6_st_c0_exe2225_fu_stall_out | ~(local_bb6_st_c0_exe2225_inputs_ready));
assign rnode_20to21_bb6_arrayidx53_0_stall_in_0_NO_SHIFT_REG = (local_bb6_st_c0_exe2225_fu_stall_out | ~(local_bb6_st_c0_exe2225_inputs_ready));
assign local_bb6_st_c0_exe2225_causedstall = (local_bb6_st_c0_exe2225_inputs_ready && (local_bb6_st_c0_exe2225_fu_stall_out && !(~(local_bb6_st_c0_exe2225_output_regs_ready))));
assign rci_rcnode_180to181_rc0_bb6__arrayidx53_0_reg_180 = rcnode_21to180_rc0_bb6__arrayidx53_0_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_st_c0_exe2225_NO_SHIFT_REG <= 'x;
		local_bb6_st_c0_exe2225_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_st_c0_exe2225_output_regs_ready)
		begin
			local_bb6_st_c0_exe2225_NO_SHIFT_REG <= local_bb6_st_c0_exe2225_lsu_wackout;
			local_bb6_st_c0_exe2225_valid_out_NO_SHIFT_REG <= local_bb6_st_c0_exe2225_fu_valid_out;
		end
		else
		begin
			if (~(local_bb6_st_c0_exe2225_stall_in))
			begin
				local_bb6_st_c0_exe2225_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_valid_out_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_stall_in_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_stall_out_reg_181_IP_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx53_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_180to181_rc0_bb6__arrayidx53_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rcnode_180to181_rc0_bb6__arrayidx53_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rcnode_180to181_rc0_bb6__arrayidx53_0_stall_out_reg_181_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_180to181_rc0_bb6__arrayidx53_0_reg_180),
	.data_out(rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_NO_SHIFT_REG)
);

defparam rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_fifo.DEPTH = 1;
defparam rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_fifo.IMPL = "ll_reg";

assign rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_inputs_ready_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx53_0_valid_out_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx53_0_stall_out_reg_181_NO_SHIFT_REG = (~(rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_inputs_ready_NO_SHIFT_REG) | rcnode_180to181_rc0_bb6__arrayidx53_0_stall_out_reg_181_IP_NO_SHIFT_REG);
assign rcnode_21to180_rc0_bb6__arrayidx53_0_stall_in_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx53_0_stall_out_reg_181_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx53_0_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx53_0_reg_181_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx53_0_stall_in_reg_181_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx53_0_stall_in_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx53_0_valid_out_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx53_0_valid_out_reg_181_NO_SHIFT_REG;

// This section implements a staging register.
// 
wire rstag_181to181_bb6_st_c0_exe2225_valid_out;
wire rstag_181to181_bb6_st_c0_exe2225_stall_in;
wire rstag_181to181_bb6_st_c0_exe2225_inputs_ready;
wire rstag_181to181_bb6_st_c0_exe2225_stall_local;
 reg rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG;
wire rstag_181to181_bb6_st_c0_exe2225_combined_valid;
 reg rstag_181to181_bb6_st_c0_exe2225_staging_reg_NO_SHIFT_REG;
wire rstag_181to181_bb6_st_c0_exe2225;

assign rstag_181to181_bb6_st_c0_exe2225_inputs_ready = local_bb6_st_c0_exe2225_valid_out_NO_SHIFT_REG;
assign rstag_181to181_bb6_st_c0_exe2225 = (rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG ? rstag_181to181_bb6_st_c0_exe2225_staging_reg_NO_SHIFT_REG : local_bb6_st_c0_exe2225_NO_SHIFT_REG);
assign rstag_181to181_bb6_st_c0_exe2225_combined_valid = (rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG | rstag_181to181_bb6_st_c0_exe2225_inputs_ready);
assign rstag_181to181_bb6_st_c0_exe2225_valid_out = rstag_181to181_bb6_st_c0_exe2225_combined_valid;
assign rstag_181to181_bb6_st_c0_exe2225_stall_local = rstag_181to181_bb6_st_c0_exe2225_stall_in;
assign local_bb6_st_c0_exe2225_stall_in = (|rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_181to181_bb6_st_c0_exe2225_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_181to181_bb6_st_c0_exe2225_stall_local)
		begin
			if (~(rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG))
			begin
				rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG <= rstag_181to181_bb6_st_c0_exe2225_inputs_ready;
			end
		end
		else
		begin
			rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_181to181_bb6_st_c0_exe2225_staging_valid_NO_SHIFT_REG))
		begin
			rstag_181to181_bb6_st_c0_exe2225_staging_reg_NO_SHIFT_REG <= local_bb6_st_c0_exe2225_NO_SHIFT_REG;
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_bb6_indvars_iv_next31_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb6_indvars_iv_next31_valid_out & rcnode_180to181_rc0_bb6__arrayidx53_0_valid_out_NO_SHIFT_REG & rstag_181to181_bb6_st_c0_exe2225_valid_out);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb6_indvars_iv_next31_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_180to181_rc0_bb6__arrayidx53_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_181to181_bb6_st_c0_exe2225_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb6_indvars_iv_next31_0 = lvb_bb6_indvars_iv_next31_0_reg_NO_SHIFT_REG;
assign lvb_bb6_indvars_iv_next31_1 = lvb_bb6_indvars_iv_next31_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_bb6_indvars_iv_next31_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb6_indvars_iv_next31_0_reg_NO_SHIFT_REG <= local_bb6_indvars_iv_next31;
			branch_compare_result_NO_SHIFT_REG <= rcnode_180to181_rc0_bb6__arrayidx53_0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_7
	(
		input 		clock,
		input 		resetn,
		input 		input_wii_cmp1017,
		input [31:0] 		input_wii_mul39,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u115,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out_0,
		input 		stall_in_0,
		output [63:0] 		lvb_bb7_indvars_iv_next34_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [63:0] 		lvb_bb7_indvars_iv_next34_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		ffwd_2_0,
		input [63:0] 		ffwd_0_0,
		input 		ffwd_6_0,
		output [31:0] 		ffwd_14_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb7_cmp190_acl_ffwd_dest_i1_2_stall_local;
wire local_bb7_cmp190_acl_ffwd_dest_i1_2;

assign local_bb7_cmp190_acl_ffwd_dest_i1_2 = ffwd_2_0;

// This section implements an unregistered operation.
// 
wire local_bb7_indvars_iv33189_acl_ffwd_dest_i64_0_stall_local;
wire [63:0] local_bb7_indvars_iv33189_acl_ffwd_dest_i64_0;

assign local_bb7_indvars_iv33189_acl_ffwd_dest_i64_0 = ffwd_0_0;

// This section implements an unregistered operation.
// 
wire local_bb7__acl_ffwd_dest_i1_6_stall_local;
wire local_bb7__acl_ffwd_dest_i1_6;

assign local_bb7__acl_ffwd_dest_i1_6 = ffwd_6_0;

// This section implements an unregistered operation.
// 
wire local_bb7_var__stall_local;
wire [31:0] local_bb7_var_;

assign local_bb7_var_[31:1] = 31'h0;
assign local_bb7_var_[0] = local_bb7_cmp190_acl_ffwd_dest_i1_2;

// This section implements an unregistered operation.
// 
wire local_bb7_indvars_iv_next34_stall_local;
wire [63:0] local_bb7_indvars_iv_next34;

assign local_bb7_indvars_iv_next34 = (local_bb7_indvars_iv33189_acl_ffwd_dest_i64_0 + 64'h1);

// This section implements an unregistered operation.
// 
wire local_bb7_came_from_for_cond_select_stall_local;
wire [31:0] local_bb7_came_from_for_cond_select;

assign local_bb7_came_from_for_cond_select = ((local_bb7_var_ & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb7_select44_stall_local;
wire [31:0] local_bb7_select44;

assign local_bb7_select44 = (local_bb7__acl_ffwd_dest_i1_6 ? 32'h2 : (local_bb7_came_from_for_cond_select & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb7_for_cond_branch_back_stall_local;
wire local_bb7_for_cond_branch_back;

assign local_bb7_for_cond_branch_back = ((local_bb7_select44 & 32'h3) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb7_for_cond_branch_back_valid_out;
wire local_bb7_for_cond_branch_back_stall_in;
wire local_bb7__select44_valid_out;
wire local_bb7__select44_stall_in;
wire local_bb7_indvars_iv_next34_valid_out;
wire local_bb7_indvars_iv_next34_stall_in;
wire local_bb7__select44_inputs_ready;
wire local_bb7__select44_stall_local;
 reg [31:0] ffwd_14_0_reg_NO_SHIFT_REG;

assign local_bb7__select44_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign ffwd_14_0 = ffwd_14_0_reg_NO_SHIFT_REG;
assign local_bb7__select44_stall_local = (local_bb7_for_cond_branch_back_stall_in | local_bb7__select44_stall_in | local_bb7_indvars_iv_next34_stall_in);
assign local_bb7_for_cond_branch_back_valid_out = local_bb7__select44_inputs_ready;
assign local_bb7__select44_valid_out = local_bb7__select44_inputs_ready;
assign local_bb7_indvars_iv_next34_valid_out = local_bb7__select44_inputs_ready;
assign merge_node_stall_in_0 = (local_bb7__select44_stall_local | ~(local_bb7__select44_inputs_ready));
assign merge_node_stall_in_2 = (local_bb7__select44_stall_local | ~(local_bb7__select44_inputs_ready));
assign merge_node_stall_in_1 = (local_bb7__select44_stall_local | ~(local_bb7__select44_inputs_ready));

always @(posedge clock)
begin
	if ((1'b1 & local_bb7__select44_inputs_ready))
	begin
		ffwd_14_0_reg_NO_SHIFT_REG <= (local_bb7_select44 & 32'h3);
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_bb7_indvars_iv_next34_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb7__select44_valid_out & local_bb7_for_cond_branch_back_valid_out & local_bb7_indvars_iv_next34_valid_out);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb7__select44_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb7_for_cond_branch_back_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb7_indvars_iv_next34_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb7_indvars_iv_next34_0 = lvb_bb7_indvars_iv_next34_0_reg_NO_SHIFT_REG;
assign lvb_bb7_indvars_iv_next34_1 = lvb_bb7_indvars_iv_next34_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_bb7_indvars_iv_next34_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb7_indvars_iv_next34_0_reg_NO_SHIFT_REG <= local_bb7_indvars_iv_next34;
			branch_compare_result_NO_SHIFT_REG <= local_bb7_for_cond_branch_back;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_8
	(
		input 		clock,
		input 		resetn,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start,
		input [31:0] 		ffwd_14_0,
		input [63:0] 		ffwd_13_0,
		input [511:0] 		avm_local_bb8_st__readdata,
		input 		avm_local_bb8_st__readdatavalid,
		input 		avm_local_bb8_st__waitrequest,
		output [32:0] 		avm_local_bb8_st__address,
		output 		avm_local_bb8_st__read,
		output 		avm_local_bb8_st__write,
		input 		avm_local_bb8_st__writeack,
		output [511:0] 		avm_local_bb8_st__writedata,
		output [63:0] 		avm_local_bb8_st__byteenable,
		output [4:0] 		avm_local_bb8_st__burstcount,
		output 		local_bb8_st__active,
		input 		clock2x
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb8_select44198_acl_ffwd_dest_i32_14_stall_local;
wire [31:0] local_bb8_select44198_acl_ffwd_dest_i32_14;

assign local_bb8_select44198_acl_ffwd_dest_i32_14 = ffwd_14_0;

// This section implements an unregistered operation.
// 
wire local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_valid_out;
wire local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_stall_in;
wire local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_inputs_ready;
wire local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_stall_local;
wire [63:0] local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13;

assign local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13 = ffwd_13_0;
assign local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_valid_out = local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_inputs_ready;
assign local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_stall_local = local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_stall_in;
assign merge_node_stall_in_1 = (|local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb8_for_cond_branch_to_dummy_valid_out;
wire local_bb8_for_cond_branch_to_dummy_stall_in;
wire local_bb8_for_cond_branch_to_dummy_inputs_ready;
wire local_bb8_for_cond_branch_to_dummy_stall_local;
wire local_bb8_for_cond_branch_to_dummy;

assign local_bb8_for_cond_branch_to_dummy_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb8_for_cond_branch_to_dummy = (local_bb8_select44198_acl_ffwd_dest_i32_14 == 32'h1);
assign local_bb8_for_cond_branch_to_dummy_valid_out = local_bb8_for_cond_branch_to_dummy_inputs_ready;
assign local_bb8_for_cond_branch_to_dummy_stall_local = local_bb8_for_cond_branch_to_dummy_stall_in;
assign merge_node_stall_in_0 = (|local_bb8_for_cond_branch_to_dummy_stall_local);

// This section implements a registered operation.
// 
wire local_bb8_st__inputs_ready;
 reg local_bb8_st__valid_out_NO_SHIFT_REG;
wire local_bb8_st__stall_in;
wire local_bb8_st__output_regs_ready;
wire local_bb8_st__fu_stall_out;
wire local_bb8_st__fu_valid_out;
wire local_bb8_st__causedstall;

lsu_top lsu_local_bb8_st_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb8_st__fu_stall_out),
	.i_valid(local_bb8_st__inputs_ready),
	.i_address(local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13),
	.i_writedata(32'h0),
	.i_cmpdata(),
	.i_predicate(local_bb8_for_cond_branch_to_dummy),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb8_st__output_regs_ready)),
	.o_valid(local_bb8_st__fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb8_st__active),
	.avm_address(avm_local_bb8_st__address),
	.avm_read(avm_local_bb8_st__read),
	.avm_readdata(avm_local_bb8_st__readdata),
	.avm_write(avm_local_bb8_st__write),
	.avm_writeack(avm_local_bb8_st__writeack),
	.avm_burstcount(avm_local_bb8_st__burstcount),
	.avm_writedata(avm_local_bb8_st__writedata),
	.avm_byteenable(avm_local_bb8_st__byteenable),
	.avm_waitrequest(avm_local_bb8_st__waitrequest),
	.avm_readdatavalid(avm_local_bb8_st__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb8_st_.AWIDTH = 33;
defparam lsu_local_bb8_st_.WIDTH_BYTES = 4;
defparam lsu_local_bb8_st_.MWIDTH_BYTES = 64;
defparam lsu_local_bb8_st_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb8_st_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb8_st_.READ = 0;
defparam lsu_local_bb8_st_.ATOMIC = 0;
defparam lsu_local_bb8_st_.WIDTH = 32;
defparam lsu_local_bb8_st_.MWIDTH = 512;
defparam lsu_local_bb8_st_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb8_st_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb8_st_.KERNEL_SIDE_MEM_LATENCY = 4;
defparam lsu_local_bb8_st_.MEMORY_SIDE_MEM_LATENCY = 10;
defparam lsu_local_bb8_st_.USE_WRITE_ACK = 0;
defparam lsu_local_bb8_st_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb8_st_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb8_st_.NUMBER_BANKS = 1;
defparam lsu_local_bb8_st_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb8_st_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb8_st_.USEINPUTFIFO = 0;
defparam lsu_local_bb8_st_.USECACHING = 0;
defparam lsu_local_bb8_st_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb8_st_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb8_st_.HIGH_FMAX = 1;
defparam lsu_local_bb8_st_.ADDRSPACE = 1;
defparam lsu_local_bb8_st_.STYLE = "BURST-COALESCED";
defparam lsu_local_bb8_st_.USE_BYTE_EN = 0;

assign local_bb8_st__inputs_ready = (local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_valid_out & local_bb8_for_cond_branch_to_dummy_valid_out);
assign local_bb8_st__output_regs_ready = (&(~(local_bb8_st__valid_out_NO_SHIFT_REG) | ~(local_bb8_st__stall_in)));
assign local_bb8_arrayidx53197_acl_ffwd_dest_p1f_13_stall_in = (local_bb8_st__fu_stall_out | ~(local_bb8_st__inputs_ready));
assign local_bb8_for_cond_branch_to_dummy_stall_in = (local_bb8_st__fu_stall_out | ~(local_bb8_st__inputs_ready));
assign local_bb8_st__causedstall = (local_bb8_st__inputs_ready && (local_bb8_st__fu_stall_out && !(~(local_bb8_st__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb8_st__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb8_st__output_regs_ready)
		begin
			local_bb8_st__valid_out_NO_SHIFT_REG <= local_bb8_st__fu_valid_out;
		end
		else
		begin
			if (~(local_bb8_st__stall_in))
			begin
				local_bb8_st__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_5to5_bb8_st__valid_out;
wire rstag_5to5_bb8_st__stall_in;
wire rstag_5to5_bb8_st__inputs_ready;
wire rstag_5to5_bb8_st__stall_local;
 reg rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb8_st__combined_valid;

assign rstag_5to5_bb8_st__inputs_ready = local_bb8_st__valid_out_NO_SHIFT_REG;
assign rstag_5to5_bb8_st__combined_valid = (rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG | rstag_5to5_bb8_st__inputs_ready);
assign rstag_5to5_bb8_st__valid_out = rstag_5to5_bb8_st__combined_valid;
assign rstag_5to5_bb8_st__stall_local = rstag_5to5_bb8_st__stall_in;
assign local_bb8_st__stall_in = (|rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (rstag_5to5_bb8_st__stall_local)
		begin
			if (~(rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG <= rstag_5to5_bb8_st__inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
wire branch_var__output_regs_ready;

assign branch_var__inputs_ready = rstag_5to5_bb8_st__valid_out;
assign branch_var__output_regs_ready = ~(stall_in);
assign rstag_5to5_bb8_st__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out = branch_var__inputs_ready;

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_function
	(
		input 		clock,
		input 		resetn,
		output 		stall_out,
		input 		valid_in,
		output 		valid_out,
		input 		stall_in,
		input [511:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [32:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [511:0] 		avm_local_bb2_ld__writedata,
		output [63:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		input [511:0] 		avm_local_bb4_ld__readdata,
		input 		avm_local_bb4_ld__readdatavalid,
		input 		avm_local_bb4_ld__waitrequest,
		output [32:0] 		avm_local_bb4_ld__address,
		output 		avm_local_bb4_ld__read,
		output 		avm_local_bb4_ld__write,
		input 		avm_local_bb4_ld__writeack,
		output [511:0] 		avm_local_bb4_ld__writedata,
		output [63:0] 		avm_local_bb4_ld__byteenable,
		output [4:0] 		avm_local_bb4_ld__burstcount,
		input [511:0] 		avm_local_bb4_ld__u28_readdata,
		input 		avm_local_bb4_ld__u28_readdatavalid,
		input 		avm_local_bb4_ld__u28_waitrequest,
		output [32:0] 		avm_local_bb4_ld__u28_address,
		output 		avm_local_bb4_ld__u28_read,
		output 		avm_local_bb4_ld__u28_write,
		input 		avm_local_bb4_ld__u28_writeack,
		output [511:0] 		avm_local_bb4_ld__u28_writedata,
		output [63:0] 		avm_local_bb4_ld__u28_byteenable,
		output [4:0] 		avm_local_bb4_ld__u28_burstcount,
		input [511:0] 		avm_local_bb4_ld__u29_readdata,
		input 		avm_local_bb4_ld__u29_readdatavalid,
		input 		avm_local_bb4_ld__u29_waitrequest,
		output [32:0] 		avm_local_bb4_ld__u29_address,
		output 		avm_local_bb4_ld__u29_read,
		output 		avm_local_bb4_ld__u29_write,
		input 		avm_local_bb4_ld__u29_writeack,
		output [511:0] 		avm_local_bb4_ld__u29_writedata,
		output [63:0] 		avm_local_bb4_ld__u29_byteenable,
		output [4:0] 		avm_local_bb4_ld__u29_burstcount,
		input [511:0] 		avm_local_bb6_st_c0_exe2225_readdata,
		input 		avm_local_bb6_st_c0_exe2225_readdatavalid,
		input 		avm_local_bb6_st_c0_exe2225_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe2225_address,
		output 		avm_local_bb6_st_c0_exe2225_read,
		output 		avm_local_bb6_st_c0_exe2225_write,
		input 		avm_local_bb6_st_c0_exe2225_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe2225_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe2225_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe2225_burstcount,
		input [511:0] 		avm_local_bb8_st__readdata,
		input 		avm_local_bb8_st__readdatavalid,
		input 		avm_local_bb8_st__waitrequest,
		output [32:0] 		avm_local_bb8_st__address,
		output 		avm_local_bb8_st__read,
		output 		avm_local_bb8_st__write,
		input 		avm_local_bb8_st__writeack,
		output [511:0] 		avm_local_bb8_st__writedata,
		output [63:0] 		avm_local_bb8_st__byteenable,
		output [4:0] 		avm_local_bb8_st__burstcount,
		input 		start,
		input [31:0] 		input_r,
		input [31:0] 		input_e_d,
		input 		clock2x,
		input [63:0] 		input_in,
		input [63:0] 		input_gaussian,
		input [63:0] 		input_out,
		output reg 		has_a_write_pending,
		output reg 		has_a_lsu_active
	);


wire [31:0] workgroup_size;
wire [31:0] cur_cycle;
wire bb_0_stall_out;
wire bb_0_valid_out;
wire bb_0_lvb_bb0_cmp1017;
wire [31:0] bb_0_lvb_bb0_mul39;
wire [63:0] bb_0_lvb_bb0_var_;
wire [63:0] bb_0_lvb_bb0_var__u0;
wire bb_1_stall_out_0;
wire bb_1_stall_out_1;
wire bb_1_valid_out;
wire [63:0] ffwd_0_0;
wire [31:0] ffwd_1_0;
wire ffwd_2_0;
wire [63:0] ffwd_3_0;
wire bb_2_stall_out_0;
wire bb_2_stall_out_1;
wire bb_2_valid_out;
wire [63:0] ffwd_4_0;
wire [31:0] ffwd_5_0;
wire [63:0] ffwd_7_0;
wire ffwd_6_0;
wire bb_2_local_bb2_ld__active;
wire [31:0] ffwd_8_0;
wire ffwd_9_0;
wire ffwd_10_0;
wire bb_3_stall_out_0;
wire bb_3_stall_out_1;
wire bb_3_valid_out;
wire [31:0] bb_3_lvb_bb3_c0_exe1;
wire [63:0] bb_3_lvb_bb3_c0_exe2;
wire bb_3_lvb_bb3_c0_exe3;
wire bb_3_lvb_bb3_c0_exe4;
wire [31:0] bb_3_lvb_bb3_t_219_pop5_;
wire [31:0] bb_3_lvb_bb3_sum_218_pop6_;
wire bb_3_feedback_stall_out_5;
wire bb_3_feedback_stall_out_6;
wire bb_3_feedback_stall_out_4;
wire bb_3_feedback_stall_out_2;
wire bb_3_feedback_stall_out_3;
wire bb_3_acl_pipelined_valid;
wire bb_3_acl_pipelined_exiting_valid;
wire bb_3_acl_pipelined_exiting_stall;
wire bb_3_feedback_valid_out_3;
wire bb_3_feedback_data_out_3;
wire bb_3_feedback_valid_out_4;
wire [63:0] bb_3_feedback_data_out_4;
wire bb_4_stall_out_0;
wire bb_4_stall_out_1;
wire bb_4_valid_out_0;
wire [319:0] bb_4_lvb_bb4_c0_exit214_c0_exi7_0;
wire bb_4_lvb_bb4_c0_exe7_0;
wire [95:0] bb_4_lvb_bb4_c1_exit_c1_exi2_0;
wire bb_4_valid_out_1;
wire [319:0] bb_4_lvb_bb4_c0_exit214_c0_exi7_1;
wire bb_4_lvb_bb4_c0_exe7_1;
wire [95:0] bb_4_lvb_bb4_c1_exit_c1_exi2_1;
wire bb_4_feedback_stall_out_7;
wire bb_4_feedback_stall_out_0;
wire bb_4_feedback_stall_out_1;
wire bb_4_acl_pipelined_valid;
wire bb_4_acl_pipelined_exiting_valid;
wire bb_4_acl_pipelined_exiting_stall;
wire bb_4_feedback_stall_out_10;
wire bb_4_feedback_stall_out_11;
wire bb_4_feedback_stall_out_12;
wire bb_4_feedback_stall_out_13;
wire bb_4_feedback_valid_out_1;
wire bb_4_feedback_data_out_1;
wire bb_4_feedback_valid_out_7;
wire [63:0] bb_4_feedback_data_out_7;
wire bb_4_feedback_valid_out_11;
wire [63:0] bb_4_feedback_data_out_11;
wire bb_4_feedback_valid_out_12;
wire bb_4_feedback_data_out_12;
wire bb_4_feedback_valid_out_13;
wire bb_4_feedback_data_out_13;
wire bb_4_feedback_valid_out_10;
wire [31:0] bb_4_feedback_data_out_10;
wire bb_4_local_bb4_ld__active;
wire bb_4_local_bb4_ld__u28_active;
wire bb_4_local_bb4_ld__u29_active;
wire bb_4_feedback_stall_out_9;
wire bb_4_feedback_stall_out_8;
wire bb_4_feedback_valid_out_9;
wire [31:0] bb_4_feedback_data_out_9;
wire [31:0] ffwd_11_0;
wire bb_4_feedback_valid_out_8;
wire [31:0] bb_4_feedback_data_out_8;
wire [31:0] ffwd_12_0;
wire bb_5_stall_out;
wire bb_5_valid_out_0;
wire bb_5_valid_out_1;
wire bb_5_feedback_valid_out_5;
wire [31:0] bb_5_feedback_data_out_5;
wire bb_5_feedback_valid_out_6;
wire [31:0] bb_5_feedback_data_out_6;
wire bb_6_stall_out;
wire bb_6_valid_out_0;
wire [63:0] bb_6_lvb_bb6_indvars_iv_next31_0;
wire bb_6_valid_out_1;
wire [63:0] bb_6_lvb_bb6_indvars_iv_next31_1;
wire [63:0] ffwd_13_0;
wire bb_6_local_bb6_st_c0_exe2225_active;
wire bb_7_stall_out;
wire bb_7_valid_out_0;
wire [63:0] bb_7_lvb_bb7_indvars_iv_next34_0;
wire bb_7_valid_out_1;
wire [63:0] bb_7_lvb_bb7_indvars_iv_next34_1;
wire [31:0] ffwd_14_0;
wire bb_8_stall_out;
wire bb_8_valid_out;
wire bb_8_local_bb8_st__active;
wire feedback_stall_3;
wire feedback_valid_3;
wire feedback_data_3;
wire feedback_stall_4;
wire feedback_valid_4;
wire [63:0] feedback_data_4;
wire feedback_stall_1;
wire feedback_valid_1;
wire feedback_data_1;
wire feedback_stall_11;
wire feedback_valid_11;
wire [63:0] feedback_data_11;
wire feedback_stall_10;
wire feedback_valid_10;
wire [31:0] feedback_data_10;
wire feedback_stall_7;
wire feedback_valid_7;
wire [63:0] feedback_data_7;
wire feedback_stall_12;
wire feedback_valid_12;
wire feedback_data_12;
wire feedback_stall_13;
wire feedback_valid_13;
wire feedback_data_13;
wire feedback_stall_9;
wire feedback_valid_9;
wire [31:0] feedback_data_9;
wire feedback_stall_8;
wire feedback_valid_8;
wire [31:0] feedback_data_8;
wire feedback_stall_6;
wire feedback_valid_6;
wire [31:0] feedback_data_6;
wire feedback_stall_5;
wire feedback_valid_5;
wire [31:0] feedback_data_5;
wire loop_limiter_1_stall_out;
wire loop_limiter_1_valid_out;
wire loop_limiter_2_stall_out;
wire loop_limiter_2_valid_out;
wire loop_limiter_3_stall_out;
wire loop_limiter_3_valid_out;
wire [1:0] writes_pending;
wire [5:0] lsus_active;

AOCbilateralFilterkernel_basic_block_0 AOCbilateralFilterkernel_basic_block_0 (
	.clock(clock),
	.resetn(resetn),
	.start(start),
	.input_r(input_r),
	.input_e_d(input_e_d),
	.valid_in(valid_in),
	.stall_out(bb_0_stall_out),
	.valid_out(bb_0_valid_out),
	.stall_in(bb_1_stall_out_1),
	.lvb_bb0_cmp1017(bb_0_lvb_bb0_cmp1017),
	.lvb_bb0_mul39(bb_0_lvb_bb0_mul39),
	.lvb_bb0_var_(bb_0_lvb_bb0_var_),
	.lvb_bb0_var__u0(bb_0_lvb_bb0_var__u0),
	.workgroup_size(workgroup_size)
);


AOCbilateralFilterkernel_basic_block_1 AOCbilateralFilterkernel_basic_block_1 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_cmp1017(bb_0_lvb_bb0_cmp1017),
	.input_wii_mul39(bb_0_lvb_bb0_mul39),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u3(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_7_valid_out_0),
	.stall_out_0(bb_1_stall_out_0),
	.input_indvars_iv33_0(bb_7_lvb_bb7_indvars_iv_next34_0),
	.valid_in_1(bb_0_valid_out),
	.stall_out_1(bb_1_stall_out_1),
	.input_indvars_iv33_1(64'h0),
	.valid_out(bb_1_valid_out),
	.stall_in(loop_limiter_1_stall_out),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_0_0(ffwd_0_0),
	.ffwd_1_0(ffwd_1_0),
	.ffwd_2_0(ffwd_2_0),
	.ffwd_3_0(ffwd_3_0)
);


AOCbilateralFilterkernel_basic_block_2 AOCbilateralFilterkernel_basic_block_2 (
	.clock(clock),
	.resetn(resetn),
	.input_in(input_in),
	.input_wii_cmp1017(bb_0_lvb_bb0_cmp1017),
	.input_wii_mul39(bb_0_lvb_bb0_mul39),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u6(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_6_valid_out_0),
	.stall_out_0(bb_2_stall_out_0),
	.input_indvars_iv30_0(bb_6_lvb_bb6_indvars_iv_next31_0),
	.valid_in_1(loop_limiter_1_valid_out),
	.stall_out_1(bb_2_stall_out_1),
	.input_indvars_iv30_1(64'h0),
	.valid_out(bb_2_valid_out),
	.stall_in(loop_limiter_2_stall_out),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_3_0(ffwd_3_0),
	.ffwd_4_0(ffwd_4_0),
	.ffwd_5_0(ffwd_5_0),
	.ffwd_2_0(ffwd_2_0),
	.ffwd_7_0(ffwd_7_0),
	.ffwd_6_0(ffwd_6_0),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__burstcount),
	.local_bb2_ld__active(bb_2_local_bb2_ld__active),
	.clock2x(clock2x),
	.ffwd_8_0(ffwd_8_0),
	.ffwd_9_0(ffwd_9_0),
	.ffwd_10_0(ffwd_10_0)
);


AOCbilateralFilterkernel_basic_block_3 AOCbilateralFilterkernel_basic_block_3 (
	.clock(clock),
	.resetn(resetn),
	.input_gaussian(input_gaussian),
	.input_r(input_r),
	.input_wii_cmp1017(bb_0_lvb_bb0_cmp1017),
	.input_wii_mul39(bb_0_lvb_bb0_mul39),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u15(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_3_acl_pipelined_valid),
	.stall_out_0(bb_3_stall_out_0),
	.input_forked_0(1'b0),
	.valid_in_1(loop_limiter_2_valid_out),
	.stall_out_1(bb_3_stall_out_1),
	.input_forked_1(1'b1),
	.valid_out(bb_3_valid_out),
	.stall_in(loop_limiter_3_stall_out),
	.lvb_bb3_c0_exe1(bb_3_lvb_bb3_c0_exe1),
	.lvb_bb3_c0_exe2(bb_3_lvb_bb3_c0_exe2),
	.lvb_bb3_c0_exe3(bb_3_lvb_bb3_c0_exe3),
	.lvb_bb3_c0_exe4(bb_3_lvb_bb3_c0_exe4),
	.lvb_bb3_t_219_pop5_(bb_3_lvb_bb3_t_219_pop5_),
	.lvb_bb3_sum_218_pop6_(bb_3_lvb_bb3_sum_218_pop6_),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_in_5(feedback_valid_5),
	.feedback_stall_out_5(feedback_stall_5),
	.feedback_data_in_5(feedback_data_5),
	.feedback_valid_in_6(feedback_valid_6),
	.feedback_stall_out_6(feedback_stall_6),
	.feedback_data_in_6(feedback_data_6),
	.feedback_valid_in_4(feedback_valid_4),
	.feedback_stall_out_4(feedback_stall_4),
	.feedback_data_in_4(feedback_data_4),
	.ffwd_10_0(ffwd_10_0),
	.feedback_stall_out_2(bb_3_feedback_stall_out_2),
	.feedback_valid_in_3(feedback_valid_3),
	.feedback_stall_out_3(feedback_stall_3),
	.feedback_data_in_3(feedback_data_3),
	.acl_pipelined_valid(bb_3_acl_pipelined_valid),
	.acl_pipelined_stall(bb_3_stall_out_0),
	.acl_pipelined_exiting_valid(bb_3_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_3_acl_pipelined_exiting_stall),
	.ffwd_5_0(ffwd_5_0),
	.feedback_valid_out_3(feedback_valid_3),
	.feedback_stall_in_3(feedback_stall_3),
	.feedback_data_out_3(feedback_data_3),
	.feedback_valid_out_4(feedback_valid_4),
	.feedback_stall_in_4(feedback_stall_4),
	.feedback_data_out_4(feedback_data_4)
);


AOCbilateralFilterkernel_basic_block_4 AOCbilateralFilterkernel_basic_block_4 (
	.clock(clock),
	.resetn(resetn),
	.input_in(input_in),
	.input_gaussian(input_gaussian),
	.input_r(input_r),
	.input_wii_cmp1017(bb_0_lvb_bb0_cmp1017),
	.input_wii_mul39(bb_0_lvb_bb0_mul39),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u19(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_4_acl_pipelined_valid),
	.stall_out_0(bb_4_stall_out_0),
	.input_t_313_0('x),
	.input_sum_312_0('x),
	.input_forked203_0(1'b0),
	.input_sub17_add16204_0('x),
	.input_arrayidx32205_0('x),
	.input_var__u20_0('x),
	.input_notexitcond201206_0('x),
	.valid_in_1(loop_limiter_3_valid_out),
	.stall_out_1(bb_4_stall_out_1),
	.input_t_313_1(bb_3_lvb_bb3_t_219_pop5_),
	.input_sum_312_1(bb_3_lvb_bb3_sum_218_pop6_),
	.input_forked203_1(1'b1),
	.input_sub17_add16204_1(bb_3_lvb_bb3_c0_exe1),
	.input_arrayidx32205_1(bb_3_lvb_bb3_c0_exe2),
	.input_var__u20_1(bb_3_lvb_bb3_c0_exe3),
	.input_notexitcond201206_1(bb_3_lvb_bb3_c0_exe4),
	.valid_out_0(bb_4_valid_out_0),
	.stall_in_0(bb_5_stall_out),
	.lvb_bb4_c0_exit214_c0_exi7_0(bb_4_lvb_bb4_c0_exit214_c0_exi7_0),
	.lvb_bb4_c0_exe7_0(bb_4_lvb_bb4_c0_exe7_0),
	.lvb_bb4_c1_exit_c1_exi2_0(bb_4_lvb_bb4_c1_exit_c1_exi2_0),
	.valid_out_1(bb_4_valid_out_1),
	.stall_in_1(1'b0),
	.lvb_bb4_c0_exit214_c0_exi7_1(bb_4_lvb_bb4_c0_exit214_c0_exi7_1),
	.lvb_bb4_c0_exe7_1(bb_4_lvb_bb4_c0_exe7_1),
	.lvb_bb4_c1_exit_c1_exi2_1(bb_4_lvb_bb4_c1_exit_c1_exi2_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_10_0(ffwd_10_0),
	.ffwd_1_0(ffwd_1_0),
	.feedback_valid_in_7(feedback_valid_7),
	.feedback_stall_out_7(feedback_stall_7),
	.feedback_data_in_7(feedback_data_7),
	.feedback_stall_out_0(bb_4_feedback_stall_out_0),
	.feedback_valid_in_1(feedback_valid_1),
	.feedback_stall_out_1(feedback_stall_1),
	.feedback_data_in_1(feedback_data_1),
	.acl_pipelined_valid(bb_4_acl_pipelined_valid),
	.acl_pipelined_stall(bb_4_stall_out_0),
	.acl_pipelined_exiting_valid(bb_4_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_4_acl_pipelined_exiting_stall),
	.feedback_valid_in_10(feedback_valid_10),
	.feedback_stall_out_10(feedback_stall_10),
	.feedback_data_in_10(feedback_data_10),
	.feedback_valid_in_11(feedback_valid_11),
	.feedback_stall_out_11(feedback_stall_11),
	.feedback_data_in_11(feedback_data_11),
	.feedback_valid_in_12(feedback_valid_12),
	.feedback_stall_out_12(feedback_stall_12),
	.feedback_data_in_12(feedback_data_12),
	.feedback_valid_in_13(feedback_valid_13),
	.feedback_stall_out_13(feedback_stall_13),
	.feedback_data_in_13(feedback_data_13),
	.feedback_valid_out_1(feedback_valid_1),
	.feedback_stall_in_1(feedback_stall_1),
	.feedback_data_out_1(feedback_data_1),
	.feedback_valid_out_7(feedback_valid_7),
	.feedback_stall_in_7(feedback_stall_7),
	.feedback_data_out_7(feedback_data_7),
	.feedback_valid_out_11(feedback_valid_11),
	.feedback_stall_in_11(feedback_stall_11),
	.feedback_data_out_11(feedback_data_11),
	.feedback_valid_out_12(feedback_valid_12),
	.feedback_stall_in_12(feedback_stall_12),
	.feedback_data_out_12(feedback_data_12),
	.feedback_valid_out_13(feedback_valid_13),
	.feedback_stall_in_13(feedback_stall_13),
	.feedback_data_out_13(feedback_data_13),
	.feedback_valid_out_10(feedback_valid_10),
	.feedback_stall_in_10(feedback_stall_10),
	.feedback_data_out_10(feedback_data_10),
	.avm_local_bb4_ld__readdata(avm_local_bb4_ld__readdata),
	.avm_local_bb4_ld__readdatavalid(avm_local_bb4_ld__readdatavalid),
	.avm_local_bb4_ld__waitrequest(avm_local_bb4_ld__waitrequest),
	.avm_local_bb4_ld__address(avm_local_bb4_ld__address),
	.avm_local_bb4_ld__read(avm_local_bb4_ld__read),
	.avm_local_bb4_ld__write(avm_local_bb4_ld__write),
	.avm_local_bb4_ld__writeack(avm_local_bb4_ld__writeack),
	.avm_local_bb4_ld__writedata(avm_local_bb4_ld__writedata),
	.avm_local_bb4_ld__byteenable(avm_local_bb4_ld__byteenable),
	.avm_local_bb4_ld__burstcount(avm_local_bb4_ld__burstcount),
	.local_bb4_ld__active(bb_4_local_bb4_ld__active),
	.clock2x(clock2x),
	.avm_local_bb4_ld__u28_readdata(avm_local_bb4_ld__u28_readdata),
	.avm_local_bb4_ld__u28_readdatavalid(avm_local_bb4_ld__u28_readdatavalid),
	.avm_local_bb4_ld__u28_waitrequest(avm_local_bb4_ld__u28_waitrequest),
	.avm_local_bb4_ld__u28_address(avm_local_bb4_ld__u28_address),
	.avm_local_bb4_ld__u28_read(avm_local_bb4_ld__u28_read),
	.avm_local_bb4_ld__u28_write(avm_local_bb4_ld__u28_write),
	.avm_local_bb4_ld__u28_writeack(avm_local_bb4_ld__u28_writeack),
	.avm_local_bb4_ld__u28_writedata(avm_local_bb4_ld__u28_writedata),
	.avm_local_bb4_ld__u28_byteenable(avm_local_bb4_ld__u28_byteenable),
	.avm_local_bb4_ld__u28_burstcount(avm_local_bb4_ld__u28_burstcount),
	.local_bb4_ld__u28_active(bb_4_local_bb4_ld__u28_active),
	.avm_local_bb4_ld__u29_readdata(avm_local_bb4_ld__u29_readdata),
	.avm_local_bb4_ld__u29_readdatavalid(avm_local_bb4_ld__u29_readdatavalid),
	.avm_local_bb4_ld__u29_waitrequest(avm_local_bb4_ld__u29_waitrequest),
	.avm_local_bb4_ld__u29_address(avm_local_bb4_ld__u29_address),
	.avm_local_bb4_ld__u29_read(avm_local_bb4_ld__u29_read),
	.avm_local_bb4_ld__u29_write(avm_local_bb4_ld__u29_write),
	.avm_local_bb4_ld__u29_writeack(avm_local_bb4_ld__u29_writeack),
	.avm_local_bb4_ld__u29_writedata(avm_local_bb4_ld__u29_writedata),
	.avm_local_bb4_ld__u29_byteenable(avm_local_bb4_ld__u29_byteenable),
	.avm_local_bb4_ld__u29_burstcount(avm_local_bb4_ld__u29_burstcount),
	.local_bb4_ld__u29_active(bb_4_local_bb4_ld__u29_active),
	.ffwd_8_0(ffwd_8_0),
	.feedback_valid_in_9(feedback_valid_9),
	.feedback_stall_out_9(feedback_stall_9),
	.feedback_data_in_9(feedback_data_9),
	.feedback_valid_in_8(feedback_valid_8),
	.feedback_stall_out_8(feedback_stall_8),
	.feedback_data_in_8(feedback_data_8),
	.feedback_valid_out_9(feedback_valid_9),
	.feedback_stall_in_9(feedback_stall_9),
	.feedback_data_out_9(feedback_data_9),
	.ffwd_11_0(ffwd_11_0),
	.feedback_valid_out_8(feedback_valid_8),
	.feedback_stall_in_8(feedback_stall_8),
	.feedback_data_out_8(feedback_data_8),
	.ffwd_12_0(ffwd_12_0)
);


AOCbilateralFilterkernel_basic_block_5 AOCbilateralFilterkernel_basic_block_5 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_cmp1017(bb_0_lvb_bb0_cmp1017),
	.input_wii_mul39(bb_0_lvb_bb0_mul39),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u111(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_4_valid_out_0),
	.stall_out(bb_5_stall_out),
	.input_c0_exit214_c0_exi7(bb_4_lvb_bb4_c0_exit214_c0_exi7_0),
	.input_c0_exe7(bb_4_lvb_bb4_c0_exe7_0),
	.input_c1_exit_c1_exi2(bb_4_lvb_bb4_c1_exit_c1_exi2_0),
	.valid_out_0(bb_5_valid_out_0),
	.stall_in_0(bb_6_stall_out),
	.valid_out_1(bb_5_valid_out_1),
	.stall_in_1(1'b0),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_out_5(feedback_valid_5),
	.feedback_stall_in_5(feedback_stall_5),
	.feedback_data_out_5(feedback_data_5),
	.feedback_valid_out_6(feedback_valid_6),
	.feedback_stall_in_6(feedback_stall_6),
	.feedback_data_out_6(feedback_data_6)
);


AOCbilateralFilterkernel_basic_block_6 AOCbilateralFilterkernel_basic_block_6 (
	.clock(clock),
	.resetn(resetn),
	.input_out(input_out),
	.input_wii_cmp1017(bb_0_lvb_bb0_cmp1017),
	.input_wii_mul39(bb_0_lvb_bb0_mul39),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u112(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_5_valid_out_0),
	.stall_out(bb_6_stall_out),
	.valid_out_0(bb_6_valid_out_0),
	.stall_in_0(bb_2_stall_out_0),
	.lvb_bb6_indvars_iv_next31_0(bb_6_lvb_bb6_indvars_iv_next31_0),
	.valid_out_1(bb_6_valid_out_1),
	.stall_in_1(bb_7_stall_out),
	.lvb_bb6_indvars_iv_next31_1(bb_6_lvb_bb6_indvars_iv_next31_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_10_0(ffwd_10_0),
	.ffwd_6_0(ffwd_6_0),
	.ffwd_12_0(ffwd_12_0),
	.ffwd_11_0(ffwd_11_0),
	.ffwd_7_0(ffwd_7_0),
	.ffwd_4_0(ffwd_4_0),
	.ffwd_9_0(ffwd_9_0),
	.ffwd_13_0(ffwd_13_0),
	.avm_local_bb6_st_c0_exe2225_readdata(avm_local_bb6_st_c0_exe2225_readdata),
	.avm_local_bb6_st_c0_exe2225_readdatavalid(avm_local_bb6_st_c0_exe2225_readdatavalid),
	.avm_local_bb6_st_c0_exe2225_waitrequest(avm_local_bb6_st_c0_exe2225_waitrequest),
	.avm_local_bb6_st_c0_exe2225_address(avm_local_bb6_st_c0_exe2225_address),
	.avm_local_bb6_st_c0_exe2225_read(avm_local_bb6_st_c0_exe2225_read),
	.avm_local_bb6_st_c0_exe2225_write(avm_local_bb6_st_c0_exe2225_write),
	.avm_local_bb6_st_c0_exe2225_writeack(avm_local_bb6_st_c0_exe2225_writeack),
	.avm_local_bb6_st_c0_exe2225_writedata(avm_local_bb6_st_c0_exe2225_writedata),
	.avm_local_bb6_st_c0_exe2225_byteenable(avm_local_bb6_st_c0_exe2225_byteenable),
	.avm_local_bb6_st_c0_exe2225_burstcount(avm_local_bb6_st_c0_exe2225_burstcount),
	.local_bb6_st_c0_exe2225_active(bb_6_local_bb6_st_c0_exe2225_active),
	.clock2x(clock2x)
);


AOCbilateralFilterkernel_basic_block_7 AOCbilateralFilterkernel_basic_block_7 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_cmp1017(bb_0_lvb_bb0_cmp1017),
	.input_wii_mul39(bb_0_lvb_bb0_mul39),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u115(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_6_valid_out_1),
	.stall_out(bb_7_stall_out),
	.valid_out_0(bb_7_valid_out_0),
	.stall_in_0(bb_1_stall_out_0),
	.lvb_bb7_indvars_iv_next34_0(bb_7_lvb_bb7_indvars_iv_next34_0),
	.valid_out_1(bb_7_valid_out_1),
	.stall_in_1(bb_8_stall_out),
	.lvb_bb7_indvars_iv_next34_1(bb_7_lvb_bb7_indvars_iv_next34_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_2_0(ffwd_2_0),
	.ffwd_0_0(ffwd_0_0),
	.ffwd_6_0(ffwd_6_0),
	.ffwd_14_0(ffwd_14_0)
);


AOCbilateralFilterkernel_basic_block_8 AOCbilateralFilterkernel_basic_block_8 (
	.clock(clock),
	.resetn(resetn),
	.valid_in(bb_7_valid_out_1),
	.stall_out(bb_8_stall_out),
	.valid_out(bb_8_valid_out),
	.stall_in(stall_in),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_14_0(ffwd_14_0),
	.ffwd_13_0(ffwd_13_0),
	.avm_local_bb8_st__readdata(avm_local_bb8_st__readdata),
	.avm_local_bb8_st__readdatavalid(avm_local_bb8_st__readdatavalid),
	.avm_local_bb8_st__waitrequest(avm_local_bb8_st__waitrequest),
	.avm_local_bb8_st__address(avm_local_bb8_st__address),
	.avm_local_bb8_st__read(avm_local_bb8_st__read),
	.avm_local_bb8_st__write(avm_local_bb8_st__write),
	.avm_local_bb8_st__writeack(avm_local_bb8_st__writeack),
	.avm_local_bb8_st__writedata(avm_local_bb8_st__writedata),
	.avm_local_bb8_st__byteenable(avm_local_bb8_st__byteenable),
	.avm_local_bb8_st__burstcount(avm_local_bb8_st__burstcount),
	.local_bb8_st__active(bb_8_local_bb8_st__active),
	.clock2x(clock2x)
);


acl_loop_limiter loop_limiter_1 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_1_valid_out),
	.i_stall(bb_2_stall_out_1),
	.i_valid_exit(bb_6_valid_out_1),
	.i_stall_exit(bb_7_stall_out),
	.o_valid(loop_limiter_1_valid_out),
	.o_stall(loop_limiter_1_stall_out)
);

defparam loop_limiter_1.ENTRY_WIDTH = 1;
defparam loop_limiter_1.EXIT_WIDTH = 1;
defparam loop_limiter_1.THRESHOLD = 772;

acl_loop_limiter loop_limiter_2 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_2_valid_out),
	.i_stall(bb_3_stall_out_1),
	.i_valid_exit(bb_3_acl_pipelined_exiting_valid),
	.i_stall_exit(bb_3_acl_pipelined_exiting_stall),
	.o_valid(loop_limiter_2_valid_out),
	.o_stall(loop_limiter_2_stall_out)
);

defparam loop_limiter_2.ENTRY_WIDTH = 1;
defparam loop_limiter_2.EXIT_WIDTH = 1;
defparam loop_limiter_2.THRESHOLD = 2;

acl_loop_limiter loop_limiter_3 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_3_valid_out),
	.i_stall(bb_4_stall_out_1),
	.i_valid_exit(bb_4_acl_pipelined_exiting_valid),
	.i_stall_exit(bb_4_acl_pipelined_exiting_stall),
	.o_valid(loop_limiter_3_valid_out),
	.o_stall(loop_limiter_3_stall_out)
);

defparam loop_limiter_3.ENTRY_WIDTH = 1;
defparam loop_limiter_3.EXIT_WIDTH = 1;
defparam loop_limiter_3.THRESHOLD = 9;

AOCbilateralFilterkernel_sys_cycle_time system_cycle_time_module (
	.clock(clock),
	.resetn(resetn),
	.cur_cycle(cur_cycle)
);


assign workgroup_size = 32'h1;
assign valid_out = bb_8_valid_out;
assign stall_out = bb_0_stall_out;
assign writes_pending[0] = bb_6_local_bb6_st_c0_exe2225_active;
assign writes_pending[1] = bb_8_local_bb8_st__active;
assign lsus_active[0] = bb_2_local_bb2_ld__active;
assign lsus_active[1] = bb_4_local_bb4_ld__active;
assign lsus_active[2] = bb_4_local_bb4_ld__u28_active;
assign lsus_active[3] = bb_4_local_bb4_ld__u29_active;
assign lsus_active[4] = bb_6_local_bb6_st_c0_exe2225_active;
assign lsus_active[5] = bb_8_local_bb8_st__active;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		has_a_write_pending <= 1'b0;
		has_a_lsu_active <= 1'b0;
	end
	else
	begin
		has_a_write_pending <= (|writes_pending);
		has_a_lsu_active <= (|lsus_active);
	end
end

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_function_wrapper
	(
		input 		clock,
		input 		resetn,
		input 		clock2x,
		input 		local_router_hang,
		input 		avs_cra_read,
		input 		avs_cra_write,
		input [4:0] 		avs_cra_address,
		input [63:0] 		avs_cra_writedata,
		input [7:0] 		avs_cra_byteenable,
		output reg [63:0] 		avs_cra_readdata,
		output reg 		avs_cra_readdatavalid,
		output 		cra_irq,
		input [511:0] 		avm_local_bb2_ld__inst0_readdata,
		input 		avm_local_bb2_ld__inst0_readdatavalid,
		input 		avm_local_bb2_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb2_ld__inst0_address,
		output 		avm_local_bb2_ld__inst0_read,
		output 		avm_local_bb2_ld__inst0_write,
		input 		avm_local_bb2_ld__inst0_writeack,
		output [511:0] 		avm_local_bb2_ld__inst0_writedata,
		output [63:0] 		avm_local_bb2_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb4_ld__inst0_readdata,
		input 		avm_local_bb4_ld__inst0_readdatavalid,
		input 		avm_local_bb4_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb4_ld__inst0_address,
		output 		avm_local_bb4_ld__inst0_read,
		output 		avm_local_bb4_ld__inst0_write,
		input 		avm_local_bb4_ld__inst0_writeack,
		output [511:0] 		avm_local_bb4_ld__inst0_writedata,
		output [63:0] 		avm_local_bb4_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb4_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb4_ld__u28_inst0_readdata,
		input 		avm_local_bb4_ld__u28_inst0_readdatavalid,
		input 		avm_local_bb4_ld__u28_inst0_waitrequest,
		output [32:0] 		avm_local_bb4_ld__u28_inst0_address,
		output 		avm_local_bb4_ld__u28_inst0_read,
		output 		avm_local_bb4_ld__u28_inst0_write,
		input 		avm_local_bb4_ld__u28_inst0_writeack,
		output [511:0] 		avm_local_bb4_ld__u28_inst0_writedata,
		output [63:0] 		avm_local_bb4_ld__u28_inst0_byteenable,
		output [4:0] 		avm_local_bb4_ld__u28_inst0_burstcount,
		input [511:0] 		avm_local_bb4_ld__u29_inst0_readdata,
		input 		avm_local_bb4_ld__u29_inst0_readdatavalid,
		input 		avm_local_bb4_ld__u29_inst0_waitrequest,
		output [32:0] 		avm_local_bb4_ld__u29_inst0_address,
		output 		avm_local_bb4_ld__u29_inst0_read,
		output 		avm_local_bb4_ld__u29_inst0_write,
		input 		avm_local_bb4_ld__u29_inst0_writeack,
		output [511:0] 		avm_local_bb4_ld__u29_inst0_writedata,
		output [63:0] 		avm_local_bb4_ld__u29_inst0_byteenable,
		output [4:0] 		avm_local_bb4_ld__u29_inst0_burstcount,
		input [511:0] 		avm_local_bb6_st_c0_exe2225_inst0_readdata,
		input 		avm_local_bb6_st_c0_exe2225_inst0_readdatavalid,
		input 		avm_local_bb6_st_c0_exe2225_inst0_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe2225_inst0_address,
		output 		avm_local_bb6_st_c0_exe2225_inst0_read,
		output 		avm_local_bb6_st_c0_exe2225_inst0_write,
		input 		avm_local_bb6_st_c0_exe2225_inst0_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe2225_inst0_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe2225_inst0_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe2225_inst0_burstcount,
		input [511:0] 		avm_local_bb8_st__inst0_readdata,
		input 		avm_local_bb8_st__inst0_readdatavalid,
		input 		avm_local_bb8_st__inst0_waitrequest,
		output [32:0] 		avm_local_bb8_st__inst0_address,
		output 		avm_local_bb8_st__inst0_read,
		output 		avm_local_bb8_st__inst0_write,
		input 		avm_local_bb8_st__inst0_writeack,
		output [511:0] 		avm_local_bb8_st__inst0_writedata,
		output [63:0] 		avm_local_bb8_st__inst0_byteenable,
		output [4:0] 		avm_local_bb8_st__inst0_burstcount
	);

// Responsible for interfacing a kernel with the outside world. It comprises a
// slave interface to specify the kernel arguments and retain kernel status. 

// This section of the wrapper implements the slave interface.
// twoXclock_consumer uses clock2x, even if nobody inside the kernel does. Keeps interface to acl_iface consistent for all kernels.
 reg start_NO_SHIFT_REG;
 reg started_NO_SHIFT_REG;
wire finish;
 reg [31:0] status_NO_SHIFT_REG;
wire has_a_write_pending;
wire has_a_lsu_active;
 reg [255:0] kernel_arguments_NO_SHIFT_REG;
 reg twoXclock_consumer_NO_SHIFT_REG /* synthesis  preserve  noprune  */;
 reg [31:0] workgroup_size_NO_SHIFT_REG;
 reg [31:0] global_size_NO_SHIFT_REG[2:0];
 reg [31:0] num_groups_NO_SHIFT_REG[2:0];
 reg [31:0] local_size_NO_SHIFT_REG[2:0];
 reg [31:0] work_dim_NO_SHIFT_REG;
 reg [31:0] global_offset_NO_SHIFT_REG[2:0];
 reg [63:0] profile_data_NO_SHIFT_REG;
 reg [31:0] profile_ctrl_NO_SHIFT_REG;
 reg [63:0] profile_start_cycle_NO_SHIFT_REG;
 reg [63:0] profile_stop_cycle_NO_SHIFT_REG;
wire dispatched_all_groups;
wire [31:0] group_id_tmp[2:0];
wire [31:0] global_id_base_out[2:0];
wire start_out;
wire [31:0] local_id[0:0][2:0];
wire [31:0] global_id[0:0][2:0];
wire [31:0] group_id[0:0][2:0];
wire iter_valid_in;
wire iter_stall_out;
wire stall_in;
wire stall_out;
wire valid_in;
wire valid_out;

always @(posedge clock2x or negedge resetn)
begin
	if (~(resetn))
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b1;
	end
end



// Work group dispatcher is responsible for issuing work-groups to id iterator(s)
acl_work_group_dispatcher group_dispatcher (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.num_groups(num_groups_NO_SHIFT_REG),
	.local_size(local_size_NO_SHIFT_REG),
	.stall_in(iter_stall_out),
	.valid_out(iter_valid_in),
	.group_id_out(group_id_tmp),
	.global_id_base_out(global_id_base_out),
	.start_out(start_out),
	.dispatched_all_groups(dispatched_all_groups)
);

defparam group_dispatcher.NUM_COPIES = 1;
defparam group_dispatcher.RUN_FOREVER = 0;


// This section of the wrapper implements an Avalon Slave Interface used to configure a kernel invocation.
// The few words words contain the status and the workgroup size registers.
// The remaining addressable space is reserved for kernel arguments.
 reg [63:0] cra_readdata_st1_NO_SHIFT_REG;
 reg [4:0] cra_addr_st1_NO_SHIFT_REG;
 reg cra_read_st1_NO_SHIFT_REG;
wire [63:0] bitenable;

assign bitenable[7:0] = (avs_cra_byteenable[0] ? 8'hFF : 8'h0);
assign bitenable[15:8] = (avs_cra_byteenable[1] ? 8'hFF : 8'h0);
assign bitenable[23:16] = (avs_cra_byteenable[2] ? 8'hFF : 8'h0);
assign bitenable[31:24] = (avs_cra_byteenable[3] ? 8'hFF : 8'h0);
assign bitenable[39:32] = (avs_cra_byteenable[4] ? 8'hFF : 8'h0);
assign bitenable[47:40] = (avs_cra_byteenable[5] ? 8'hFF : 8'h0);
assign bitenable[55:48] = (avs_cra_byteenable[6] ? 8'hFF : 8'h0);
assign bitenable[63:56] = (avs_cra_byteenable[7] ? 8'hFF : 8'h0);
assign cra_irq = (status_NO_SHIFT_REG[1] | status_NO_SHIFT_REG[3]);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		start_NO_SHIFT_REG <= 1'b0;
		started_NO_SHIFT_REG <= 1'b0;
		kernel_arguments_NO_SHIFT_REG <= 256'h0;
		status_NO_SHIFT_REG <= 32'h30000;
		profile_ctrl_NO_SHIFT_REG <= 32'h4;
		profile_start_cycle_NO_SHIFT_REG <= 64'h0;
		profile_stop_cycle_NO_SHIFT_REG <= 64'hFFFFFFFFFFFFFFFF;
		work_dim_NO_SHIFT_REG <= 32'h0;
		workgroup_size_NO_SHIFT_REG <= 32'h0;
		global_size_NO_SHIFT_REG[0] <= 32'h0;
		global_size_NO_SHIFT_REG[1] <= 32'h0;
		global_size_NO_SHIFT_REG[2] <= 32'h0;
		num_groups_NO_SHIFT_REG[0] <= 32'h0;
		num_groups_NO_SHIFT_REG[1] <= 32'h0;
		num_groups_NO_SHIFT_REG[2] <= 32'h0;
		local_size_NO_SHIFT_REG[0] <= 32'h0;
		local_size_NO_SHIFT_REG[1] <= 32'h0;
		local_size_NO_SHIFT_REG[2] <= 32'h0;
		global_offset_NO_SHIFT_REG[0] <= 32'h0;
		global_offset_NO_SHIFT_REG[1] <= 32'h0;
		global_offset_NO_SHIFT_REG[2] <= 32'h0;
	end
	else
	begin
		if (avs_cra_write)
		begin
			case (avs_cra_address)
				5'h0:
				begin
					status_NO_SHIFT_REG[31:16] <= 16'h3;
					status_NO_SHIFT_REG[15:0] <= ((status_NO_SHIFT_REG[15:0] & ~(bitenable[15:0])) | (avs_cra_writedata[15:0] & bitenable[15:0]));
				end

				5'h1:
				begin
					profile_ctrl_NO_SHIFT_REG <= ((profile_ctrl_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h3:
				begin
					profile_start_cycle_NO_SHIFT_REG[31:0] <= ((profile_start_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_start_cycle_NO_SHIFT_REG[63:32] <= ((profile_start_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h4:
				begin
					profile_stop_cycle_NO_SHIFT_REG[31:0] <= ((profile_stop_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_stop_cycle_NO_SHIFT_REG[63:32] <= ((profile_stop_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h5:
				begin
					work_dim_NO_SHIFT_REG <= ((work_dim_NO_SHIFT_REG & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					workgroup_size_NO_SHIFT_REG <= ((workgroup_size_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h6:
				begin
					global_size_NO_SHIFT_REG[0] <= ((global_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_size_NO_SHIFT_REG[1] <= ((global_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h7:
				begin
					global_size_NO_SHIFT_REG[2] <= ((global_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[0] <= ((num_groups_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h8:
				begin
					num_groups_NO_SHIFT_REG[1] <= ((num_groups_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[2] <= ((num_groups_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h9:
				begin
					local_size_NO_SHIFT_REG[0] <= ((local_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					local_size_NO_SHIFT_REG[1] <= ((local_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hA:
				begin
					local_size_NO_SHIFT_REG[2] <= ((local_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[0] <= ((global_offset_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hB:
				begin
					global_offset_NO_SHIFT_REG[1] <= ((global_offset_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[2] <= ((global_offset_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hC:
				begin
					kernel_arguments_NO_SHIFT_REG[31:0] <= ((kernel_arguments_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[63:32] <= ((kernel_arguments_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hD:
				begin
					kernel_arguments_NO_SHIFT_REG[95:64] <= ((kernel_arguments_NO_SHIFT_REG[95:64] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[127:96] <= ((kernel_arguments_NO_SHIFT_REG[127:96] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hE:
				begin
					kernel_arguments_NO_SHIFT_REG[159:128] <= ((kernel_arguments_NO_SHIFT_REG[159:128] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[191:160] <= ((kernel_arguments_NO_SHIFT_REG[191:160] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hF:
				begin
					kernel_arguments_NO_SHIFT_REG[223:192] <= ((kernel_arguments_NO_SHIFT_REG[223:192] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[255:224] <= ((kernel_arguments_NO_SHIFT_REG[255:224] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				default:
				begin
				end

			endcase
		end
		else
		begin
			if (status_NO_SHIFT_REG[0])
			begin
				start_NO_SHIFT_REG <= 1'b1;
			end
			if (start_NO_SHIFT_REG)
			begin
				status_NO_SHIFT_REG[0] <= 1'b0;
				started_NO_SHIFT_REG <= 1'b1;
			end
			if (started_NO_SHIFT_REG)
			begin
				start_NO_SHIFT_REG <= 1'b0;
			end
			if (finish)
			begin
				status_NO_SHIFT_REG[1] <= 1'b1;
				started_NO_SHIFT_REG <= 1'b0;
			end
		end
		status_NO_SHIFT_REG[11] <= 1'b0;
		status_NO_SHIFT_REG[12] <= (|has_a_lsu_active);
		status_NO_SHIFT_REG[13] <= (|has_a_write_pending);
		status_NO_SHIFT_REG[14] <= (|valid_in);
		status_NO_SHIFT_REG[15] <= started_NO_SHIFT_REG;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cra_read_st1_NO_SHIFT_REG <= 1'b0;
		cra_addr_st1_NO_SHIFT_REG <= 5'h0;
		cra_readdata_st1_NO_SHIFT_REG <= 64'h0;
	end
	else
	begin
		cra_read_st1_NO_SHIFT_REG <= avs_cra_read;
		cra_addr_st1_NO_SHIFT_REG <= avs_cra_address;
		case (avs_cra_address)
			5'h0:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= status_NO_SHIFT_REG;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			5'h1:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= 'x;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			5'h2:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			5'h3:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			5'h4:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			default:
			begin
				cra_readdata_st1_NO_SHIFT_REG <= status_NO_SHIFT_REG;
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		avs_cra_readdatavalid <= 1'b0;
		avs_cra_readdata <= 64'h0;
	end
	else
	begin
		avs_cra_readdatavalid <= cra_read_st1_NO_SHIFT_REG;
		case (cra_addr_st1_NO_SHIFT_REG)
			5'h2:
			begin
				avs_cra_readdata[63:0] <= profile_data_NO_SHIFT_REG;
			end

			default:
			begin
				avs_cra_readdata <= cra_readdata_st1_NO_SHIFT_REG;
			end

		endcase
	end
end


// Handshaking signals used to control data through the pipeline

// Determine when the kernel is finished.
acl_kernel_finish_detector kernel_finish_detector (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.wg_size(workgroup_size_NO_SHIFT_REG),
	.wg_dispatch_valid_out(iter_valid_in),
	.wg_dispatch_stall_in(iter_stall_out),
	.dispatched_all_groups(dispatched_all_groups),
	.kernel_copy_valid_out(valid_out),
	.kernel_copy_stall_in(stall_in),
	.pending_writes(has_a_write_pending),
	.finish(finish)
);

defparam kernel_finish_detector.TESSELLATION_SIZE = 0;
defparam kernel_finish_detector.NUM_COPIES = 1;
defparam kernel_finish_detector.WG_SIZE_W = 32;

assign stall_in = 1'b0;

// Creating ID iterator and kernel instance for every requested kernel copy

// ID iterator is responsible for iterating over all local ids for given work-groups
acl_id_iterator id_iter_inst0 (
	.clock(clock),
	.resetn(resetn),
	.start(start_out),
	.valid_in(iter_valid_in),
	.stall_out(iter_stall_out),
	.stall_in(stall_out),
	.valid_out(valid_in),
	.group_id_in(group_id_tmp),
	.global_id_base_in(global_id_base_out),
	.local_size(local_size_NO_SHIFT_REG),
	.global_size(global_size_NO_SHIFT_REG),
	.local_id(local_id[0]),
	.global_id(global_id[0]),
	.group_id(group_id[0])
);



// This section instantiates a kernel function block
AOCbilateralFilterkernel_function AOCbilateralFilterkernel_function_inst0 (
	.clock(clock),
	.resetn(resetn),
	.stall_out(stall_out),
	.valid_in(valid_in),
	.valid_out(valid_out),
	.stall_in(stall_in),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__inst0_readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__inst0_readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__inst0_waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__inst0_address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__inst0_read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__inst0_write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__inst0_writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__inst0_writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__inst0_byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__inst0_burstcount),
	.avm_local_bb4_ld__readdata(avm_local_bb4_ld__inst0_readdata),
	.avm_local_bb4_ld__readdatavalid(avm_local_bb4_ld__inst0_readdatavalid),
	.avm_local_bb4_ld__waitrequest(avm_local_bb4_ld__inst0_waitrequest),
	.avm_local_bb4_ld__address(avm_local_bb4_ld__inst0_address),
	.avm_local_bb4_ld__read(avm_local_bb4_ld__inst0_read),
	.avm_local_bb4_ld__write(avm_local_bb4_ld__inst0_write),
	.avm_local_bb4_ld__writeack(avm_local_bb4_ld__inst0_writeack),
	.avm_local_bb4_ld__writedata(avm_local_bb4_ld__inst0_writedata),
	.avm_local_bb4_ld__byteenable(avm_local_bb4_ld__inst0_byteenable),
	.avm_local_bb4_ld__burstcount(avm_local_bb4_ld__inst0_burstcount),
	.avm_local_bb4_ld__u28_readdata(avm_local_bb4_ld__u28_inst0_readdata),
	.avm_local_bb4_ld__u28_readdatavalid(avm_local_bb4_ld__u28_inst0_readdatavalid),
	.avm_local_bb4_ld__u28_waitrequest(avm_local_bb4_ld__u28_inst0_waitrequest),
	.avm_local_bb4_ld__u28_address(avm_local_bb4_ld__u28_inst0_address),
	.avm_local_bb4_ld__u28_read(avm_local_bb4_ld__u28_inst0_read),
	.avm_local_bb4_ld__u28_write(avm_local_bb4_ld__u28_inst0_write),
	.avm_local_bb4_ld__u28_writeack(avm_local_bb4_ld__u28_inst0_writeack),
	.avm_local_bb4_ld__u28_writedata(avm_local_bb4_ld__u28_inst0_writedata),
	.avm_local_bb4_ld__u28_byteenable(avm_local_bb4_ld__u28_inst0_byteenable),
	.avm_local_bb4_ld__u28_burstcount(avm_local_bb4_ld__u28_inst0_burstcount),
	.avm_local_bb4_ld__u29_readdata(avm_local_bb4_ld__u29_inst0_readdata),
	.avm_local_bb4_ld__u29_readdatavalid(avm_local_bb4_ld__u29_inst0_readdatavalid),
	.avm_local_bb4_ld__u29_waitrequest(avm_local_bb4_ld__u29_inst0_waitrequest),
	.avm_local_bb4_ld__u29_address(avm_local_bb4_ld__u29_inst0_address),
	.avm_local_bb4_ld__u29_read(avm_local_bb4_ld__u29_inst0_read),
	.avm_local_bb4_ld__u29_write(avm_local_bb4_ld__u29_inst0_write),
	.avm_local_bb4_ld__u29_writeack(avm_local_bb4_ld__u29_inst0_writeack),
	.avm_local_bb4_ld__u29_writedata(avm_local_bb4_ld__u29_inst0_writedata),
	.avm_local_bb4_ld__u29_byteenable(avm_local_bb4_ld__u29_inst0_byteenable),
	.avm_local_bb4_ld__u29_burstcount(avm_local_bb4_ld__u29_inst0_burstcount),
	.avm_local_bb6_st_c0_exe2225_readdata(avm_local_bb6_st_c0_exe2225_inst0_readdata),
	.avm_local_bb6_st_c0_exe2225_readdatavalid(avm_local_bb6_st_c0_exe2225_inst0_readdatavalid),
	.avm_local_bb6_st_c0_exe2225_waitrequest(avm_local_bb6_st_c0_exe2225_inst0_waitrequest),
	.avm_local_bb6_st_c0_exe2225_address(avm_local_bb6_st_c0_exe2225_inst0_address),
	.avm_local_bb6_st_c0_exe2225_read(avm_local_bb6_st_c0_exe2225_inst0_read),
	.avm_local_bb6_st_c0_exe2225_write(avm_local_bb6_st_c0_exe2225_inst0_write),
	.avm_local_bb6_st_c0_exe2225_writeack(avm_local_bb6_st_c0_exe2225_inst0_writeack),
	.avm_local_bb6_st_c0_exe2225_writedata(avm_local_bb6_st_c0_exe2225_inst0_writedata),
	.avm_local_bb6_st_c0_exe2225_byteenable(avm_local_bb6_st_c0_exe2225_inst0_byteenable),
	.avm_local_bb6_st_c0_exe2225_burstcount(avm_local_bb6_st_c0_exe2225_inst0_burstcount),
	.avm_local_bb8_st__readdata(avm_local_bb8_st__inst0_readdata),
	.avm_local_bb8_st__readdatavalid(avm_local_bb8_st__inst0_readdatavalid),
	.avm_local_bb8_st__waitrequest(avm_local_bb8_st__inst0_waitrequest),
	.avm_local_bb8_st__address(avm_local_bb8_st__inst0_address),
	.avm_local_bb8_st__read(avm_local_bb8_st__inst0_read),
	.avm_local_bb8_st__write(avm_local_bb8_st__inst0_write),
	.avm_local_bb8_st__writeack(avm_local_bb8_st__inst0_writeack),
	.avm_local_bb8_st__writedata(avm_local_bb8_st__inst0_writedata),
	.avm_local_bb8_st__byteenable(avm_local_bb8_st__inst0_byteenable),
	.avm_local_bb8_st__burstcount(avm_local_bb8_st__inst0_burstcount),
	.start(start_out),
	.input_r(kernel_arguments_NO_SHIFT_REG[255:224]),
	.input_e_d(kernel_arguments_NO_SHIFT_REG[223:192]),
	.clock2x(clock2x),
	.input_in(kernel_arguments_NO_SHIFT_REG[127:64]),
	.input_gaussian(kernel_arguments_NO_SHIFT_REG[191:128]),
	.input_out(kernel_arguments_NO_SHIFT_REG[63:0]),
	.has_a_write_pending(has_a_write_pending),
	.has_a_lsu_active(has_a_lsu_active)
);



endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_sys_cycle_time
	(
		input 		clock,
		input 		resetn,
		output [31:0] 		cur_cycle
	);


 reg [31:0] cur_count_NO_SHIFT_REG;

assign cur_cycle = cur_count_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cur_count_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		cur_count_NO_SHIFT_REG <= (cur_count_NO_SHIFT_REG + 32'h1);
	end
end

endmodule

