// (C) 1992-2015 Altera Corporation. All rights reserved.                         
// Your use of Altera Corporation's design tools, logic functions and other       
// software and tools, and its AMPP partner logic functions, and any output       
// files any of the foregoing (including device programming or simulation         
// files), and any associated documentation or information are expressly subject  
// to the terms and conditions of the Altera Program License Subscription         
// Agreement, Altera MegaCore Function License Agreement, or other applicable     
// license agreement, including, without limitation, that your use is for the     
// sole purpose of programming logic devices manufactured by Altera and sold by   
// Altera or its authorized distributors.  Please refer to the applicable         
// agreement for further details.                                                 
    

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_0
	(
		input 		clock,
		input 		resetn,
		input 		start,
		input [31:0] 		input_inSize_x,
		input [31:0] 		input_inSize_y,
		input [31:0] 		input_r,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out,
		input 		stall_in,
		output [31:0] 		lvb_bb0_div,
		output [31:0] 		lvb_bb0_div1,
		output 		lvb_bb0_cmp19,
		output [31:0] 		lvb_bb0_add7,
		output [31:0] 		lvb_bb0_sub20,
		output [31:0] 		lvb_bb0_sub22,
		output 		lvb_bb0_var_,
		output 		lvb_bb0_var__u0,
		output 		lvb_bb0_var__u1,
		output 		lvb_bb0_var__u2,
		input [31:0] 		workgroup_size
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb0_div_inputs_ready;
 reg local_bb0_div_wii_reg_NO_SHIFT_REG;
 reg local_bb0_div_valid_out_NO_SHIFT_REG;
wire local_bb0_div_stall_in;
wire local_bb0_div_output_regs_ready;
 reg [31:0] local_bb0_div_NO_SHIFT_REG;
wire local_bb0_div_causedstall;

assign local_bb0_div_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb0_div_output_regs_ready = (~(local_bb0_div_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_div_valid_out_NO_SHIFT_REG) | ~(local_bb0_div_stall_in))));
assign merge_node_stall_in_0 = (~(local_bb0_div_wii_reg_NO_SHIFT_REG) & (~(local_bb0_div_output_regs_ready) | ~(local_bb0_div_inputs_ready)));
assign local_bb0_div_causedstall = (local_bb0_div_inputs_ready && (~(local_bb0_div_output_regs_ready) && !(~(local_bb0_div_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_div_NO_SHIFT_REG <= 'x;
		local_bb0_div_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_div_NO_SHIFT_REG <= 'x;
			local_bb0_div_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_div_output_regs_ready)
			begin
				local_bb0_div_NO_SHIFT_REG <= (input_inSize_x >> 32'h1);
				local_bb0_div_valid_out_NO_SHIFT_REG <= local_bb0_div_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_div_stall_in))
				begin
					local_bb0_div_valid_out_NO_SHIFT_REG <= local_bb0_div_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_div_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_div_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_div_inputs_ready)
			begin
				local_bb0_div_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_div1_inputs_ready;
 reg local_bb0_div1_wii_reg_NO_SHIFT_REG;
 reg local_bb0_div1_valid_out_NO_SHIFT_REG;
wire local_bb0_div1_stall_in;
wire local_bb0_div1_output_regs_ready;
 reg [31:0] local_bb0_div1_NO_SHIFT_REG;
wire local_bb0_div1_causedstall;

assign local_bb0_div1_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb0_div1_output_regs_ready = (~(local_bb0_div1_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_div1_valid_out_NO_SHIFT_REG) | ~(local_bb0_div1_stall_in))));
assign merge_node_stall_in_1 = (~(local_bb0_div1_wii_reg_NO_SHIFT_REG) & (~(local_bb0_div1_output_regs_ready) | ~(local_bb0_div1_inputs_ready)));
assign local_bb0_div1_causedstall = (local_bb0_div1_inputs_ready && (~(local_bb0_div1_output_regs_ready) && !(~(local_bb0_div1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_div1_NO_SHIFT_REG <= 'x;
		local_bb0_div1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_div1_NO_SHIFT_REG <= 'x;
			local_bb0_div1_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_div1_output_regs_ready)
			begin
				local_bb0_div1_NO_SHIFT_REG <= (input_inSize_y >> 32'h1);
				local_bb0_div1_valid_out_NO_SHIFT_REG <= local_bb0_div1_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_div1_stall_in))
				begin
					local_bb0_div1_valid_out_NO_SHIFT_REG <= local_bb0_div1_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_div1_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_div1_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_div1_inputs_ready)
			begin
				local_bb0_div1_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_add7_inputs_ready;
 reg local_bb0_add7_wii_reg_NO_SHIFT_REG;
 reg local_bb0_add7_valid_out_NO_SHIFT_REG;
wire local_bb0_add7_stall_in;
wire local_bb0_add7_output_regs_ready;
 reg [31:0] local_bb0_add7_NO_SHIFT_REG;
wire local_bb0_add7_causedstall;

assign local_bb0_add7_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign local_bb0_add7_output_regs_ready = (~(local_bb0_add7_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_add7_valid_out_NO_SHIFT_REG) | ~(local_bb0_add7_stall_in))));
assign merge_node_stall_in_2 = (~(local_bb0_add7_wii_reg_NO_SHIFT_REG) & (~(local_bb0_add7_output_regs_ready) | ~(local_bb0_add7_inputs_ready)));
assign local_bb0_add7_causedstall = (local_bb0_add7_inputs_ready && (~(local_bb0_add7_output_regs_ready) && !(~(local_bb0_add7_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add7_NO_SHIFT_REG <= 'x;
		local_bb0_add7_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add7_NO_SHIFT_REG <= 'x;
			local_bb0_add7_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add7_output_regs_ready)
			begin
				local_bb0_add7_NO_SHIFT_REG <= (32'h1 - input_r);
				local_bb0_add7_valid_out_NO_SHIFT_REG <= local_bb0_add7_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_add7_stall_in))
				begin
					local_bb0_add7_valid_out_NO_SHIFT_REG <= local_bb0_add7_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add7_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add7_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add7_inputs_ready)
			begin
				local_bb0_add7_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub20_inputs_ready;
 reg local_bb0_sub20_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub20_valid_out_NO_SHIFT_REG;
wire local_bb0_sub20_stall_in;
wire local_bb0_sub20_output_regs_ready;
 reg [31:0] local_bb0_sub20_NO_SHIFT_REG;
wire local_bb0_sub20_causedstall;

assign local_bb0_sub20_inputs_ready = merge_node_valid_out_4_NO_SHIFT_REG;
assign local_bb0_sub20_output_regs_ready = (~(local_bb0_sub20_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_sub20_valid_out_NO_SHIFT_REG) | ~(local_bb0_sub20_stall_in))));
assign merge_node_stall_in_4 = (~(local_bb0_sub20_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub20_output_regs_ready) | ~(local_bb0_sub20_inputs_ready)));
assign local_bb0_sub20_causedstall = (local_bb0_sub20_inputs_ready && (~(local_bb0_sub20_output_regs_ready) && !(~(local_bb0_sub20_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub20_NO_SHIFT_REG <= 'x;
		local_bb0_sub20_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub20_NO_SHIFT_REG <= 'x;
			local_bb0_sub20_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub20_output_regs_ready)
			begin
				local_bb0_sub20_NO_SHIFT_REG <= (input_inSize_x + 32'hFFFFFFFF);
				local_bb0_sub20_valid_out_NO_SHIFT_REG <= local_bb0_sub20_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub20_stall_in))
				begin
					local_bb0_sub20_valid_out_NO_SHIFT_REG <= local_bb0_sub20_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub20_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub20_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub20_inputs_ready)
			begin
				local_bb0_sub20_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub22_inputs_ready;
 reg local_bb0_sub22_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub22_valid_out_NO_SHIFT_REG;
wire local_bb0_sub22_stall_in;
wire local_bb0_sub22_output_regs_ready;
 reg [31:0] local_bb0_sub22_NO_SHIFT_REG;
wire local_bb0_sub22_causedstall;

assign local_bb0_sub22_inputs_ready = merge_node_valid_out_5_NO_SHIFT_REG;
assign local_bb0_sub22_output_regs_ready = (~(local_bb0_sub22_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_sub22_valid_out_NO_SHIFT_REG) | ~(local_bb0_sub22_stall_in))));
assign merge_node_stall_in_5 = (~(local_bb0_sub22_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub22_output_regs_ready) | ~(local_bb0_sub22_inputs_ready)));
assign local_bb0_sub22_causedstall = (local_bb0_sub22_inputs_ready && (~(local_bb0_sub22_output_regs_ready) && !(~(local_bb0_sub22_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub22_NO_SHIFT_REG <= 'x;
		local_bb0_sub22_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub22_NO_SHIFT_REG <= 'x;
			local_bb0_sub22_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub22_output_regs_ready)
			begin
				local_bb0_sub22_NO_SHIFT_REG <= (input_inSize_y + 32'hFFFFFFFF);
				local_bb0_sub22_valid_out_NO_SHIFT_REG <= local_bb0_sub22_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub22_stall_in))
				begin
					local_bb0_sub22_valid_out_NO_SHIFT_REG <= local_bb0_sub22_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub22_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub22_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub22_inputs_ready)
			begin
				local_bb0_sub22_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_3to3_bb0_div_valid_out_0;
wire rstag_3to3_bb0_div_stall_in_0;
wire rstag_3to3_bb0_div_valid_out_1;
wire rstag_3to3_bb0_div_stall_in_1;
wire rstag_3to3_bb0_div_inputs_ready;
wire rstag_3to3_bb0_div_stall_local;
 reg rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG;
wire rstag_3to3_bb0_div_combined_valid;
 reg [31:0] rstag_3to3_bb0_div_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_3to3_bb0_div;
 reg rstag_3to3_bb0_div_consumed_0_NO_SHIFT_REG;
 reg rstag_3to3_bb0_div_consumed_1_NO_SHIFT_REG;

assign rstag_3to3_bb0_div_inputs_ready = local_bb0_div_valid_out_NO_SHIFT_REG;
assign rstag_3to3_bb0_div = (rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG ? rstag_3to3_bb0_div_staging_reg_NO_SHIFT_REG : (local_bb0_div_NO_SHIFT_REG & 32'h7FFFFFFF));
assign rstag_3to3_bb0_div_combined_valid = (rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG | rstag_3to3_bb0_div_inputs_ready);
assign rstag_3to3_bb0_div_stall_local = ((rstag_3to3_bb0_div_stall_in_0 & ~(rstag_3to3_bb0_div_consumed_0_NO_SHIFT_REG)) | (rstag_3to3_bb0_div_stall_in_1 & ~(rstag_3to3_bb0_div_consumed_1_NO_SHIFT_REG)));
assign rstag_3to3_bb0_div_valid_out_0 = (rstag_3to3_bb0_div_combined_valid & ~(rstag_3to3_bb0_div_consumed_0_NO_SHIFT_REG));
assign rstag_3to3_bb0_div_valid_out_1 = (rstag_3to3_bb0_div_combined_valid & ~(rstag_3to3_bb0_div_consumed_1_NO_SHIFT_REG));
assign local_bb0_div_stall_in = (|rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb0_div_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_3to3_bb0_div_stall_local)
			begin
				if (~(rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG))
				begin
					rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG <= rstag_3to3_bb0_div_inputs_ready;
				end
			end
			else
			begin
				rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_3to3_bb0_div_staging_valid_NO_SHIFT_REG))
		begin
			rstag_3to3_bb0_div_staging_reg_NO_SHIFT_REG <= (local_bb0_div_NO_SHIFT_REG & 32'h7FFFFFFF);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb0_div_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb0_div_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_3to3_bb0_div_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_3to3_bb0_div_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_3to3_bb0_div_consumed_0_NO_SHIFT_REG <= (rstag_3to3_bb0_div_combined_valid & (rstag_3to3_bb0_div_consumed_0_NO_SHIFT_REG | ~(rstag_3to3_bb0_div_stall_in_0)) & rstag_3to3_bb0_div_stall_local);
			rstag_3to3_bb0_div_consumed_1_NO_SHIFT_REG <= (rstag_3to3_bb0_div_combined_valid & (rstag_3to3_bb0_div_consumed_1_NO_SHIFT_REG | ~(rstag_3to3_bb0_div_stall_in_1)) & rstag_3to3_bb0_div_stall_local);
		end
	end
end


// This section implements a staging register.
// 
wire rstag_2to2_bb0_div1_valid_out_0;
wire rstag_2to2_bb0_div1_stall_in_0;
wire rstag_2to2_bb0_div1_valid_out_1;
wire rstag_2to2_bb0_div1_stall_in_1;
wire rstag_2to2_bb0_div1_inputs_ready;
wire rstag_2to2_bb0_div1_stall_local;
 reg rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG;
wire rstag_2to2_bb0_div1_combined_valid;
 reg [31:0] rstag_2to2_bb0_div1_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_2to2_bb0_div1;
 reg rstag_2to2_bb0_div1_consumed_0_NO_SHIFT_REG;
 reg rstag_2to2_bb0_div1_consumed_1_NO_SHIFT_REG;

assign rstag_2to2_bb0_div1_inputs_ready = local_bb0_div1_valid_out_NO_SHIFT_REG;
assign rstag_2to2_bb0_div1 = (rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG ? rstag_2to2_bb0_div1_staging_reg_NO_SHIFT_REG : (local_bb0_div1_NO_SHIFT_REG & 32'h7FFFFFFF));
assign rstag_2to2_bb0_div1_combined_valid = (rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG | rstag_2to2_bb0_div1_inputs_ready);
assign rstag_2to2_bb0_div1_stall_local = ((rstag_2to2_bb0_div1_stall_in_0 & ~(rstag_2to2_bb0_div1_consumed_0_NO_SHIFT_REG)) | (rstag_2to2_bb0_div1_stall_in_1 & ~(rstag_2to2_bb0_div1_consumed_1_NO_SHIFT_REG)));
assign rstag_2to2_bb0_div1_valid_out_0 = (rstag_2to2_bb0_div1_combined_valid & ~(rstag_2to2_bb0_div1_consumed_0_NO_SHIFT_REG));
assign rstag_2to2_bb0_div1_valid_out_1 = (rstag_2to2_bb0_div1_combined_valid & ~(rstag_2to2_bb0_div1_consumed_1_NO_SHIFT_REG));
assign local_bb0_div1_stall_in = (|rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_div1_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_2to2_bb0_div1_stall_local)
			begin
				if (~(rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG))
				begin
					rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG <= rstag_2to2_bb0_div1_inputs_ready;
				end
			end
			else
			begin
				rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_2to2_bb0_div1_staging_valid_NO_SHIFT_REG))
		begin
			rstag_2to2_bb0_div1_staging_reg_NO_SHIFT_REG <= (local_bb0_div1_NO_SHIFT_REG & 32'h7FFFFFFF);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_div1_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_div1_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_div1_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_2to2_bb0_div1_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_2to2_bb0_div1_consumed_0_NO_SHIFT_REG <= (rstag_2to2_bb0_div1_combined_valid & (rstag_2to2_bb0_div1_consumed_0_NO_SHIFT_REG | ~(rstag_2to2_bb0_div1_stall_in_0)) & rstag_2to2_bb0_div1_stall_local);
			rstag_2to2_bb0_div1_consumed_1_NO_SHIFT_REG <= (rstag_2to2_bb0_div1_combined_valid & (rstag_2to2_bb0_div1_consumed_1_NO_SHIFT_REG | ~(rstag_2to2_bb0_div1_stall_in_1)) & rstag_2to2_bb0_div1_stall_local);
		end
	end
end


// This section implements a staging register.
// 
wire rstag_3to3_bb0_add7_valid_out_0;
wire rstag_3to3_bb0_add7_stall_in_0;
wire rstag_3to3_bb0_add7_valid_out_1;
wire rstag_3to3_bb0_add7_stall_in_1;
wire rstag_3to3_bb0_add7_inputs_ready;
wire rstag_3to3_bb0_add7_stall_local;
 reg rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG;
wire rstag_3to3_bb0_add7_combined_valid;
 reg [31:0] rstag_3to3_bb0_add7_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_3to3_bb0_add7;
 reg rstag_3to3_bb0_add7_consumed_0_NO_SHIFT_REG;
 reg rstag_3to3_bb0_add7_consumed_1_NO_SHIFT_REG;

assign rstag_3to3_bb0_add7_inputs_ready = local_bb0_add7_valid_out_NO_SHIFT_REG;
assign rstag_3to3_bb0_add7 = (rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG ? rstag_3to3_bb0_add7_staging_reg_NO_SHIFT_REG : local_bb0_add7_NO_SHIFT_REG);
assign rstag_3to3_bb0_add7_combined_valid = (rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG | rstag_3to3_bb0_add7_inputs_ready);
assign rstag_3to3_bb0_add7_stall_local = ((rstag_3to3_bb0_add7_stall_in_0 & ~(rstag_3to3_bb0_add7_consumed_0_NO_SHIFT_REG)) | (rstag_3to3_bb0_add7_stall_in_1 & ~(rstag_3to3_bb0_add7_consumed_1_NO_SHIFT_REG)));
assign rstag_3to3_bb0_add7_valid_out_0 = (rstag_3to3_bb0_add7_combined_valid & ~(rstag_3to3_bb0_add7_consumed_0_NO_SHIFT_REG));
assign rstag_3to3_bb0_add7_valid_out_1 = (rstag_3to3_bb0_add7_combined_valid & ~(rstag_3to3_bb0_add7_consumed_1_NO_SHIFT_REG));
assign local_bb0_add7_stall_in = (|rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb0_add7_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_3to3_bb0_add7_stall_local)
			begin
				if (~(rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG))
				begin
					rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG <= rstag_3to3_bb0_add7_inputs_ready;
				end
			end
			else
			begin
				rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_3to3_bb0_add7_staging_valid_NO_SHIFT_REG))
		begin
			rstag_3to3_bb0_add7_staging_reg_NO_SHIFT_REG <= local_bb0_add7_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb0_add7_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb0_add7_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_3to3_bb0_add7_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_3to3_bb0_add7_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_3to3_bb0_add7_consumed_0_NO_SHIFT_REG <= (rstag_3to3_bb0_add7_combined_valid & (rstag_3to3_bb0_add7_consumed_0_NO_SHIFT_REG | ~(rstag_3to3_bb0_add7_stall_in_0)) & rstag_3to3_bb0_add7_stall_local);
			rstag_3to3_bb0_add7_consumed_1_NO_SHIFT_REG <= (rstag_3to3_bb0_add7_combined_valid & (rstag_3to3_bb0_add7_consumed_1_NO_SHIFT_REG | ~(rstag_3to3_bb0_add7_stall_in_1)) & rstag_3to3_bb0_add7_stall_local);
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_cmp315_valid_out;
wire local_bb0_cmp315_stall_in;
wire local_bb0_cmp315_inputs_ready;
wire local_bb0_cmp315_stall_local;
wire local_bb0_cmp315;

assign local_bb0_cmp315_inputs_ready = rstag_3to3_bb0_div_valid_out_1;
assign local_bb0_cmp315 = ((rstag_3to3_bb0_div & 32'h7FFFFFFF) == 32'h0);
assign local_bb0_cmp315_valid_out = local_bb0_cmp315_inputs_ready;
assign local_bb0_cmp315_stall_local = local_bb0_cmp315_stall_in;
assign rstag_3to3_bb0_div_stall_in_1 = (|local_bb0_cmp315_stall_local);

// This section implements a registered operation.
// 
wire local_bb0_cmp19_inputs_ready;
 reg local_bb0_cmp19_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp19_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp19_stall_in;
wire local_bb0_cmp19_output_regs_ready;
 reg local_bb0_cmp19_NO_SHIFT_REG;
wire local_bb0_cmp19_causedstall;

assign local_bb0_cmp19_inputs_ready = rstag_2to2_bb0_div1_valid_out_1;
assign local_bb0_cmp19_output_regs_ready = (~(local_bb0_cmp19_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp19_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp19_stall_in))));
assign rstag_2to2_bb0_div1_stall_in_1 = (~(local_bb0_cmp19_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp19_output_regs_ready) | ~(local_bb0_cmp19_inputs_ready)));
assign local_bb0_cmp19_causedstall = (local_bb0_cmp19_inputs_ready && (~(local_bb0_cmp19_output_regs_ready) && !(~(local_bb0_cmp19_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp19_NO_SHIFT_REG <= 'x;
		local_bb0_cmp19_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp19_NO_SHIFT_REG <= 'x;
			local_bb0_cmp19_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp19_output_regs_ready)
			begin
				local_bb0_cmp19_NO_SHIFT_REG <= ((rstag_2to2_bb0_div1 & 32'h7FFFFFFF) == 32'h0);
				local_bb0_cmp19_valid_out_NO_SHIFT_REG <= local_bb0_cmp19_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp19_stall_in))
				begin
					local_bb0_cmp19_valid_out_NO_SHIFT_REG <= local_bb0_cmp19_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp19_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp19_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp19_inputs_ready)
			begin
				local_bb0_cmp19_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp98_inputs_ready;
 reg local_bb0_cmp98_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp98_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp98_stall_in;
wire local_bb0_cmp98_output_regs_ready;
 reg local_bb0_cmp98_NO_SHIFT_REG;
wire local_bb0_cmp98_causedstall;

assign local_bb0_cmp98_inputs_ready = (merge_node_valid_out_3_NO_SHIFT_REG & rstag_3to3_bb0_add7_valid_out_1);
assign local_bb0_cmp98_output_regs_ready = (~(local_bb0_cmp98_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp98_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp98_stall_in))));
assign merge_node_stall_in_3 = (~(local_bb0_cmp98_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp98_output_regs_ready) | ~(local_bb0_cmp98_inputs_ready)));
assign rstag_3to3_bb0_add7_stall_in_1 = (~(local_bb0_cmp98_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp98_output_regs_ready) | ~(local_bb0_cmp98_inputs_ready)));
assign local_bb0_cmp98_causedstall = (local_bb0_cmp98_inputs_ready && (~(local_bb0_cmp98_output_regs_ready) && !(~(local_bb0_cmp98_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp98_NO_SHIFT_REG <= 'x;
		local_bb0_cmp98_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp98_NO_SHIFT_REG <= 'x;
			local_bb0_cmp98_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp98_output_regs_ready)
			begin
				local_bb0_cmp98_NO_SHIFT_REG <= ($signed(rstag_3to3_bb0_add7) > $signed(input_r));
				local_bb0_cmp98_valid_out_NO_SHIFT_REG <= local_bb0_cmp98_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp98_stall_in))
				begin
					local_bb0_cmp98_valid_out_NO_SHIFT_REG <= local_bb0_cmp98_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp98_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp98_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp98_inputs_ready)
			begin
				local_bb0_cmp98_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_3to3_bb0_cmp19_valid_out_0;
wire rstag_3to3_bb0_cmp19_stall_in_0;
wire rstag_3to3_bb0_cmp19_valid_out_1;
wire rstag_3to3_bb0_cmp19_stall_in_1;
wire rstag_3to3_bb0_cmp19_valid_out_2;
wire rstag_3to3_bb0_cmp19_stall_in_2;
wire rstag_3to3_bb0_cmp19_inputs_ready;
wire rstag_3to3_bb0_cmp19_stall_local;
 reg rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG;
wire rstag_3to3_bb0_cmp19_combined_valid;
 reg rstag_3to3_bb0_cmp19_staging_reg_NO_SHIFT_REG;
wire rstag_3to3_bb0_cmp19;
 reg rstag_3to3_bb0_cmp19_consumed_0_NO_SHIFT_REG;
 reg rstag_3to3_bb0_cmp19_consumed_1_NO_SHIFT_REG;
 reg rstag_3to3_bb0_cmp19_consumed_2_NO_SHIFT_REG;

assign rstag_3to3_bb0_cmp19_inputs_ready = local_bb0_cmp19_valid_out_NO_SHIFT_REG;
assign rstag_3to3_bb0_cmp19 = (rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG ? rstag_3to3_bb0_cmp19_staging_reg_NO_SHIFT_REG : local_bb0_cmp19_NO_SHIFT_REG);
assign rstag_3to3_bb0_cmp19_combined_valid = (rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG | rstag_3to3_bb0_cmp19_inputs_ready);
assign rstag_3to3_bb0_cmp19_stall_local = ((rstag_3to3_bb0_cmp19_stall_in_0 & ~(rstag_3to3_bb0_cmp19_consumed_0_NO_SHIFT_REG)) | (rstag_3to3_bb0_cmp19_stall_in_1 & ~(rstag_3to3_bb0_cmp19_consumed_1_NO_SHIFT_REG)) | (rstag_3to3_bb0_cmp19_stall_in_2 & ~(rstag_3to3_bb0_cmp19_consumed_2_NO_SHIFT_REG)));
assign rstag_3to3_bb0_cmp19_valid_out_0 = (rstag_3to3_bb0_cmp19_combined_valid & ~(rstag_3to3_bb0_cmp19_consumed_0_NO_SHIFT_REG));
assign rstag_3to3_bb0_cmp19_valid_out_1 = (rstag_3to3_bb0_cmp19_combined_valid & ~(rstag_3to3_bb0_cmp19_consumed_1_NO_SHIFT_REG));
assign rstag_3to3_bb0_cmp19_valid_out_2 = (rstag_3to3_bb0_cmp19_combined_valid & ~(rstag_3to3_bb0_cmp19_consumed_2_NO_SHIFT_REG));
assign local_bb0_cmp19_stall_in = (|rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb0_cmp19_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_3to3_bb0_cmp19_stall_local)
			begin
				if (~(rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG))
				begin
					rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG <= rstag_3to3_bb0_cmp19_inputs_ready;
				end
			end
			else
			begin
				rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_3to3_bb0_cmp19_staging_valid_NO_SHIFT_REG))
		begin
			rstag_3to3_bb0_cmp19_staging_reg_NO_SHIFT_REG <= local_bb0_cmp19_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb0_cmp19_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb0_cmp19_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb0_cmp19_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_3to3_bb0_cmp19_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_3to3_bb0_cmp19_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_3to3_bb0_cmp19_consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_3to3_bb0_cmp19_consumed_0_NO_SHIFT_REG <= (rstag_3to3_bb0_cmp19_combined_valid & (rstag_3to3_bb0_cmp19_consumed_0_NO_SHIFT_REG | ~(rstag_3to3_bb0_cmp19_stall_in_0)) & rstag_3to3_bb0_cmp19_stall_local);
			rstag_3to3_bb0_cmp19_consumed_1_NO_SHIFT_REG <= (rstag_3to3_bb0_cmp19_combined_valid & (rstag_3to3_bb0_cmp19_consumed_1_NO_SHIFT_REG | ~(rstag_3to3_bb0_cmp19_stall_in_1)) & rstag_3to3_bb0_cmp19_stall_local);
			rstag_3to3_bb0_cmp19_consumed_2_NO_SHIFT_REG <= (rstag_3to3_bb0_cmp19_combined_valid & (rstag_3to3_bb0_cmp19_consumed_2_NO_SHIFT_REG | ~(rstag_3to3_bb0_cmp19_stall_in_2)) & rstag_3to3_bb0_cmp19_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u2_inputs_ready;
 reg local_bb0_var__u2_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u2_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u2_stall_in;
wire local_bb0_var__u2_output_regs_ready;
 reg local_bb0_var__u2_NO_SHIFT_REG;
wire local_bb0_var__u2_causedstall;

assign local_bb0_var__u2_inputs_ready = rstag_3to3_bb0_cmp19_valid_out_1;
assign local_bb0_var__u2_output_regs_ready = (~(local_bb0_var__u2_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u2_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u2_stall_in))));
assign rstag_3to3_bb0_cmp19_stall_in_1 = (~(local_bb0_var__u2_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u2_output_regs_ready) | ~(local_bb0_var__u2_inputs_ready)));
assign local_bb0_var__u2_causedstall = (local_bb0_var__u2_inputs_ready && (~(local_bb0_var__u2_output_regs_ready) && !(~(local_bb0_var__u2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u2_NO_SHIFT_REG <= 'x;
		local_bb0_var__u2_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u2_NO_SHIFT_REG <= 'x;
			local_bb0_var__u2_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u2_output_regs_ready)
			begin
				local_bb0_var__u2_NO_SHIFT_REG <= (rstag_3to3_bb0_cmp19 ^ 1'b1);
				local_bb0_var__u2_valid_out_NO_SHIFT_REG <= local_bb0_var__u2_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u2_stall_in))
				begin
					local_bb0_var__u2_valid_out_NO_SHIFT_REG <= local_bb0_var__u2_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u2_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u2_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u2_inputs_ready)
			begin
				local_bb0_var__u2_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__inputs_ready;
 reg local_bb0_var__wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__valid_out_NO_SHIFT_REG;
wire local_bb0_var__stall_in;
wire local_bb0_var__output_regs_ready;
 reg local_bb0_var__NO_SHIFT_REG;
wire local_bb0_var__causedstall;

assign local_bb0_var__inputs_ready = (local_bb0_cmp315_valid_out & rstag_3to3_bb0_cmp19_valid_out_2);
assign local_bb0_var__output_regs_ready = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__valid_out_NO_SHIFT_REG) | ~(local_bb0_var__stall_in))));
assign local_bb0_cmp315_stall_in = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__output_regs_ready) | ~(local_bb0_var__inputs_ready)));
assign rstag_3to3_bb0_cmp19_stall_in_2 = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__output_regs_ready) | ~(local_bb0_var__inputs_ready)));
assign local_bb0_var__causedstall = (local_bb0_var__inputs_ready && (~(local_bb0_var__output_regs_ready) && !(~(local_bb0_var__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__NO_SHIFT_REG <= 'x;
		local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__NO_SHIFT_REG <= 'x;
			local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__output_regs_ready)
			begin
				local_bb0_var__NO_SHIFT_REG <= (rstag_3to3_bb0_cmp19 | local_bb0_cmp315);
				local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__stall_in))
				begin
					local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__inputs_ready)
			begin
				local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_4to4_bb0_var__valid_out_0;
wire rstag_4to4_bb0_var__stall_in_0;
wire rstag_4to4_bb0_var__valid_out_1;
wire rstag_4to4_bb0_var__stall_in_1;
wire rstag_4to4_bb0_var__valid_out_2;
wire rstag_4to4_bb0_var__stall_in_2;
wire rstag_4to4_bb0_var__inputs_ready;
wire rstag_4to4_bb0_var__stall_local;
 reg rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG;
wire rstag_4to4_bb0_var__combined_valid;
 reg rstag_4to4_bb0_var__staging_reg_NO_SHIFT_REG;
wire rstag_4to4_bb0_var_;
 reg rstag_4to4_bb0_var__consumed_0_NO_SHIFT_REG;
 reg rstag_4to4_bb0_var__consumed_1_NO_SHIFT_REG;
 reg rstag_4to4_bb0_var__consumed_2_NO_SHIFT_REG;

assign rstag_4to4_bb0_var__inputs_ready = local_bb0_var__valid_out_NO_SHIFT_REG;
assign rstag_4to4_bb0_var_ = (rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG ? rstag_4to4_bb0_var__staging_reg_NO_SHIFT_REG : local_bb0_var__NO_SHIFT_REG);
assign rstag_4to4_bb0_var__combined_valid = (rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG | rstag_4to4_bb0_var__inputs_ready);
assign rstag_4to4_bb0_var__stall_local = ((rstag_4to4_bb0_var__stall_in_0 & ~(rstag_4to4_bb0_var__consumed_0_NO_SHIFT_REG)) | (rstag_4to4_bb0_var__stall_in_1 & ~(rstag_4to4_bb0_var__consumed_1_NO_SHIFT_REG)) | (rstag_4to4_bb0_var__stall_in_2 & ~(rstag_4to4_bb0_var__consumed_2_NO_SHIFT_REG)));
assign rstag_4to4_bb0_var__valid_out_0 = (rstag_4to4_bb0_var__combined_valid & ~(rstag_4to4_bb0_var__consumed_0_NO_SHIFT_REG));
assign rstag_4to4_bb0_var__valid_out_1 = (rstag_4to4_bb0_var__combined_valid & ~(rstag_4to4_bb0_var__consumed_1_NO_SHIFT_REG));
assign rstag_4to4_bb0_var__valid_out_2 = (rstag_4to4_bb0_var__combined_valid & ~(rstag_4to4_bb0_var__consumed_2_NO_SHIFT_REG));
assign local_bb0_var__stall_in = (|rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_var__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_4to4_bb0_var__stall_local)
			begin
				if (~(rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG))
				begin
					rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG <= rstag_4to4_bb0_var__inputs_ready;
				end
			end
			else
			begin
				rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_4to4_bb0_var__staging_valid_NO_SHIFT_REG))
		begin
			rstag_4to4_bb0_var__staging_reg_NO_SHIFT_REG <= local_bb0_var__NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_var__consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_var__consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_var__consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_var__consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_var__consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_var__consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_4to4_bb0_var__consumed_0_NO_SHIFT_REG <= (rstag_4to4_bb0_var__combined_valid & (rstag_4to4_bb0_var__consumed_0_NO_SHIFT_REG | ~(rstag_4to4_bb0_var__stall_in_0)) & rstag_4to4_bb0_var__stall_local);
			rstag_4to4_bb0_var__consumed_1_NO_SHIFT_REG <= (rstag_4to4_bb0_var__combined_valid & (rstag_4to4_bb0_var__consumed_1_NO_SHIFT_REG | ~(rstag_4to4_bb0_var__stall_in_1)) & rstag_4to4_bb0_var__stall_local);
			rstag_4to4_bb0_var__consumed_2_NO_SHIFT_REG <= (rstag_4to4_bb0_var__combined_valid & (rstag_4to4_bb0_var__consumed_2_NO_SHIFT_REG | ~(rstag_4to4_bb0_var__stall_in_2)) & rstag_4to4_bb0_var__stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u1_inputs_ready;
 reg local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u1_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u1_stall_in;
wire local_bb0_var__u1_output_regs_ready;
 reg local_bb0_var__u1_NO_SHIFT_REG;
wire local_bb0_var__u1_causedstall;

assign local_bb0_var__u1_inputs_ready = rstag_4to4_bb0_var__valid_out_1;
assign local_bb0_var__u1_output_regs_ready = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u1_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u1_stall_in))));
assign rstag_4to4_bb0_var__stall_in_1 = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u1_output_regs_ready) | ~(local_bb0_var__u1_inputs_ready)));
assign local_bb0_var__u1_causedstall = (local_bb0_var__u1_inputs_ready && (~(local_bb0_var__u1_output_regs_ready) && !(~(local_bb0_var__u1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_NO_SHIFT_REG <= 'x;
		local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_NO_SHIFT_REG <= 'x;
			local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_output_regs_ready)
			begin
				local_bb0_var__u1_NO_SHIFT_REG <= (rstag_4to4_bb0_var_ ^ 1'b1);
				local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u1_stall_in))
				begin
					local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_inputs_ready)
			begin
				local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u0_inputs_ready;
 reg local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u0_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u0_stall_in;
wire local_bb0_var__u0_output_regs_ready;
 reg local_bb0_var__u0_NO_SHIFT_REG;
wire local_bb0_var__u0_causedstall;

assign local_bb0_var__u0_inputs_ready = (local_bb0_cmp98_valid_out_NO_SHIFT_REG & rstag_4to4_bb0_var__valid_out_2);
assign local_bb0_var__u0_output_regs_ready = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u0_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u0_stall_in))));
assign local_bb0_cmp98_stall_in = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u0_output_regs_ready) | ~(local_bb0_var__u0_inputs_ready)));
assign rstag_4to4_bb0_var__stall_in_2 = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u0_output_regs_ready) | ~(local_bb0_var__u0_inputs_ready)));
assign local_bb0_var__u0_causedstall = (local_bb0_var__u0_inputs_ready && (~(local_bb0_var__u0_output_regs_ready) && !(~(local_bb0_var__u0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_NO_SHIFT_REG <= 'x;
		local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_NO_SHIFT_REG <= 'x;
			local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_output_regs_ready)
			begin
				local_bb0_var__u0_NO_SHIFT_REG <= (rstag_4to4_bb0_var_ | local_bb0_cmp98_NO_SHIFT_REG);
				local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u0_stall_in))
				begin
					local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_inputs_ready)
			begin
				local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [31:0] lvb_bb0_div_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_div1_reg_NO_SHIFT_REG;
 reg lvb_bb0_cmp19_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_add7_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_sub20_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_sub22_reg_NO_SHIFT_REG;
 reg lvb_bb0_var__reg_NO_SHIFT_REG;
 reg lvb_bb0_var__u0_reg_NO_SHIFT_REG;
 reg lvb_bb0_var__u1_reg_NO_SHIFT_REG;
 reg lvb_bb0_var__u2_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb0_var__u2_valid_out_NO_SHIFT_REG & local_bb0_var__u1_valid_out_NO_SHIFT_REG & local_bb0_var__u0_valid_out_NO_SHIFT_REG & local_bb0_sub22_valid_out_NO_SHIFT_REG & local_bb0_sub20_valid_out_NO_SHIFT_REG & merge_node_valid_out_6_NO_SHIFT_REG & rstag_4to4_bb0_var__valid_out_0 & rstag_3to3_bb0_cmp19_valid_out_0 & rstag_3to3_bb0_add7_valid_out_0 & rstag_2to2_bb0_div1_valid_out_0 & rstag_3to3_bb0_div_valid_out_0);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb0_var__u2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_var__u1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_var__u0_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_sub22_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_sub20_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign merge_node_stall_in_6 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_4to4_bb0_var__stall_in_0 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_3to3_bb0_cmp19_stall_in_0 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_3to3_bb0_add7_stall_in_0 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_2to2_bb0_div1_stall_in_0 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_3to3_bb0_div_stall_in_0 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb0_div = lvb_bb0_div_reg_NO_SHIFT_REG;
assign lvb_bb0_div1 = lvb_bb0_div1_reg_NO_SHIFT_REG;
assign lvb_bb0_cmp19 = lvb_bb0_cmp19_reg_NO_SHIFT_REG;
assign lvb_bb0_add7 = lvb_bb0_add7_reg_NO_SHIFT_REG;
assign lvb_bb0_sub20 = lvb_bb0_sub20_reg_NO_SHIFT_REG;
assign lvb_bb0_sub22 = lvb_bb0_sub22_reg_NO_SHIFT_REG;
assign lvb_bb0_var_ = lvb_bb0_var__reg_NO_SHIFT_REG;
assign lvb_bb0_var__u0 = lvb_bb0_var__u0_reg_NO_SHIFT_REG;
assign lvb_bb0_var__u1 = lvb_bb0_var__u1_reg_NO_SHIFT_REG;
assign lvb_bb0_var__u2 = lvb_bb0_var__u2_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb0_div_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_div1_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_cmp19_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_add7_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_sub20_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_sub22_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__u0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__u1_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__u2_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb0_div_reg_NO_SHIFT_REG <= (rstag_3to3_bb0_div & 32'h7FFFFFFF);
			lvb_bb0_div1_reg_NO_SHIFT_REG <= (rstag_2to2_bb0_div1 & 32'h7FFFFFFF);
			lvb_bb0_cmp19_reg_NO_SHIFT_REG <= rstag_3to3_bb0_cmp19;
			lvb_bb0_add7_reg_NO_SHIFT_REG <= rstag_3to3_bb0_add7;
			lvb_bb0_sub20_reg_NO_SHIFT_REG <= local_bb0_sub20_NO_SHIFT_REG;
			lvb_bb0_sub22_reg_NO_SHIFT_REG <= local_bb0_sub22_NO_SHIFT_REG;
			lvb_bb0_var__reg_NO_SHIFT_REG <= rstag_4to4_bb0_var_;
			lvb_bb0_var__u0_reg_NO_SHIFT_REG <= local_bb0_var__u0_NO_SHIFT_REG;
			lvb_bb0_var__u1_reg_NO_SHIFT_REG <= local_bb0_var__u1_NO_SHIFT_REG;
			lvb_bb0_var__u2_reg_NO_SHIFT_REG <= local_bb0_var__u2_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_1
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_wii_div,
		input [31:0] 		input_wii_div1,
		input 		input_wii_cmp19,
		input [31:0] 		input_wii_add7,
		input [31:0] 		input_wii_sub20,
		input [31:0] 		input_wii_sub22,
		input 		input_wii_var_,
		input 		input_wii_var__u3,
		input 		input_wii_var__u4,
		input 		input_wii_var__u5,
		input 		valid_in_0,
		output 		stall_out_0,
		input 		input_forked17_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input 		input_forked17_1,
		output 		valid_out,
		input 		stall_in,
		output [31:0] 		lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0,
		output [31:0] 		lvb_bb1_mul37,
		output 		lvb_bb1_notcmp11,
		output 		lvb_bb1_notexitcond14_,
		output 		lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		feedback_valid_in_8,
		output 		feedback_stall_out_8,
		input [31:0] 		feedback_data_in_8,
		input 		feedback_valid_in_9,
		output 		feedback_stall_out_9,
		input 		feedback_data_in_9,
		output 		feedback_stall_out_6,
		input 		feedback_valid_in_7,
		output 		feedback_stall_out_7,
		input 		feedback_data_in_7,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		output 		feedback_valid_out_8,
		input 		feedback_stall_in_8,
		output [31:0] 		feedback_data_out_8,
		output 		feedback_valid_out_7,
		input 		feedback_stall_in_7,
		output 		feedback_data_out_7
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg input_forked17_0_staging_reg_NO_SHIFT_REG;
 reg local_lvm_forked17_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg input_forked17_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_forked17_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_forked17_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_forked17_0_staging_reg_NO_SHIFT_REG <= input_forked17_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_forked17_1_staging_reg_NO_SHIFT_REG <= input_forked17_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_local;
wire [31:0] local_bb1_pixel_y_020_pop8_acl_pop_i32_0;
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_fu_valid_out;
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_fu_stall_out;
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_inputs_ready;

acl_pop local_bb1_pixel_y_020_pop8_acl_pop_i32_0_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_forked17_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(32'h0),
	.stall_out(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_fu_stall_out),
	.valid_in(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_inputs_ready),
	.valid_out(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_fu_valid_out),
	.stall_in(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_local),
	.data_out(local_bb1_pixel_y_020_pop8_acl_pop_i32_0),
	.feedback_in(feedback_data_in_8),
	.feedback_valid_in(feedback_valid_in_8),
	.feedback_stall_out(feedback_stall_out_8)
);

defparam local_bb1_pixel_y_020_pop8_acl_pop_i32_0_feedback.COALESCE_DISTANCE = 1;
defparam local_bb1_pixel_y_020_pop8_acl_pop_i32_0_feedback.DATA_WIDTH = 32;
defparam local_bb1_pixel_y_020_pop8_acl_pop_i32_0_feedback.STYLE = "REGULAR";


// This section implements a registered operation.
// 
wire local_bb1_memdep_phi1_pop9_acl_pop_i1_0_inputs_ready;
 reg local_bb1_memdep_phi1_pop9_acl_pop_i1_0_valid_out_NO_SHIFT_REG;
wire local_bb1_memdep_phi1_pop9_acl_pop_i1_0_stall_in;
wire local_bb1_memdep_phi1_pop9_acl_pop_i1_0_output_regs_ready;
wire local_bb1_memdep_phi1_pop9_acl_pop_i1_0_result;
wire local_bb1_memdep_phi1_pop9_acl_pop_i1_0_fu_valid_out;
wire local_bb1_memdep_phi1_pop9_acl_pop_i1_0_fu_stall_out;
 reg local_bb1_memdep_phi1_pop9_acl_pop_i1_0_NO_SHIFT_REG;
wire local_bb1_memdep_phi1_pop9_acl_pop_i1_0_causedstall;

acl_pop local_bb1_memdep_phi1_pop9_acl_pop_i1_0_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_forked17_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(1'b0),
	.stall_out(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_fu_stall_out),
	.valid_in(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_inputs_ready),
	.valid_out(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_fu_valid_out),
	.stall_in(~(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_output_regs_ready)),
	.data_out(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_result),
	.feedback_in(feedback_data_in_9),
	.feedback_valid_in(feedback_valid_in_9),
	.feedback_stall_out(feedback_stall_out_9)
);

defparam local_bb1_memdep_phi1_pop9_acl_pop_i1_0_feedback.COALESCE_DISTANCE = 1;
defparam local_bb1_memdep_phi1_pop9_acl_pop_i1_0_feedback.DATA_WIDTH = 1;
defparam local_bb1_memdep_phi1_pop9_acl_pop_i1_0_feedback.STYLE = "REGULAR";

assign local_bb1_memdep_phi1_pop9_acl_pop_i1_0_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb1_memdep_phi1_pop9_acl_pop_i1_0_output_regs_ready = (&(~(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_valid_out_NO_SHIFT_REG) | ~(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_stall_in)));
assign merge_node_stall_in_1 = (local_bb1_memdep_phi1_pop9_acl_pop_i1_0_fu_stall_out | ~(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_inputs_ready));
assign local_bb1_memdep_phi1_pop9_acl_pop_i1_0_causedstall = (local_bb1_memdep_phi1_pop9_acl_pop_i1_0_inputs_ready && (local_bb1_memdep_phi1_pop9_acl_pop_i1_0_fu_stall_out && !(~(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_memdep_phi1_pop9_acl_pop_i1_0_NO_SHIFT_REG <= 'x;
		local_bb1_memdep_phi1_pop9_acl_pop_i1_0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_memdep_phi1_pop9_acl_pop_i1_0_output_regs_ready)
		begin
			local_bb1_memdep_phi1_pop9_acl_pop_i1_0_NO_SHIFT_REG <= local_bb1_memdep_phi1_pop9_acl_pop_i1_0_result;
			local_bb1_memdep_phi1_pop9_acl_pop_i1_0_valid_out_NO_SHIFT_REG <= local_bb1_memdep_phi1_pop9_acl_pop_i1_0_fu_valid_out;
		end
		else
		begin
			if (~(local_bb1_memdep_phi1_pop9_acl_pop_i1_0_stall_in))
			begin
				local_bb1_memdep_phi1_pop9_acl_pop_i1_0_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_fifo.DATA_WIDTH = 0;
defparam rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_reg_2_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign merge_node_stall_in_2 = rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_valid_out_reg_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb1_inc45_stall_local;
wire [31:0] local_bb1_inc45;

assign local_bb1_inc45 = (local_bb1_pixel_y_020_pop8_acl_pop_i32_0 + 32'h1);

// This section implements a registered operation.
// 
wire local_bb1_keep_going13_acl_pipeline_1_inputs_ready;
 reg local_bb1_keep_going13_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb1_keep_going13_acl_pipeline_1_stall_in;
wire local_bb1_keep_going13_acl_pipeline_1_output_regs_ready;
wire local_bb1_keep_going13_acl_pipeline_1_keep_going;
wire local_bb1_keep_going13_acl_pipeline_1_fu_valid_out;
wire local_bb1_keep_going13_acl_pipeline_1_fu_stall_out;
 reg local_bb1_keep_going13_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb1_keep_going13_acl_pipeline_1_feedback_pipelined;
wire local_bb1_keep_going13_acl_pipeline_1_causedstall;

acl_pipeline local_bb1_keep_going13_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb1_keep_going13_acl_pipeline_1_fu_stall_out),
	.valid_in(local_bb1_keep_going13_acl_pipeline_1_inputs_ready),
	.valid_out(local_bb1_keep_going13_acl_pipeline_1_fu_valid_out),
	.stall_in(~(local_bb1_keep_going13_acl_pipeline_1_output_regs_ready)),
	.data_out(local_bb1_keep_going13_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_6),
	.not_exitcond_in(feedback_data_in_7),
	.not_exitcond_valid_in(feedback_valid_in_7),
	.not_exitcond_stall_out(feedback_stall_out_7),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb1_keep_going13_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb1_keep_going13_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb1_keep_going13_acl_pipeline_1_inputs_ready = rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
assign local_bb1_keep_going13_acl_pipeline_1_output_regs_ready = (&(~(local_bb1_keep_going13_acl_pipeline_1_valid_out_NO_SHIFT_REG) | ~(local_bb1_keep_going13_acl_pipeline_1_stall_in)));
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign rnode_1to2_bb1_keep_going13_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = (local_bb1_keep_going13_acl_pipeline_1_fu_stall_out | ~(local_bb1_keep_going13_acl_pipeline_1_inputs_ready));
assign local_bb1_keep_going13_acl_pipeline_1_causedstall = (local_bb1_keep_going13_acl_pipeline_1_inputs_ready && (local_bb1_keep_going13_acl_pipeline_1_fu_stall_out && !(~(local_bb1_keep_going13_acl_pipeline_1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_keep_going13_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb1_keep_going13_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_keep_going13_acl_pipeline_1_output_regs_ready)
		begin
			local_bb1_keep_going13_acl_pipeline_1_NO_SHIFT_REG <= local_bb1_keep_going13_acl_pipeline_1_keep_going;
			local_bb1_keep_going13_acl_pipeline_1_valid_out_NO_SHIFT_REG <= local_bb1_keep_going13_acl_pipeline_1_fu_valid_out;
		end
		else
		begin
			if (~(local_bb1_keep_going13_acl_pipeline_1_stall_in))
			begin
				local_bb1_keep_going13_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1_cmp_stall_local;
wire [32:0] cmprep_local_bb1_cmp;
wire local_bb1_cmp;

assign cmprep_local_bb1_cmp = (local_bb1_inc45 - (input_wii_div1 & 32'h7FFFFFFF));
assign local_bb1_cmp = cmprep_local_bb1_cmp[32];

// This section implements an unregistered operation.
// 
wire local_bb1_var__stall_local;
wire local_bb1_var_;

assign local_bb1_var_ = (local_bb1_cmp & input_wii_var__u5);

// This section implements an unregistered operation.
// 
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_valid_out_0;
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_0;
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_valid_out_2;
wire local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_2;
wire local_bb1_inc45_valid_out_1;
wire local_bb1_inc45_stall_in_1;
wire local_bb1_var__valid_out;
wire local_bb1_var__stall_in;
wire local_bb1_cmp_not_valid_out;
wire local_bb1_cmp_not_stall_in;
wire local_bb1_cmp_not_inputs_ready;
wire local_bb1_cmp_not_stall_local;
wire local_bb1_cmp_not;
wire local_bb1_cmp_not_stall_out_local_or;
wire local_bb1_cmp_not_stall_local_fanout;
wire local_bb1_cmp_not_fu_valid_out_and;
 reg local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_0_NO_SHIFT_REG;
 reg local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_2_NO_SHIFT_REG;
 reg local_bb1_inc45_consumed_1_NO_SHIFT_REG;
 reg local_bb1_var__consumed_0_NO_SHIFT_REG;
 reg local_bb1_cmp_not_consumed_0_NO_SHIFT_REG;

assign local_bb1_cmp_not_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb1_pixel_y_020_pop8_acl_pop_i32_0_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb1_cmp_not = (local_bb1_cmp ^ 1'b1);
assign local_bb1_cmp_not_stall_out_local_or = local_bb1_pixel_y_020_pop8_acl_pop_i32_0_fu_stall_out;
assign local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_local = local_bb1_cmp_not_stall_local_fanout;
assign local_bb1_cmp_not_fu_valid_out_and = local_bb1_pixel_y_020_pop8_acl_pop_i32_0_fu_valid_out;
assign local_bb1_cmp_not_stall_local_fanout = ((local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_0 & ~(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_0_NO_SHIFT_REG)) | (local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_2 & ~(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_2_NO_SHIFT_REG)) | (local_bb1_inc45_stall_in_1 & ~(local_bb1_inc45_consumed_1_NO_SHIFT_REG)) | (local_bb1_var__stall_in & ~(local_bb1_var__consumed_0_NO_SHIFT_REG)) | (local_bb1_cmp_not_stall_in & ~(local_bb1_cmp_not_consumed_0_NO_SHIFT_REG)));
assign local_bb1_pixel_y_020_pop8_acl_pop_i32_0_valid_out_0 = (local_bb1_cmp_not_fu_valid_out_and & ~(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_0_NO_SHIFT_REG));
assign local_bb1_pixel_y_020_pop8_acl_pop_i32_0_valid_out_2 = (local_bb1_cmp_not_fu_valid_out_and & ~(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_2_NO_SHIFT_REG));
assign local_bb1_inc45_valid_out_1 = (local_bb1_cmp_not_fu_valid_out_and & ~(local_bb1_inc45_consumed_1_NO_SHIFT_REG));
assign local_bb1_var__valid_out = (local_bb1_cmp_not_fu_valid_out_and & ~(local_bb1_var__consumed_0_NO_SHIFT_REG));
assign local_bb1_cmp_not_valid_out = (local_bb1_cmp_not_fu_valid_out_and & ~(local_bb1_cmp_not_consumed_0_NO_SHIFT_REG));
assign merge_node_stall_in_0 = (|local_bb1_cmp_not_stall_out_local_or);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb1_inc45_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb1_var__consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb1_cmp_not_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_0_NO_SHIFT_REG <= (local_bb1_cmp_not_fu_valid_out_and & (local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_0_NO_SHIFT_REG | ~(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_0)) & local_bb1_cmp_not_stall_local_fanout);
		local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_2_NO_SHIFT_REG <= (local_bb1_cmp_not_fu_valid_out_and & (local_bb1_pixel_y_020_pop8_acl_pop_i32_0_consumed_2_NO_SHIFT_REG | ~(local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_2)) & local_bb1_cmp_not_stall_local_fanout);
		local_bb1_inc45_consumed_1_NO_SHIFT_REG <= (local_bb1_cmp_not_fu_valid_out_and & (local_bb1_inc45_consumed_1_NO_SHIFT_REG | ~(local_bb1_inc45_stall_in_1)) & local_bb1_cmp_not_stall_local_fanout);
		local_bb1_var__consumed_0_NO_SHIFT_REG <= (local_bb1_cmp_not_fu_valid_out_and & (local_bb1_var__consumed_0_NO_SHIFT_REG | ~(local_bb1_var__stall_in)) & local_bb1_cmp_not_stall_local_fanout);
		local_bb1_cmp_not_consumed_0_NO_SHIFT_REG <= (local_bb1_cmp_not_fu_valid_out_and & (local_bb1_cmp_not_consumed_0_NO_SHIFT_REG | ~(local_bb1_cmp_not_stall_in)) & local_bb1_cmp_not_stall_local_fanout);
	end
end


// This section implements a registered operation.
// 
wire local_bb1_mul37_inputs_ready;
 reg local_bb1_mul37_valid_out_NO_SHIFT_REG;
wire local_bb1_mul37_stall_in;
wire local_bb1_mul37_output_regs_ready;
wire [31:0] local_bb1_mul37;
 reg local_bb1_mul37_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb1_mul37_valid_pipe_1_NO_SHIFT_REG;
wire local_bb1_mul37_causedstall;

acl_int_mult int_module_local_bb1_mul37 (
	.clock(clock),
	.dataa(local_bb1_pixel_y_020_pop8_acl_pop_i32_0),
	.datab((input_wii_div & 32'h7FFFFFFF)),
	.enable(local_bb1_mul37_output_regs_ready),
	.result(local_bb1_mul37)
);

defparam int_module_local_bb1_mul37.INPUT1_WIDTH = 32;
defparam int_module_local_bb1_mul37.INPUT2_WIDTH = 31;
defparam int_module_local_bb1_mul37.OUTPUT_WIDTH = 32;
defparam int_module_local_bb1_mul37.LATENCY = 3;
defparam int_module_local_bb1_mul37.SIGNED = 0;

assign local_bb1_mul37_inputs_ready = local_bb1_pixel_y_020_pop8_acl_pop_i32_0_valid_out_0;
assign local_bb1_mul37_output_regs_ready = (&(~(local_bb1_mul37_valid_out_NO_SHIFT_REG) | ~(local_bb1_mul37_stall_in)));
assign local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_0 = (~(local_bb1_mul37_output_regs_ready) | ~(local_bb1_mul37_inputs_ready));
assign local_bb1_mul37_causedstall = (local_bb1_mul37_inputs_ready && (~(local_bb1_mul37_output_regs_ready) && !(~(local_bb1_mul37_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul37_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb1_mul37_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul37_output_regs_ready)
		begin
			local_bb1_mul37_valid_pipe_0_NO_SHIFT_REG <= local_bb1_mul37_inputs_ready;
			local_bb1_mul37_valid_pipe_1_NO_SHIFT_REG <= local_bb1_mul37_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul37_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul37_output_regs_ready)
		begin
			local_bb1_mul37_valid_out_NO_SHIFT_REG <= local_bb1_mul37_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb1_mul37_stall_in))
			begin
				local_bb1_mul37_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_NO_SHIFT_REG;
 logic rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb1_pixel_y_020_pop8_acl_pop_i32_0),
	.data_out(rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb1_pixel_y_020_pop8_acl_pop_i32_0_valid_out_2;
assign local_bb1_pixel_y_020_pop8_acl_pop_i32_0_stall_in_2 = rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_NO_SHIFT_REG = rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_reg_4_NO_SHIFT_REG;
assign rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_in_reg_4_NO_SHIFT_REG = rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_in_NO_SHIFT_REG;
assign rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_valid_out_NO_SHIFT_REG = rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_valid_out_reg_4_NO_SHIFT_REG;

// This section implements a staging register.
// 
wire rstag_1to1_bb1_var__valid_out_0;
wire rstag_1to1_bb1_var__stall_in_0;
wire rstag_1to1_bb1_var__valid_out_1;
wire rstag_1to1_bb1_var__stall_in_1;
wire rstag_1to1_bb1_var__inputs_ready;
wire rstag_1to1_bb1_var__stall_local;
 reg rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG;
wire rstag_1to1_bb1_var__combined_valid;
 reg rstag_1to1_bb1_var__staging_reg_NO_SHIFT_REG;
wire rstag_1to1_bb1_var_;
 reg rstag_1to1_bb1_var__consumed_0_NO_SHIFT_REG;
 reg rstag_1to1_bb1_var__consumed_1_NO_SHIFT_REG;

assign rstag_1to1_bb1_var__inputs_ready = local_bb1_var__valid_out;
assign rstag_1to1_bb1_var_ = (rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG ? rstag_1to1_bb1_var__staging_reg_NO_SHIFT_REG : local_bb1_var_);
assign rstag_1to1_bb1_var__combined_valid = (rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG | rstag_1to1_bb1_var__inputs_ready);
assign rstag_1to1_bb1_var__stall_local = ((rstag_1to1_bb1_var__stall_in_0 & ~(rstag_1to1_bb1_var__consumed_0_NO_SHIFT_REG)) | (rstag_1to1_bb1_var__stall_in_1 & ~(rstag_1to1_bb1_var__consumed_1_NO_SHIFT_REG)));
assign rstag_1to1_bb1_var__valid_out_0 = (rstag_1to1_bb1_var__combined_valid & ~(rstag_1to1_bb1_var__consumed_0_NO_SHIFT_REG));
assign rstag_1to1_bb1_var__valid_out_1 = (rstag_1to1_bb1_var__combined_valid & ~(rstag_1to1_bb1_var__consumed_1_NO_SHIFT_REG));
assign local_bb1_var__stall_in = (|rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_1to1_bb1_var__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_1to1_bb1_var__stall_local)
		begin
			if (~(rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG))
			begin
				rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG <= rstag_1to1_bb1_var__inputs_ready;
			end
		end
		else
		begin
			rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_1to1_bb1_var__staging_valid_NO_SHIFT_REG))
		begin
			rstag_1to1_bb1_var__staging_reg_NO_SHIFT_REG <= local_bb1_var_;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_1to1_bb1_var__consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_1to1_bb1_var__consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_1to1_bb1_var__consumed_0_NO_SHIFT_REG <= (rstag_1to1_bb1_var__combined_valid & (rstag_1to1_bb1_var__consumed_0_NO_SHIFT_REG | ~(rstag_1to1_bb1_var__stall_in_0)) & rstag_1to1_bb1_var__stall_local);
		rstag_1to1_bb1_var__consumed_1_NO_SHIFT_REG <= (rstag_1to1_bb1_var__combined_valid & (rstag_1to1_bb1_var__consumed_1_NO_SHIFT_REG | ~(rstag_1to1_bb1_var__stall_in_1)) & rstag_1to1_bb1_var__stall_local);
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_bb1_cmp_not_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to4_bb1_cmp_not_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to4_bb1_cmp_not_0_NO_SHIFT_REG;
 logic rnode_1to4_bb1_cmp_not_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to4_bb1_cmp_not_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1_cmp_not_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1_cmp_not_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1_cmp_not_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_1to4_bb1_cmp_not_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_bb1_cmp_not_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_bb1_cmp_not_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_bb1_cmp_not_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_bb1_cmp_not_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb1_cmp_not),
	.data_out(rnode_1to4_bb1_cmp_not_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_bb1_cmp_not_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_bb1_cmp_not_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_1to4_bb1_cmp_not_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_bb1_cmp_not_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_bb1_cmp_not_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb1_cmp_not_valid_out;
assign local_bb1_cmp_not_stall_in = rnode_1to4_bb1_cmp_not_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_bb1_cmp_not_0_NO_SHIFT_REG = rnode_1to4_bb1_cmp_not_0_reg_4_NO_SHIFT_REG;
assign rnode_1to4_bb1_cmp_not_0_stall_in_reg_4_NO_SHIFT_REG = rnode_1to4_bb1_cmp_not_0_stall_in_NO_SHIFT_REG;
assign rnode_1to4_bb1_cmp_not_0_valid_out_NO_SHIFT_REG = rnode_1to4_bb1_cmp_not_0_valid_out_reg_4_NO_SHIFT_REG;

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_4to4_bb1_mul37_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul37_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb1_mul37_0_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul37_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb1_mul37_0_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul37_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul37_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul37_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_4to4_bb1_mul37_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to4_bb1_mul37_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to4_bb1_mul37_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_4to4_bb1_mul37_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_4to4_bb1_mul37_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb1_mul37),
	.data_out(rnode_4to4_bb1_mul37_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_4to4_bb1_mul37_0_reg_4_fifo.DEPTH = 3;
defparam rnode_4to4_bb1_mul37_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_4to4_bb1_mul37_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to4_bb1_mul37_0_reg_4_fifo.IMPL = "zl_reg";

assign rnode_4to4_bb1_mul37_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb1_mul37_valid_out_NO_SHIFT_REG;
assign local_bb1_mul37_stall_in = rnode_4to4_bb1_mul37_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb1_mul37_0_NO_SHIFT_REG = rnode_4to4_bb1_mul37_0_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb1_mul37_0_stall_in_reg_4_NO_SHIFT_REG = rnode_4to4_bb1_mul37_0_stall_in_NO_SHIFT_REG;
assign rnode_4to4_bb1_mul37_0_valid_out_NO_SHIFT_REG = rnode_4to4_bb1_mul37_0_valid_out_reg_4_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb1_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb1_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb1_var__0_NO_SHIFT_REG;
 logic rnode_1to2_bb1_var__0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb1_var__0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_var__0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_var__0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_var__0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb1_var__0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb1_var__0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb1_var__0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb1_var__0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb1_var__0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(rstag_1to1_bb1_var_),
	.data_out(rnode_1to2_bb1_var__0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb1_var__0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb1_var__0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb1_var__0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb1_var__0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb1_var__0_reg_2_inputs_ready_NO_SHIFT_REG = rstag_1to1_bb1_var__valid_out_0;
assign rstag_1to1_bb1_var__stall_in_0 = rnode_1to2_bb1_var__0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb1_var__0_NO_SHIFT_REG = rnode_1to2_bb1_var__0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb1_var__0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb1_var__0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb1_var__0_valid_out_NO_SHIFT_REG = rnode_1to2_bb1_var__0_valid_out_reg_2_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb1_pixel_y_020_push8_inc45_inputs_ready;
 reg local_bb1_pixel_y_020_push8_inc45_valid_out_NO_SHIFT_REG;
wire local_bb1_pixel_y_020_push8_inc45_stall_in;
wire local_bb1_pixel_y_020_push8_inc45_output_regs_ready;
wire [31:0] local_bb1_pixel_y_020_push8_inc45_result;
wire local_bb1_pixel_y_020_push8_inc45_fu_valid_out;
wire local_bb1_pixel_y_020_push8_inc45_fu_stall_out;
 reg [31:0] local_bb1_pixel_y_020_push8_inc45_NO_SHIFT_REG;
wire local_bb1_pixel_y_020_push8_inc45_causedstall;

acl_push local_bb1_pixel_y_020_push8_inc45_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rstag_1to1_bb1_var_),
	.predicate(1'b0),
	.data_in(local_bb1_inc45),
	.stall_out(local_bb1_pixel_y_020_push8_inc45_fu_stall_out),
	.valid_in(local_bb1_pixel_y_020_push8_inc45_inputs_ready),
	.valid_out(local_bb1_pixel_y_020_push8_inc45_fu_valid_out),
	.stall_in(~(local_bb1_pixel_y_020_push8_inc45_output_regs_ready)),
	.data_out(local_bb1_pixel_y_020_push8_inc45_result),
	.feedback_out(feedback_data_out_8),
	.feedback_valid_out(feedback_valid_out_8),
	.feedback_stall_in(feedback_stall_in_8)
);

defparam local_bb1_pixel_y_020_push8_inc45_feedback.STALLFREE = 0;
defparam local_bb1_pixel_y_020_push8_inc45_feedback.DATA_WIDTH = 32;
defparam local_bb1_pixel_y_020_push8_inc45_feedback.FIFO_DEPTH = 4;
defparam local_bb1_pixel_y_020_push8_inc45_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb1_pixel_y_020_push8_inc45_feedback.STYLE = "REGULAR";

assign local_bb1_pixel_y_020_push8_inc45_inputs_ready = (local_bb1_inc45_valid_out_1 & rstag_1to1_bb1_var__valid_out_1);
assign local_bb1_pixel_y_020_push8_inc45_output_regs_ready = (&(~(local_bb1_pixel_y_020_push8_inc45_valid_out_NO_SHIFT_REG) | ~(local_bb1_pixel_y_020_push8_inc45_stall_in)));
assign local_bb1_inc45_stall_in_1 = (local_bb1_pixel_y_020_push8_inc45_fu_stall_out | ~(local_bb1_pixel_y_020_push8_inc45_inputs_ready));
assign rstag_1to1_bb1_var__stall_in_1 = (local_bb1_pixel_y_020_push8_inc45_fu_stall_out | ~(local_bb1_pixel_y_020_push8_inc45_inputs_ready));
assign local_bb1_pixel_y_020_push8_inc45_causedstall = (local_bb1_pixel_y_020_push8_inc45_inputs_ready && (local_bb1_pixel_y_020_push8_inc45_fu_stall_out && !(~(local_bb1_pixel_y_020_push8_inc45_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_pixel_y_020_push8_inc45_NO_SHIFT_REG <= 'x;
		local_bb1_pixel_y_020_push8_inc45_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_pixel_y_020_push8_inc45_output_regs_ready)
		begin
			local_bb1_pixel_y_020_push8_inc45_NO_SHIFT_REG <= local_bb1_pixel_y_020_push8_inc45_result;
			local_bb1_pixel_y_020_push8_inc45_valid_out_NO_SHIFT_REG <= local_bb1_pixel_y_020_push8_inc45_fu_valid_out;
		end
		else
		begin
			if (~(local_bb1_pixel_y_020_push8_inc45_stall_in))
			begin
				local_bb1_pixel_y_020_push8_inc45_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1_notcmp11_valid_out;
wire local_bb1_notcmp11_stall_in;
wire local_bb1_notcmp11_inputs_ready;
wire local_bb1_notcmp11_stall_local;
wire local_bb1_notcmp11;

assign local_bb1_notcmp11_inputs_ready = rnode_1to4_bb1_cmp_not_0_valid_out_NO_SHIFT_REG;
assign local_bb1_notcmp11 = (input_wii_cmp19 | rnode_1to4_bb1_cmp_not_0_NO_SHIFT_REG);
assign local_bb1_notcmp11_valid_out = local_bb1_notcmp11_inputs_ready;
assign local_bb1_notcmp11_stall_local = local_bb1_notcmp11_stall_in;
assign rnode_1to4_bb1_cmp_not_0_stall_in_NO_SHIFT_REG = (|local_bb1_notcmp11_stall_local);

// This section implements a registered operation.
// 
wire local_bb1_notexitcond14__inputs_ready;
 reg local_bb1_notexitcond14__valid_out_NO_SHIFT_REG;
wire local_bb1_notexitcond14__stall_in;
wire local_bb1_notexitcond14__output_regs_ready;
wire local_bb1_notexitcond14__result;
wire local_bb1_notexitcond14__fu_valid_out;
wire local_bb1_notexitcond14__fu_stall_out;
 reg local_bb1_notexitcond14__NO_SHIFT_REG;
wire local_bb1_notexitcond14__causedstall;
wire [32:0] rci_rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_2;

acl_push local_bb1_notexitcond14__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(rnode_1to2_bb1_var__0_NO_SHIFT_REG),
	.stall_out(local_bb1_notexitcond14__fu_stall_out),
	.valid_in(local_bb1_notexitcond14__inputs_ready),
	.valid_out(local_bb1_notexitcond14__fu_valid_out),
	.stall_in(~(local_bb1_notexitcond14__output_regs_ready)),
	.data_out(local_bb1_notexitcond14__result),
	.feedback_out(feedback_data_out_7),
	.feedback_valid_out(feedback_valid_out_7),
	.feedback_stall_in(feedback_stall_in_7)
);

defparam local_bb1_notexitcond14__feedback.STALLFREE = 0;
defparam local_bb1_notexitcond14__feedback.DATA_WIDTH = 1;
defparam local_bb1_notexitcond14__feedback.FIFO_DEPTH = 2;
defparam local_bb1_notexitcond14__feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb1_notexitcond14__feedback.STYLE = "REGULAR";

assign local_bb1_notexitcond14__inputs_ready = rnode_1to2_bb1_var__0_valid_out_NO_SHIFT_REG;
assign local_bb1_notexitcond14__output_regs_ready = (&(~(local_bb1_notexitcond14__valid_out_NO_SHIFT_REG) | ~(local_bb1_notexitcond14__stall_in)));
assign rnode_1to2_bb1_var__0_stall_in_NO_SHIFT_REG = (local_bb1_notexitcond14__fu_stall_out | ~(local_bb1_notexitcond14__inputs_ready));
assign local_bb1_notexitcond14__causedstall = (local_bb1_notexitcond14__inputs_ready && (local_bb1_notexitcond14__fu_stall_out && !(~(local_bb1_notexitcond14__output_regs_ready))));
assign rci_rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_2[0] = local_bb1_memdep_phi1_pop9_acl_pop_i1_0_NO_SHIFT_REG;
assign rci_rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_2[32:1] = local_bb1_pixel_y_020_push8_inc45_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_notexitcond14__NO_SHIFT_REG <= 'x;
		local_bb1_notexitcond14__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_notexitcond14__output_regs_ready)
		begin
			local_bb1_notexitcond14__NO_SHIFT_REG <= local_bb1_notexitcond14__result;
			local_bb1_notexitcond14__valid_out_NO_SHIFT_REG <= local_bb1_notexitcond14__fu_valid_out;
		end
		else
		begin
			if (~(local_bb1_notexitcond14__stall_in))
			begin
				local_bb1_notexitcond14__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_valid_out_NO_SHIFT_REG;
 logic rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_in_NO_SHIFT_REG;
 logic [32:0] rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_NO_SHIFT_REG;
 logic rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [32:0] rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_NO_SHIFT_REG;
 logic rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_out_0_reg_4_IP_NO_SHIFT_REG;
 logic rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_out_0_reg_4_NO_SHIFT_REG;
wire [1:0] rci_rcnode_3to4_rc0_bb1_notexitcond14__0_reg_3;

acl_data_fifo rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_out_0_reg_4_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_2),
	.data_out(rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_NO_SHIFT_REG)
);

defparam rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_fifo.DEPTH = 3;
defparam rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_fifo.DATA_WIDTH = 33;
defparam rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_fifo.IMPL = "ll_reg";

assign rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_inputs_ready_NO_SHIFT_REG = (local_bb1_memdep_phi1_pop9_acl_pop_i1_0_valid_out_NO_SHIFT_REG & local_bb1_pixel_y_020_push8_inc45_valid_out_NO_SHIFT_REG);
assign rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_out_0_reg_4_NO_SHIFT_REG = (~(rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_inputs_ready_NO_SHIFT_REG) | rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_out_0_reg_4_IP_NO_SHIFT_REG);
assign local_bb1_memdep_phi1_pop9_acl_pop_i1_0_stall_in = rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_out_0_reg_4_NO_SHIFT_REG;
assign local_bb1_pixel_y_020_push8_inc45_stall_in = rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_out_0_reg_4_NO_SHIFT_REG;
assign rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_NO_SHIFT_REG = rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_reg_4_NO_SHIFT_REG;
assign rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_in_reg_4_NO_SHIFT_REG = rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_in_NO_SHIFT_REG;
assign rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_valid_out_NO_SHIFT_REG = rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_valid_out_reg_4_NO_SHIFT_REG;
assign rci_rcnode_3to4_rc0_bb1_notexitcond14__0_reg_3[0] = local_bb1_notexitcond14__NO_SHIFT_REG;
assign rci_rcnode_3to4_rc0_bb1_notexitcond14__0_reg_3[1] = local_bb1_keep_going13_acl_pipeline_1_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_3to4_rc0_bb1_notexitcond14__0_valid_out_NO_SHIFT_REG;
 logic rcnode_3to4_rc0_bb1_notexitcond14__0_stall_in_NO_SHIFT_REG;
 logic [1:0] rcnode_3to4_rc0_bb1_notexitcond14__0_NO_SHIFT_REG;
 logic rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [1:0] rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_NO_SHIFT_REG;
 logic rcnode_3to4_rc0_bb1_notexitcond14__0_valid_out_reg_4_NO_SHIFT_REG;
 logic rcnode_3to4_rc0_bb1_notexitcond14__0_stall_in_reg_4_NO_SHIFT_REG;
 logic rcnode_3to4_rc0_bb1_notexitcond14__0_stall_out_0_reg_4_IP_NO_SHIFT_REG;
 logic rcnode_3to4_rc0_bb1_notexitcond14__0_stall_out_0_reg_4_NO_SHIFT_REG;

acl_data_fifo rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_3to4_rc0_bb1_notexitcond14__0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rcnode_3to4_rc0_bb1_notexitcond14__0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rcnode_3to4_rc0_bb1_notexitcond14__0_stall_out_0_reg_4_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_3to4_rc0_bb1_notexitcond14__0_reg_3),
	.data_out(rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_NO_SHIFT_REG)
);

defparam rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_fifo.DEPTH = 1;
defparam rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_fifo.DATA_WIDTH = 2;
defparam rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_fifo.IMPL = "ll_reg";

assign rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_inputs_ready_NO_SHIFT_REG = (local_bb1_notexitcond14__valid_out_NO_SHIFT_REG & local_bb1_keep_going13_acl_pipeline_1_valid_out_NO_SHIFT_REG);
assign rcnode_3to4_rc0_bb1_notexitcond14__0_stall_out_0_reg_4_NO_SHIFT_REG = (~(rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_inputs_ready_NO_SHIFT_REG) | rcnode_3to4_rc0_bb1_notexitcond14__0_stall_out_0_reg_4_IP_NO_SHIFT_REG);
assign local_bb1_notexitcond14__stall_in = rcnode_3to4_rc0_bb1_notexitcond14__0_stall_out_0_reg_4_NO_SHIFT_REG;
assign local_bb1_keep_going13_acl_pipeline_1_stall_in = rcnode_3to4_rc0_bb1_notexitcond14__0_stall_out_0_reg_4_NO_SHIFT_REG;
assign rcnode_3to4_rc0_bb1_notexitcond14__0_NO_SHIFT_REG = rcnode_3to4_rc0_bb1_notexitcond14__0_reg_4_NO_SHIFT_REG;
assign rcnode_3to4_rc0_bb1_notexitcond14__0_stall_in_reg_4_NO_SHIFT_REG = rcnode_3to4_rc0_bb1_notexitcond14__0_stall_in_NO_SHIFT_REG;
assign rcnode_3to4_rc0_bb1_notexitcond14__0_valid_out_NO_SHIFT_REG = rcnode_3to4_rc0_bb1_notexitcond14__0_valid_out_reg_4_NO_SHIFT_REG;

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [31:0] lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb1_mul37_reg_NO_SHIFT_REG;
 reg lvb_bb1_notcmp11_reg_NO_SHIFT_REG;
 reg lvb_bb1_notexitcond14__reg_NO_SHIFT_REG;
 reg lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb1_notcmp11_valid_out & rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_valid_out_NO_SHIFT_REG & rnode_4to4_bb1_mul37_0_valid_out_NO_SHIFT_REG & rcnode_3to4_rc0_bb1_notexitcond14__0_valid_out_NO_SHIFT_REG & rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb1_notcmp11_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_4to4_bb1_mul37_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_3to4_rc0_bb1_notexitcond14__0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0 = lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0_reg_NO_SHIFT_REG;
assign lvb_bb1_mul37 = lvb_bb1_mul37_reg_NO_SHIFT_REG;
assign lvb_bb1_notcmp11 = lvb_bb1_notcmp11_reg_NO_SHIFT_REG;
assign lvb_bb1_notexitcond14_ = lvb_bb1_notexitcond14__reg_NO_SHIFT_REG;
assign lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0 = lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb1_mul37_reg_NO_SHIFT_REG <= 'x;
		lvb_bb1_notcmp11_reg_NO_SHIFT_REG <= 'x;
		lvb_bb1_notexitcond14__reg_NO_SHIFT_REG <= 'x;
		lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0_reg_NO_SHIFT_REG <= rnode_1to4_bb1_pixel_y_020_pop8_acl_pop_i32_0_0_NO_SHIFT_REG;
			lvb_bb1_mul37_reg_NO_SHIFT_REG <= rnode_4to4_bb1_mul37_0_NO_SHIFT_REG;
			lvb_bb1_notcmp11_reg_NO_SHIFT_REG <= local_bb1_notcmp11;
			lvb_bb1_notexitcond14__reg_NO_SHIFT_REG <= rcnode_3to4_rc0_bb1_notexitcond14__0_NO_SHIFT_REG[0];
			lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0_reg_NO_SHIFT_REG <= rcnode_2to4_rc0_bb1_memdep_phi1_pop9_acl_pop_i1_0_0_NO_SHIFT_REG[0];
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_2
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_inSize_x,
		input [63:0] 		input_in,
		input [31:0] 		input_wii_div,
		input [31:0] 		input_wii_div1,
		input 		input_wii_cmp19,
		input [31:0] 		input_wii_add7,
		input [31:0] 		input_wii_sub20,
		input [31:0] 		input_wii_sub22,
		input 		input_wii_var_,
		input 		input_wii_var__u6,
		input 		input_wii_var__u7,
		input 		input_wii_var__u8,
		input 		valid_in_0,
		output 		stall_out_0,
		input 		input_forked18_0,
		input [31:0] 		input_pixel_y_020_pop819_0,
		input [31:0] 		input_mul3722_0,
		input 		input_notcmp1125_0,
		input 		input_notexitcond1428_0,
		input 		input_memdep_phi1_pop931_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input 		input_forked18_1,
		input [31:0] 		input_pixel_y_020_pop819_1,
		input [31:0] 		input_mul3722_1,
		input 		input_notcmp1125_1,
		input 		input_notexitcond1428_1,
		input 		input_memdep_phi1_pop931_1,
		output 		valid_out,
		input 		stall_in,
		output [31:0] 		lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819,
		output [31:0] 		lvb_bb2_mul5,
		output [63:0] 		lvb_bb2_indvars_iv_pop10_acl_pop_i64_0,
		output [31:0] 		lvb_bb2_var_,
		output 		lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931,
		output 		lvb_bb2_memdep_phi1_or,
		output [31:0] 		lvb_bb2_ld_,
		output 		lvb_bb2_notcmp,
		output 		lvb_bb2_notexitcond9_,
		output [31:0] 		lvb_bb2_mul3722_pop13_mul3722,
		output 		lvb_bb2_notcmp1125_pop14_notcmp1125,
		output 		lvb_bb2_notexitcond1428_pop15_notexitcond1428,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		feedback_valid_in_12,
		output 		feedback_stall_out_12,
		input [31:0] 		feedback_data_in_12,
		input 		feedback_valid_in_10,
		output 		feedback_stall_out_10,
		input [63:0] 		feedback_data_in_10,
		output 		feedback_stall_out_4,
		input 		feedback_valid_in_5,
		output 		feedback_stall_out_5,
		input 		feedback_data_in_5,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		input 		feedback_valid_in_11,
		output 		feedback_stall_out_11,
		input 		feedback_data_in_11,
		input 		feedback_valid_in_16,
		output 		feedback_stall_out_16,
		input 		feedback_data_in_16,
		input 		feedback_valid_in_13,
		output 		feedback_stall_out_13,
		input [31:0] 		feedback_data_in_13,
		input 		feedback_valid_in_14,
		output 		feedback_stall_out_14,
		input 		feedback_data_in_14,
		input 		feedback_valid_in_15,
		output 		feedback_stall_out_15,
		input 		feedback_data_in_15,
		output 		feedback_valid_out_10,
		input 		feedback_stall_in_10,
		output [63:0] 		feedback_data_out_10,
		output 		feedback_valid_out_5,
		input 		feedback_stall_in_5,
		output 		feedback_data_out_5,
		output 		feedback_valid_out_12,
		input 		feedback_stall_in_12,
		output [31:0] 		feedback_data_out_12,
		output 		feedback_valid_out_16,
		input 		feedback_stall_in_16,
		output 		feedback_data_out_16,
		output 		feedback_valid_out_13,
		input 		feedback_stall_in_13,
		output [31:0] 		feedback_data_out_13,
		output 		feedback_valid_out_14,
		input 		feedback_stall_in_14,
		output 		feedback_data_out_14,
		output 		feedback_valid_out_15,
		input 		feedback_stall_in_15,
		output 		feedback_data_out_15,
		input [511:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [32:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [511:0] 		avm_local_bb2_ld__writedata,
		output [63:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		output 		local_bb2_ld__active,
		input 		clock2x
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_node_stall_in_8;
 reg merge_node_valid_out_8_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg input_forked18_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pixel_y_020_pop819_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul3722_0_staging_reg_NO_SHIFT_REG;
 reg input_notcmp1125_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1428_0_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_pop931_0_staging_reg_NO_SHIFT_REG;
 reg local_lvm_forked18_NO_SHIFT_REG;
 reg [31:0] local_lvm_pixel_y_020_pop819_NO_SHIFT_REG;
 reg [31:0] local_lvm_mul3722_NO_SHIFT_REG;
 reg local_lvm_notcmp1125_NO_SHIFT_REG;
 reg local_lvm_notexitcond1428_NO_SHIFT_REG;
 reg local_lvm_memdep_phi1_pop931_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg input_forked18_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pixel_y_020_pop819_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul3722_1_staging_reg_NO_SHIFT_REG;
 reg input_notcmp1125_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1428_1_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_pop931_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG) | (merge_node_stall_in_8 & merge_node_valid_out_8_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_forked18_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_pixel_y_020_pop819_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul3722_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp1125_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1428_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_pop931_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_forked18_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_pixel_y_020_pop819_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul3722_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp1125_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1428_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_pop931_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_forked18_0_staging_reg_NO_SHIFT_REG <= input_forked18_0;
				input_pixel_y_020_pop819_0_staging_reg_NO_SHIFT_REG <= input_pixel_y_020_pop819_0;
				input_mul3722_0_staging_reg_NO_SHIFT_REG <= input_mul3722_0;
				input_notcmp1125_0_staging_reg_NO_SHIFT_REG <= input_notcmp1125_0;
				input_notexitcond1428_0_staging_reg_NO_SHIFT_REG <= input_notexitcond1428_0;
				input_memdep_phi1_pop931_0_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_pop931_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_forked18_1_staging_reg_NO_SHIFT_REG <= input_forked18_1;
				input_pixel_y_020_pop819_1_staging_reg_NO_SHIFT_REG <= input_pixel_y_020_pop819_1;
				input_mul3722_1_staging_reg_NO_SHIFT_REG <= input_mul3722_1;
				input_notcmp1125_1_staging_reg_NO_SHIFT_REG <= input_notcmp1125_1;
				input_notexitcond1428_1_staging_reg_NO_SHIFT_REG <= input_notexitcond1428_1;
				input_memdep_phi1_pop931_1_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_pop931_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked18_NO_SHIFT_REG <= input_forked18_0_staging_reg_NO_SHIFT_REG;
					local_lvm_pixel_y_020_pop819_NO_SHIFT_REG <= input_pixel_y_020_pop819_0_staging_reg_NO_SHIFT_REG;
					local_lvm_mul3722_NO_SHIFT_REG <= input_mul3722_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp1125_NO_SHIFT_REG <= input_notcmp1125_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1428_NO_SHIFT_REG <= input_notexitcond1428_0_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_pop931_NO_SHIFT_REG <= input_memdep_phi1_pop931_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked18_NO_SHIFT_REG <= input_forked18_0;
					local_lvm_pixel_y_020_pop819_NO_SHIFT_REG <= input_pixel_y_020_pop819_0;
					local_lvm_mul3722_NO_SHIFT_REG <= input_mul3722_0;
					local_lvm_notcmp1125_NO_SHIFT_REG <= input_notcmp1125_0;
					local_lvm_notexitcond1428_NO_SHIFT_REG <= input_notexitcond1428_0;
					local_lvm_memdep_phi1_pop931_NO_SHIFT_REG <= input_memdep_phi1_pop931_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked18_NO_SHIFT_REG <= input_forked18_1_staging_reg_NO_SHIFT_REG;
					local_lvm_pixel_y_020_pop819_NO_SHIFT_REG <= input_pixel_y_020_pop819_1_staging_reg_NO_SHIFT_REG;
					local_lvm_mul3722_NO_SHIFT_REG <= input_mul3722_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp1125_NO_SHIFT_REG <= input_notcmp1125_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1428_NO_SHIFT_REG <= input_notexitcond1428_1_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_pop931_NO_SHIFT_REG <= input_memdep_phi1_pop931_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked18_NO_SHIFT_REG <= input_forked18_1;
					local_lvm_pixel_y_020_pop819_NO_SHIFT_REG <= input_pixel_y_020_pop819_1;
					local_lvm_mul3722_NO_SHIFT_REG <= input_mul3722_1;
					local_lvm_notcmp1125_NO_SHIFT_REG <= input_notcmp1125_1;
					local_lvm_notexitcond1428_NO_SHIFT_REG <= input_notexitcond1428_1;
					local_lvm_memdep_phi1_pop931_NO_SHIFT_REG <= input_memdep_phi1_pop931_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_8_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_8))
			begin
				merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_inputs_ready;
 reg local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_0_NO_SHIFT_REG;
wire local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_0;
 reg local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_1_NO_SHIFT_REG;
wire local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_1;
wire local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_output_regs_ready;
wire [31:0] local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_result;
wire local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_valid_out;
wire local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_stall_out;
 reg [31:0] local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_NO_SHIFT_REG;
wire local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_causedstall;

acl_pop local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_forked18_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_lvm_pixel_y_020_pop819_NO_SHIFT_REG),
	.stall_out(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_stall_out),
	.valid_in(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_inputs_ready),
	.valid_out(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_valid_out),
	.stall_in(~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_output_regs_ready)),
	.data_out(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_result),
	.feedback_in(feedback_data_in_12),
	.feedback_valid_in(feedback_valid_in_12),
	.feedback_stall_out(feedback_stall_out_12)
);

defparam local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_feedback.COALESCE_DISTANCE = 1;
defparam local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_feedback.DATA_WIDTH = 32;
defparam local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_feedback.STYLE = "REGULAR";

assign local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_output_regs_ready = ((~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_0_NO_SHIFT_REG) | ~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_0)) & (~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_1_NO_SHIFT_REG) | ~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_1)));
assign merge_node_stall_in_0 = (local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_stall_out | ~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_inputs_ready));
assign local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_causedstall = (local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_inputs_ready && (local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_stall_out && !(~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_NO_SHIFT_REG <= 'x;
		local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_output_regs_ready)
		begin
			local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_NO_SHIFT_REG <= local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_result;
			local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_0_NO_SHIFT_REG <= local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_valid_out;
			local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_1_NO_SHIFT_REG <= local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_0))
			begin
				local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_1))
			begin
				local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_indvars_iv_pop10_acl_pop_i64_0_stall_local;
wire [63:0] local_bb2_indvars_iv_pop10_acl_pop_i64_0;
wire local_bb2_indvars_iv_pop10_acl_pop_i64_0_fu_valid_out;
wire local_bb2_indvars_iv_pop10_acl_pop_i64_0_fu_stall_out;
wire local_bb2_indvars_iv_pop10_acl_pop_i64_0_inputs_ready;

acl_pop local_bb2_indvars_iv_pop10_acl_pop_i64_0_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_forked18_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(64'h0),
	.stall_out(local_bb2_indvars_iv_pop10_acl_pop_i64_0_fu_stall_out),
	.valid_in(local_bb2_indvars_iv_pop10_acl_pop_i64_0_inputs_ready),
	.valid_out(local_bb2_indvars_iv_pop10_acl_pop_i64_0_fu_valid_out),
	.stall_in(local_bb2_indvars_iv_pop10_acl_pop_i64_0_stall_local),
	.data_out(local_bb2_indvars_iv_pop10_acl_pop_i64_0),
	.feedback_in(feedback_data_in_10),
	.feedback_valid_in(feedback_valid_in_10),
	.feedback_stall_out(feedback_stall_out_10)
);

defparam local_bb2_indvars_iv_pop10_acl_pop_i64_0_feedback.COALESCE_DISTANCE = 1;
defparam local_bb2_indvars_iv_pop10_acl_pop_i64_0_feedback.DATA_WIDTH = 64;
defparam local_bb2_indvars_iv_pop10_acl_pop_i64_0_feedback.STYLE = "REGULAR";


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_fifo.DATA_WIDTH = 0;
defparam rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_reg_2_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign merge_node_stall_in_2 = rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_valid_out_reg_2_NO_SHIFT_REG;

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_1to6_forked18_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to6_forked18_1_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_1to6_forked18_2_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_1to6_forked18_3_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_stall_in_4_NO_SHIFT_REG;
 logic rnode_1to6_forked18_4_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_forked18_0_stall_out_reg_6_NO_SHIFT_REG;
 reg rnode_1to6_forked18_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to6_forked18_0_consumed_1_NO_SHIFT_REG;
 reg rnode_1to6_forked18_0_consumed_2_NO_SHIFT_REG;
 reg rnode_1to6_forked18_0_consumed_3_NO_SHIFT_REG;
 reg rnode_1to6_forked18_0_consumed_4_NO_SHIFT_REG;

acl_data_fifo rnode_1to6_forked18_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to6_forked18_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_1to6_forked18_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_lvm_forked18_NO_SHIFT_REG),
	.data_out(rnode_1to6_forked18_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_1to6_forked18_0_reg_6_fifo.DEPTH = 6;
defparam rnode_1to6_forked18_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_1to6_forked18_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to6_forked18_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_1to6_forked18_0_reg_6_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_3_NO_SHIFT_REG;
assign merge_node_stall_in_3 = rnode_1to6_forked18_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG = ((rnode_1to6_forked18_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to6_forked18_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_1_NO_SHIFT_REG)) | (rnode_1to6_forked18_0_stall_in_2_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_2_NO_SHIFT_REG)) | (rnode_1to6_forked18_0_stall_in_3_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_3_NO_SHIFT_REG)) | (rnode_1to6_forked18_0_stall_in_4_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_4_NO_SHIFT_REG)));
assign rnode_1to6_forked18_0_valid_out_0_NO_SHIFT_REG = (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to6_forked18_0_valid_out_1_NO_SHIFT_REG = (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to6_forked18_0_valid_out_2_NO_SHIFT_REG = (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_2_NO_SHIFT_REG));
assign rnode_1to6_forked18_0_valid_out_3_NO_SHIFT_REG = (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_3_NO_SHIFT_REG));
assign rnode_1to6_forked18_0_valid_out_4_NO_SHIFT_REG = (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & ~(rnode_1to6_forked18_0_consumed_4_NO_SHIFT_REG));
assign rnode_1to6_forked18_0_NO_SHIFT_REG = rnode_1to6_forked18_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_forked18_1_NO_SHIFT_REG = rnode_1to6_forked18_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_forked18_2_NO_SHIFT_REG = rnode_1to6_forked18_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_forked18_3_NO_SHIFT_REG = rnode_1to6_forked18_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_forked18_4_NO_SHIFT_REG = rnode_1to6_forked18_0_reg_6_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to6_forked18_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to6_forked18_0_consumed_1_NO_SHIFT_REG <= 1'b0;
		rnode_1to6_forked18_0_consumed_2_NO_SHIFT_REG <= 1'b0;
		rnode_1to6_forked18_0_consumed_3_NO_SHIFT_REG <= 1'b0;
		rnode_1to6_forked18_0_consumed_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to6_forked18_0_consumed_0_NO_SHIFT_REG <= (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & (rnode_1to6_forked18_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to6_forked18_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG);
		rnode_1to6_forked18_0_consumed_1_NO_SHIFT_REG <= (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & (rnode_1to6_forked18_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to6_forked18_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG);
		rnode_1to6_forked18_0_consumed_2_NO_SHIFT_REG <= (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & (rnode_1to6_forked18_0_consumed_2_NO_SHIFT_REG | ~(rnode_1to6_forked18_0_stall_in_2_NO_SHIFT_REG)) & rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG);
		rnode_1to6_forked18_0_consumed_3_NO_SHIFT_REG <= (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & (rnode_1to6_forked18_0_consumed_3_NO_SHIFT_REG | ~(rnode_1to6_forked18_0_stall_in_3_NO_SHIFT_REG)) & rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG);
		rnode_1to6_forked18_0_consumed_4_NO_SHIFT_REG <= (rnode_1to6_forked18_0_valid_out_0_reg_6_NO_SHIFT_REG & (rnode_1to6_forked18_0_consumed_4_NO_SHIFT_REG | ~(rnode_1to6_forked18_0_stall_in_4_NO_SHIFT_REG)) & rnode_1to6_forked18_0_stall_in_0_reg_6_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_1to6_memdep_phi1_pop931_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to6_memdep_phi1_pop931_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to6_memdep_phi1_pop931_0_NO_SHIFT_REG;
 logic rnode_1to6_memdep_phi1_pop931_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to6_memdep_phi1_pop931_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_memdep_phi1_pop931_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_memdep_phi1_pop931_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_memdep_phi1_pop931_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_1to6_memdep_phi1_pop931_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to6_memdep_phi1_pop931_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to6_memdep_phi1_pop931_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_1to6_memdep_phi1_pop931_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_1to6_memdep_phi1_pop931_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_lvm_memdep_phi1_pop931_NO_SHIFT_REG),
	.data_out(rnode_1to6_memdep_phi1_pop931_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_1to6_memdep_phi1_pop931_0_reg_6_fifo.DEPTH = 6;
defparam rnode_1to6_memdep_phi1_pop931_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_1to6_memdep_phi1_pop931_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to6_memdep_phi1_pop931_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_1to6_memdep_phi1_pop931_0_reg_6_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_4_NO_SHIFT_REG;
assign merge_node_stall_in_4 = rnode_1to6_memdep_phi1_pop931_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_1to6_memdep_phi1_pop931_0_NO_SHIFT_REG = rnode_1to6_memdep_phi1_pop931_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_memdep_phi1_pop931_0_stall_in_reg_6_NO_SHIFT_REG = rnode_1to6_memdep_phi1_pop931_0_stall_in_NO_SHIFT_REG;
assign rnode_1to6_memdep_phi1_pop931_0_valid_out_NO_SHIFT_REG = rnode_1to6_memdep_phi1_pop931_0_valid_out_reg_6_NO_SHIFT_REG;

// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_1to7_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_1to7_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_1to7_var__0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to7_var__0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_1to7_var__0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_1to7_var__0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_1to7_var__0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to7_var__0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to7_var__0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_1to7_var__0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_1to7_var__0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to7_var__0_reg_7_fifo.DEPTH = 7;
defparam rnode_1to7_var__0_reg_7_fifo.DATA_WIDTH = 0;
defparam rnode_1to7_var__0_reg_7_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to7_var__0_reg_7_fifo.IMPL = "ll_reg";

assign rnode_1to7_var__0_reg_7_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign merge_node_stall_in_5 = rnode_1to7_var__0_stall_out_reg_7_NO_SHIFT_REG;
assign rnode_1to7_var__0_stall_in_reg_7_NO_SHIFT_REG = rnode_1to7_var__0_stall_in_NO_SHIFT_REG;
assign rnode_1to7_var__0_valid_out_NO_SHIFT_REG = rnode_1to7_var__0_valid_out_reg_7_NO_SHIFT_REG;

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_1to6_mul3722_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to6_mul3722_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to6_mul3722_0_NO_SHIFT_REG;
 logic rnode_1to6_mul3722_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to6_mul3722_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_mul3722_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_mul3722_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_mul3722_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_1to6_mul3722_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to6_mul3722_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to6_mul3722_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_1to6_mul3722_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_1to6_mul3722_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_lvm_mul3722_NO_SHIFT_REG),
	.data_out(rnode_1to6_mul3722_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_1to6_mul3722_0_reg_6_fifo.DEPTH = 6;
defparam rnode_1to6_mul3722_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_1to6_mul3722_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to6_mul3722_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_1to6_mul3722_0_reg_6_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_6_NO_SHIFT_REG;
assign merge_node_stall_in_6 = rnode_1to6_mul3722_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_1to6_mul3722_0_NO_SHIFT_REG = rnode_1to6_mul3722_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_mul3722_0_stall_in_reg_6_NO_SHIFT_REG = rnode_1to6_mul3722_0_stall_in_NO_SHIFT_REG;
assign rnode_1to6_mul3722_0_valid_out_NO_SHIFT_REG = rnode_1to6_mul3722_0_valid_out_reg_6_NO_SHIFT_REG;

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_1to6_notcmp1125_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to6_notcmp1125_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to6_notcmp1125_0_NO_SHIFT_REG;
 logic rnode_1to6_notcmp1125_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to6_notcmp1125_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_notcmp1125_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_notcmp1125_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_notcmp1125_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_1to6_notcmp1125_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to6_notcmp1125_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to6_notcmp1125_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_1to6_notcmp1125_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_1to6_notcmp1125_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_lvm_notcmp1125_NO_SHIFT_REG),
	.data_out(rnode_1to6_notcmp1125_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_1to6_notcmp1125_0_reg_6_fifo.DEPTH = 6;
defparam rnode_1to6_notcmp1125_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_1to6_notcmp1125_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to6_notcmp1125_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_1to6_notcmp1125_0_reg_6_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_7_NO_SHIFT_REG;
assign merge_node_stall_in_7 = rnode_1to6_notcmp1125_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_1to6_notcmp1125_0_NO_SHIFT_REG = rnode_1to6_notcmp1125_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_notcmp1125_0_stall_in_reg_6_NO_SHIFT_REG = rnode_1to6_notcmp1125_0_stall_in_NO_SHIFT_REG;
assign rnode_1to6_notcmp1125_0_valid_out_NO_SHIFT_REG = rnode_1to6_notcmp1125_0_valid_out_reg_6_NO_SHIFT_REG;

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_1to6_notexitcond1428_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to6_notexitcond1428_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to6_notexitcond1428_0_NO_SHIFT_REG;
 logic rnode_1to6_notexitcond1428_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to6_notexitcond1428_0_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_notexitcond1428_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_notexitcond1428_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_1to6_notexitcond1428_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_1to6_notexitcond1428_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to6_notexitcond1428_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to6_notexitcond1428_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_1to6_notexitcond1428_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_1to6_notexitcond1428_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_lvm_notexitcond1428_NO_SHIFT_REG),
	.data_out(rnode_1to6_notexitcond1428_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_1to6_notexitcond1428_0_reg_6_fifo.DEPTH = 6;
defparam rnode_1to6_notexitcond1428_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_1to6_notexitcond1428_0_reg_6_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to6_notexitcond1428_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_1to6_notexitcond1428_0_reg_6_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_8_NO_SHIFT_REG;
assign merge_node_stall_in_8 = rnode_1to6_notexitcond1428_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_1to6_notexitcond1428_0_NO_SHIFT_REG = rnode_1to6_notexitcond1428_0_reg_6_NO_SHIFT_REG;
assign rnode_1to6_notexitcond1428_0_stall_in_reg_6_NO_SHIFT_REG = rnode_1to6_notexitcond1428_0_stall_in_NO_SHIFT_REG;
assign rnode_1to6_notexitcond1428_0_valid_out_NO_SHIFT_REG = rnode_1to6_notexitcond1428_0_valid_out_reg_6_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_mul5_valid_out_0;
wire local_bb2_mul5_stall_in_0;
wire local_bb2_mul5_valid_out_1;
wire local_bb2_mul5_stall_in_1;
wire local_bb2_mul5_inputs_ready;
wire local_bb2_mul5_stall_local;
wire [31:0] local_bb2_mul5;
 reg local_bb2_mul5_consumed_0_NO_SHIFT_REG;
 reg local_bb2_mul5_consumed_1_NO_SHIFT_REG;

assign local_bb2_mul5_inputs_ready = local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_0_NO_SHIFT_REG;
assign local_bb2_mul5 = (local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_NO_SHIFT_REG << 32'h1);
assign local_bb2_mul5_stall_local = ((local_bb2_mul5_stall_in_0 & ~(local_bb2_mul5_consumed_0_NO_SHIFT_REG)) | (local_bb2_mul5_stall_in_1 & ~(local_bb2_mul5_consumed_1_NO_SHIFT_REG)));
assign local_bb2_mul5_valid_out_0 = (local_bb2_mul5_inputs_ready & ~(local_bb2_mul5_consumed_0_NO_SHIFT_REG));
assign local_bb2_mul5_valid_out_1 = (local_bb2_mul5_inputs_ready & ~(local_bb2_mul5_consumed_1_NO_SHIFT_REG));
assign local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_0 = (|local_bb2_mul5_stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul5_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul5_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_mul5_consumed_0_NO_SHIFT_REG <= (local_bb2_mul5_inputs_ready & (local_bb2_mul5_consumed_0_NO_SHIFT_REG | ~(local_bb2_mul5_stall_in_0)) & local_bb2_mul5_stall_local);
		local_bb2_mul5_consumed_1_NO_SHIFT_REG <= (local_bb2_mul5_inputs_ready & (local_bb2_mul5_consumed_1_NO_SHIFT_REG | ~(local_bb2_mul5_stall_in_1)) & local_bb2_mul5_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_NO_SHIFT_REG;
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_1_NO_SHIFT_REG;
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_reg_3_NO_SHIFT_REG;
 reg rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_0_NO_SHIFT_REG;
 reg rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_NO_SHIFT_REG),
	.data_out(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_valid_out_1_NO_SHIFT_REG;
assign local_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_stall_in_1 = rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_reg_3_NO_SHIFT_REG = ((rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_NO_SHIFT_REG & ~(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_0_NO_SHIFT_REG)) | (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_1_NO_SHIFT_REG & ~(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_1_NO_SHIFT_REG)));
assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_NO_SHIFT_REG = (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_reg_3_NO_SHIFT_REG & ~(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_0_NO_SHIFT_REG));
assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_1_NO_SHIFT_REG = (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_reg_3_NO_SHIFT_REG & ~(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_1_NO_SHIFT_REG));
assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_NO_SHIFT_REG = rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_1_NO_SHIFT_REG = rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_0_NO_SHIFT_REG <= (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_reg_3_NO_SHIFT_REG & (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_0_NO_SHIFT_REG | ~(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_NO_SHIFT_REG)) & rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_reg_3_NO_SHIFT_REG);
		rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_1_NO_SHIFT_REG <= (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_reg_3_NO_SHIFT_REG & (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_consumed_1_NO_SHIFT_REG | ~(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_1_NO_SHIFT_REG)) & rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_reg_3_NO_SHIFT_REG);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_indvars_iv_next_stall_local;
wire [63:0] local_bb2_indvars_iv_next;

assign local_bb2_indvars_iv_next = (local_bb2_indvars_iv_pop10_acl_pop_i64_0 + 64'h1);

// This section implements a registered operation.
// 
wire local_bb2_keep_going8_acl_pipeline_1_inputs_ready;
 reg local_bb2_keep_going8_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb2_keep_going8_acl_pipeline_1_stall_in;
wire local_bb2_keep_going8_acl_pipeline_1_output_regs_ready;
wire local_bb2_keep_going8_acl_pipeline_1_keep_going;
wire local_bb2_keep_going8_acl_pipeline_1_fu_valid_out;
wire local_bb2_keep_going8_acl_pipeline_1_fu_stall_out;
 reg local_bb2_keep_going8_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb2_keep_going8_acl_pipeline_1_feedback_pipelined;
wire local_bb2_keep_going8_acl_pipeline_1_causedstall;

acl_pipeline local_bb2_keep_going8_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb2_keep_going8_acl_pipeline_1_fu_stall_out),
	.valid_in(local_bb2_keep_going8_acl_pipeline_1_inputs_ready),
	.valid_out(local_bb2_keep_going8_acl_pipeline_1_fu_valid_out),
	.stall_in(~(local_bb2_keep_going8_acl_pipeline_1_output_regs_ready)),
	.data_out(local_bb2_keep_going8_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_4),
	.not_exitcond_in(feedback_data_in_5),
	.not_exitcond_valid_in(feedback_valid_in_5),
	.not_exitcond_stall_out(feedback_stall_out_5),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb2_keep_going8_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb2_keep_going8_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb2_keep_going8_acl_pipeline_1_inputs_ready = rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
assign local_bb2_keep_going8_acl_pipeline_1_output_regs_ready = (&(~(local_bb2_keep_going8_acl_pipeline_1_valid_out_NO_SHIFT_REG) | ~(local_bb2_keep_going8_acl_pipeline_1_stall_in)));
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign rnode_1to2_bb2_keep_going8_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = (local_bb2_keep_going8_acl_pipeline_1_fu_stall_out | ~(local_bb2_keep_going8_acl_pipeline_1_inputs_ready));
assign local_bb2_keep_going8_acl_pipeline_1_causedstall = (local_bb2_keep_going8_acl_pipeline_1_inputs_ready && (local_bb2_keep_going8_acl_pipeline_1_fu_stall_out && !(~(local_bb2_keep_going8_acl_pipeline_1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_keep_going8_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb2_keep_going8_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_keep_going8_acl_pipeline_1_output_regs_ready)
		begin
			local_bb2_keep_going8_acl_pipeline_1_NO_SHIFT_REG <= local_bb2_keep_going8_acl_pipeline_1_keep_going;
			local_bb2_keep_going8_acl_pipeline_1_valid_out_NO_SHIFT_REG <= local_bb2_keep_going8_acl_pipeline_1_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_keep_going8_acl_pipeline_1_stall_in))
			begin
				local_bb2_keep_going8_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_memdep_phi_pop11_acl_pop_i1_0_inputs_ready;
 reg local_bb2_memdep_phi_pop11_acl_pop_i1_0_valid_out_NO_SHIFT_REG;
wire local_bb2_memdep_phi_pop11_acl_pop_i1_0_stall_in;
wire local_bb2_memdep_phi_pop11_acl_pop_i1_0_output_regs_ready;
wire local_bb2_memdep_phi_pop11_acl_pop_i1_0_result;
wire local_bb2_memdep_phi_pop11_acl_pop_i1_0_fu_valid_out;
wire local_bb2_memdep_phi_pop11_acl_pop_i1_0_fu_stall_out;
 reg local_bb2_memdep_phi_pop11_acl_pop_i1_0_NO_SHIFT_REG;
wire local_bb2_memdep_phi_pop11_acl_pop_i1_0_causedstall;

acl_pop local_bb2_memdep_phi_pop11_acl_pop_i1_0_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to6_forked18_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(1'b0),
	.stall_out(local_bb2_memdep_phi_pop11_acl_pop_i1_0_fu_stall_out),
	.valid_in(local_bb2_memdep_phi_pop11_acl_pop_i1_0_inputs_ready),
	.valid_out(local_bb2_memdep_phi_pop11_acl_pop_i1_0_fu_valid_out),
	.stall_in(~(local_bb2_memdep_phi_pop11_acl_pop_i1_0_output_regs_ready)),
	.data_out(local_bb2_memdep_phi_pop11_acl_pop_i1_0_result),
	.feedback_in(feedback_data_in_11),
	.feedback_valid_in(feedback_valid_in_11),
	.feedback_stall_out(feedback_stall_out_11)
);

defparam local_bb2_memdep_phi_pop11_acl_pop_i1_0_feedback.COALESCE_DISTANCE = 1;
defparam local_bb2_memdep_phi_pop11_acl_pop_i1_0_feedback.DATA_WIDTH = 1;
defparam local_bb2_memdep_phi_pop11_acl_pop_i1_0_feedback.STYLE = "REGULAR";

assign local_bb2_memdep_phi_pop11_acl_pop_i1_0_inputs_ready = rnode_1to6_forked18_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_memdep_phi_pop11_acl_pop_i1_0_output_regs_ready = (&(~(local_bb2_memdep_phi_pop11_acl_pop_i1_0_valid_out_NO_SHIFT_REG) | ~(local_bb2_memdep_phi_pop11_acl_pop_i1_0_stall_in)));
assign rnode_1to6_forked18_0_stall_in_0_NO_SHIFT_REG = (local_bb2_memdep_phi_pop11_acl_pop_i1_0_fu_stall_out | ~(local_bb2_memdep_phi_pop11_acl_pop_i1_0_inputs_ready));
assign local_bb2_memdep_phi_pop11_acl_pop_i1_0_causedstall = (local_bb2_memdep_phi_pop11_acl_pop_i1_0_inputs_ready && (local_bb2_memdep_phi_pop11_acl_pop_i1_0_fu_stall_out && !(~(local_bb2_memdep_phi_pop11_acl_pop_i1_0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_memdep_phi_pop11_acl_pop_i1_0_NO_SHIFT_REG <= 'x;
		local_bb2_memdep_phi_pop11_acl_pop_i1_0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_memdep_phi_pop11_acl_pop_i1_0_output_regs_ready)
		begin
			local_bb2_memdep_phi_pop11_acl_pop_i1_0_NO_SHIFT_REG <= local_bb2_memdep_phi_pop11_acl_pop_i1_0_result;
			local_bb2_memdep_phi_pop11_acl_pop_i1_0_valid_out_NO_SHIFT_REG <= local_bb2_memdep_phi_pop11_acl_pop_i1_0_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_memdep_phi_pop11_acl_pop_i1_0_stall_in))
			begin
				local_bb2_memdep_phi_pop11_acl_pop_i1_0_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_inputs_ready;
 reg local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_0_NO_SHIFT_REG;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_0;
 reg local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_1_NO_SHIFT_REG;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_1;
 reg local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_2_NO_SHIFT_REG;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_2;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_output_regs_ready;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_result;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_valid_out;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_stall_out;
 reg local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_NO_SHIFT_REG;
wire local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_causedstall;

acl_pop local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to6_forked18_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to6_memdep_phi1_pop931_0_NO_SHIFT_REG),
	.stall_out(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_stall_out),
	.valid_in(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_inputs_ready),
	.valid_out(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_valid_out),
	.stall_in(~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_output_regs_ready)),
	.data_out(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_result),
	.feedback_in(feedback_data_in_16),
	.feedback_valid_in(feedback_valid_in_16),
	.feedback_stall_out(feedback_stall_out_16)
);

defparam local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_feedback.COALESCE_DISTANCE = 1;
defparam local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_feedback.DATA_WIDTH = 1;
defparam local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_feedback.STYLE = "REGULAR";

assign local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_inputs_ready = (rnode_1to6_memdep_phi1_pop931_0_valid_out_NO_SHIFT_REG & rnode_1to6_forked18_0_valid_out_1_NO_SHIFT_REG);
assign local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_output_regs_ready = ((~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_0_NO_SHIFT_REG) | ~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_0)) & (~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_1_NO_SHIFT_REG) | ~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_1)) & (~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_2_NO_SHIFT_REG) | ~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_2)));
assign rnode_1to6_memdep_phi1_pop931_0_stall_in_NO_SHIFT_REG = (local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_stall_out | ~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_inputs_ready));
assign rnode_1to6_forked18_0_stall_in_1_NO_SHIFT_REG = (local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_stall_out | ~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_inputs_ready));
assign local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_causedstall = (local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_inputs_ready && (local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_stall_out && !(~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_NO_SHIFT_REG <= 'x;
		local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_output_regs_ready)
		begin
			local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_NO_SHIFT_REG <= local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_result;
			local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_0_NO_SHIFT_REG <= local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_valid_out;
			local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_1_NO_SHIFT_REG <= local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_valid_out;
			local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_2_NO_SHIFT_REG <= local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_0))
			begin
				local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_1))
			begin
				local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_2))
			begin
				local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul3722_pop13_mul3722_inputs_ready;
 reg local_bb2_mul3722_pop13_mul3722_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul3722_pop13_mul3722_stall_in_0;
 reg local_bb2_mul3722_pop13_mul3722_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul3722_pop13_mul3722_stall_in_1;
wire local_bb2_mul3722_pop13_mul3722_output_regs_ready;
wire [31:0] local_bb2_mul3722_pop13_mul3722_result;
wire local_bb2_mul3722_pop13_mul3722_fu_valid_out;
wire local_bb2_mul3722_pop13_mul3722_fu_stall_out;
 reg [31:0] local_bb2_mul3722_pop13_mul3722_NO_SHIFT_REG;
wire local_bb2_mul3722_pop13_mul3722_causedstall;

acl_pop local_bb2_mul3722_pop13_mul3722_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to6_forked18_2_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to6_mul3722_0_NO_SHIFT_REG),
	.stall_out(local_bb2_mul3722_pop13_mul3722_fu_stall_out),
	.valid_in(local_bb2_mul3722_pop13_mul3722_inputs_ready),
	.valid_out(local_bb2_mul3722_pop13_mul3722_fu_valid_out),
	.stall_in(~(local_bb2_mul3722_pop13_mul3722_output_regs_ready)),
	.data_out(local_bb2_mul3722_pop13_mul3722_result),
	.feedback_in(feedback_data_in_13),
	.feedback_valid_in(feedback_valid_in_13),
	.feedback_stall_out(feedback_stall_out_13)
);

defparam local_bb2_mul3722_pop13_mul3722_feedback.COALESCE_DISTANCE = 1;
defparam local_bb2_mul3722_pop13_mul3722_feedback.DATA_WIDTH = 32;
defparam local_bb2_mul3722_pop13_mul3722_feedback.STYLE = "REGULAR";

assign local_bb2_mul3722_pop13_mul3722_inputs_ready = (rnode_1to6_mul3722_0_valid_out_NO_SHIFT_REG & rnode_1to6_forked18_0_valid_out_2_NO_SHIFT_REG);
assign local_bb2_mul3722_pop13_mul3722_output_regs_ready = ((~(local_bb2_mul3722_pop13_mul3722_valid_out_0_NO_SHIFT_REG) | ~(local_bb2_mul3722_pop13_mul3722_stall_in_0)) & (~(local_bb2_mul3722_pop13_mul3722_valid_out_1_NO_SHIFT_REG) | ~(local_bb2_mul3722_pop13_mul3722_stall_in_1)));
assign rnode_1to6_mul3722_0_stall_in_NO_SHIFT_REG = (local_bb2_mul3722_pop13_mul3722_fu_stall_out | ~(local_bb2_mul3722_pop13_mul3722_inputs_ready));
assign rnode_1to6_forked18_0_stall_in_2_NO_SHIFT_REG = (local_bb2_mul3722_pop13_mul3722_fu_stall_out | ~(local_bb2_mul3722_pop13_mul3722_inputs_ready));
assign local_bb2_mul3722_pop13_mul3722_causedstall = (local_bb2_mul3722_pop13_mul3722_inputs_ready && (local_bb2_mul3722_pop13_mul3722_fu_stall_out && !(~(local_bb2_mul3722_pop13_mul3722_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul3722_pop13_mul3722_NO_SHIFT_REG <= 'x;
		local_bb2_mul3722_pop13_mul3722_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul3722_pop13_mul3722_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul3722_pop13_mul3722_output_regs_ready)
		begin
			local_bb2_mul3722_pop13_mul3722_NO_SHIFT_REG <= local_bb2_mul3722_pop13_mul3722_result;
			local_bb2_mul3722_pop13_mul3722_valid_out_0_NO_SHIFT_REG <= local_bb2_mul3722_pop13_mul3722_fu_valid_out;
			local_bb2_mul3722_pop13_mul3722_valid_out_1_NO_SHIFT_REG <= local_bb2_mul3722_pop13_mul3722_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_mul3722_pop13_mul3722_stall_in_0))
			begin
				local_bb2_mul3722_pop13_mul3722_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul3722_pop13_mul3722_stall_in_1))
			begin
				local_bb2_mul3722_pop13_mul3722_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_notcmp1125_pop14_notcmp1125_inputs_ready;
 reg local_bb2_notcmp1125_pop14_notcmp1125_valid_out_0_NO_SHIFT_REG;
wire local_bb2_notcmp1125_pop14_notcmp1125_stall_in_0;
 reg local_bb2_notcmp1125_pop14_notcmp1125_valid_out_1_NO_SHIFT_REG;
wire local_bb2_notcmp1125_pop14_notcmp1125_stall_in_1;
wire local_bb2_notcmp1125_pop14_notcmp1125_output_regs_ready;
wire local_bb2_notcmp1125_pop14_notcmp1125_result;
wire local_bb2_notcmp1125_pop14_notcmp1125_fu_valid_out;
wire local_bb2_notcmp1125_pop14_notcmp1125_fu_stall_out;
 reg local_bb2_notcmp1125_pop14_notcmp1125_NO_SHIFT_REG;
wire local_bb2_notcmp1125_pop14_notcmp1125_causedstall;

acl_pop local_bb2_notcmp1125_pop14_notcmp1125_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to6_forked18_3_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to6_notcmp1125_0_NO_SHIFT_REG),
	.stall_out(local_bb2_notcmp1125_pop14_notcmp1125_fu_stall_out),
	.valid_in(local_bb2_notcmp1125_pop14_notcmp1125_inputs_ready),
	.valid_out(local_bb2_notcmp1125_pop14_notcmp1125_fu_valid_out),
	.stall_in(~(local_bb2_notcmp1125_pop14_notcmp1125_output_regs_ready)),
	.data_out(local_bb2_notcmp1125_pop14_notcmp1125_result),
	.feedback_in(feedback_data_in_14),
	.feedback_valid_in(feedback_valid_in_14),
	.feedback_stall_out(feedback_stall_out_14)
);

defparam local_bb2_notcmp1125_pop14_notcmp1125_feedback.COALESCE_DISTANCE = 1;
defparam local_bb2_notcmp1125_pop14_notcmp1125_feedback.DATA_WIDTH = 1;
defparam local_bb2_notcmp1125_pop14_notcmp1125_feedback.STYLE = "REGULAR";

assign local_bb2_notcmp1125_pop14_notcmp1125_inputs_ready = (rnode_1to6_notcmp1125_0_valid_out_NO_SHIFT_REG & rnode_1to6_forked18_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_notcmp1125_pop14_notcmp1125_output_regs_ready = ((~(local_bb2_notcmp1125_pop14_notcmp1125_valid_out_0_NO_SHIFT_REG) | ~(local_bb2_notcmp1125_pop14_notcmp1125_stall_in_0)) & (~(local_bb2_notcmp1125_pop14_notcmp1125_valid_out_1_NO_SHIFT_REG) | ~(local_bb2_notcmp1125_pop14_notcmp1125_stall_in_1)));
assign rnode_1to6_notcmp1125_0_stall_in_NO_SHIFT_REG = (local_bb2_notcmp1125_pop14_notcmp1125_fu_stall_out | ~(local_bb2_notcmp1125_pop14_notcmp1125_inputs_ready));
assign rnode_1to6_forked18_0_stall_in_3_NO_SHIFT_REG = (local_bb2_notcmp1125_pop14_notcmp1125_fu_stall_out | ~(local_bb2_notcmp1125_pop14_notcmp1125_inputs_ready));
assign local_bb2_notcmp1125_pop14_notcmp1125_causedstall = (local_bb2_notcmp1125_pop14_notcmp1125_inputs_ready && (local_bb2_notcmp1125_pop14_notcmp1125_fu_stall_out && !(~(local_bb2_notcmp1125_pop14_notcmp1125_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_notcmp1125_pop14_notcmp1125_NO_SHIFT_REG <= 'x;
		local_bb2_notcmp1125_pop14_notcmp1125_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_notcmp1125_pop14_notcmp1125_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_notcmp1125_pop14_notcmp1125_output_regs_ready)
		begin
			local_bb2_notcmp1125_pop14_notcmp1125_NO_SHIFT_REG <= local_bb2_notcmp1125_pop14_notcmp1125_result;
			local_bb2_notcmp1125_pop14_notcmp1125_valid_out_0_NO_SHIFT_REG <= local_bb2_notcmp1125_pop14_notcmp1125_fu_valid_out;
			local_bb2_notcmp1125_pop14_notcmp1125_valid_out_1_NO_SHIFT_REG <= local_bb2_notcmp1125_pop14_notcmp1125_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_notcmp1125_pop14_notcmp1125_stall_in_0))
			begin
				local_bb2_notcmp1125_pop14_notcmp1125_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_notcmp1125_pop14_notcmp1125_stall_in_1))
			begin
				local_bb2_notcmp1125_pop14_notcmp1125_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_notexitcond1428_pop15_notexitcond1428_inputs_ready;
 reg local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_0_NO_SHIFT_REG;
wire local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_0;
 reg local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_1_NO_SHIFT_REG;
wire local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_1;
wire local_bb2_notexitcond1428_pop15_notexitcond1428_output_regs_ready;
wire local_bb2_notexitcond1428_pop15_notexitcond1428_result;
wire local_bb2_notexitcond1428_pop15_notexitcond1428_fu_valid_out;
wire local_bb2_notexitcond1428_pop15_notexitcond1428_fu_stall_out;
 reg local_bb2_notexitcond1428_pop15_notexitcond1428_NO_SHIFT_REG;
wire local_bb2_notexitcond1428_pop15_notexitcond1428_causedstall;

acl_pop local_bb2_notexitcond1428_pop15_notexitcond1428_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to6_forked18_4_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to6_notexitcond1428_0_NO_SHIFT_REG),
	.stall_out(local_bb2_notexitcond1428_pop15_notexitcond1428_fu_stall_out),
	.valid_in(local_bb2_notexitcond1428_pop15_notexitcond1428_inputs_ready),
	.valid_out(local_bb2_notexitcond1428_pop15_notexitcond1428_fu_valid_out),
	.stall_in(~(local_bb2_notexitcond1428_pop15_notexitcond1428_output_regs_ready)),
	.data_out(local_bb2_notexitcond1428_pop15_notexitcond1428_result),
	.feedback_in(feedback_data_in_15),
	.feedback_valid_in(feedback_valid_in_15),
	.feedback_stall_out(feedback_stall_out_15)
);

defparam local_bb2_notexitcond1428_pop15_notexitcond1428_feedback.COALESCE_DISTANCE = 1;
defparam local_bb2_notexitcond1428_pop15_notexitcond1428_feedback.DATA_WIDTH = 1;
defparam local_bb2_notexitcond1428_pop15_notexitcond1428_feedback.STYLE = "REGULAR";

assign local_bb2_notexitcond1428_pop15_notexitcond1428_inputs_ready = (rnode_1to6_notexitcond1428_0_valid_out_NO_SHIFT_REG & rnode_1to6_forked18_0_valid_out_4_NO_SHIFT_REG);
assign local_bb2_notexitcond1428_pop15_notexitcond1428_output_regs_ready = ((~(local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_0_NO_SHIFT_REG) | ~(local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_0)) & (~(local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_1_NO_SHIFT_REG) | ~(local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_1)));
assign rnode_1to6_notexitcond1428_0_stall_in_NO_SHIFT_REG = (local_bb2_notexitcond1428_pop15_notexitcond1428_fu_stall_out | ~(local_bb2_notexitcond1428_pop15_notexitcond1428_inputs_ready));
assign rnode_1to6_forked18_0_stall_in_4_NO_SHIFT_REG = (local_bb2_notexitcond1428_pop15_notexitcond1428_fu_stall_out | ~(local_bb2_notexitcond1428_pop15_notexitcond1428_inputs_ready));
assign local_bb2_notexitcond1428_pop15_notexitcond1428_causedstall = (local_bb2_notexitcond1428_pop15_notexitcond1428_inputs_ready && (local_bb2_notexitcond1428_pop15_notexitcond1428_fu_stall_out && !(~(local_bb2_notexitcond1428_pop15_notexitcond1428_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_notexitcond1428_pop15_notexitcond1428_NO_SHIFT_REG <= 'x;
		local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_notexitcond1428_pop15_notexitcond1428_output_regs_ready)
		begin
			local_bb2_notexitcond1428_pop15_notexitcond1428_NO_SHIFT_REG <= local_bb2_notexitcond1428_pop15_notexitcond1428_result;
			local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_0_NO_SHIFT_REG <= local_bb2_notexitcond1428_pop15_notexitcond1428_fu_valid_out;
			local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_1_NO_SHIFT_REG <= local_bb2_notexitcond1428_pop15_notexitcond1428_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_0))
			begin
				local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_1))
			begin
				local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul6_inputs_ready;
 reg local_bb2_mul6_valid_out_NO_SHIFT_REG;
wire local_bb2_mul6_stall_in;
wire local_bb2_mul6_output_regs_ready;
wire [31:0] local_bb2_mul6;
 reg local_bb2_mul6_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul6_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul6_causedstall;

acl_int_mult int_module_local_bb2_mul6 (
	.clock(clock),
	.dataa((local_bb2_mul5 & 32'hFFFFFFFE)),
	.datab(input_inSize_x),
	.enable(local_bb2_mul6_output_regs_ready),
	.result(local_bb2_mul6)
);

defparam int_module_local_bb2_mul6.INPUT1_WIDTH = 32;
defparam int_module_local_bb2_mul6.INPUT2_WIDTH = 32;
defparam int_module_local_bb2_mul6.OUTPUT_WIDTH = 32;
defparam int_module_local_bb2_mul6.LATENCY = 3;
defparam int_module_local_bb2_mul6.SIGNED = 0;

assign local_bb2_mul6_inputs_ready = local_bb2_mul5_valid_out_0;
assign local_bb2_mul6_output_regs_ready = (&(~(local_bb2_mul6_valid_out_NO_SHIFT_REG) | ~(local_bb2_mul6_stall_in)));
assign local_bb2_mul5_stall_in_0 = (~(local_bb2_mul6_output_regs_ready) | ~(local_bb2_mul6_inputs_ready));
assign local_bb2_mul6_causedstall = (local_bb2_mul6_inputs_ready && (~(local_bb2_mul6_output_regs_ready) && !(~(local_bb2_mul6_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul6_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul6_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul6_output_regs_ready)
		begin
			local_bb2_mul6_valid_pipe_0_NO_SHIFT_REG <= local_bb2_mul6_inputs_ready;
			local_bb2_mul6_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul6_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul6_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul6_output_regs_ready)
		begin
			local_bb2_mul6_valid_out_NO_SHIFT_REG <= local_bb2_mul6_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb2_mul6_stall_in))
			begin
				local_bb2_mul6_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__u9_stall_local;
wire [31:0] local_bb2_var__u9;
wire [32:0] rci_rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3;

assign local_bb2_var__u9 = local_bb2_indvars_iv_next[31:0];
assign rci_rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3[31:0] = rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_1_NO_SHIFT_REG;
assign rci_rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3[32] = local_bb2_keep_going8_acl_pipeline_1_NO_SHIFT_REG;

// Register node:
//  * latency = 163
//  * capacity = 163
 logic rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_NO_SHIFT_REG;
 logic rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_NO_SHIFT_REG;
 logic [32:0] rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_NO_SHIFT_REG;
 logic rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic [32:0] rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_NO_SHIFT_REG;
 logic rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_3),
	.data_out(rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_NO_SHIFT_REG)
);

defparam rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_fifo.DEPTH = 164;
defparam rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_fifo.DATA_WIDTH = 33;
defparam rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_fifo.IMPL = "ram";

assign rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_inputs_ready_NO_SHIFT_REG = (rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_1_NO_SHIFT_REG & local_bb2_keep_going8_acl_pipeline_1_valid_out_NO_SHIFT_REG);
assign rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_1_NO_SHIFT_REG = rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_keep_going8_acl_pipeline_1_stall_in = rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_NO_SHIFT_REG = rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_reg_166_NO_SHIFT_REG;
assign rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_NO_SHIFT_REG;
assign rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_NO_SHIFT_REG = rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_memdep_phi1_or_valid_out;
wire local_bb2_memdep_phi1_or_stall_in;
wire local_bb2_memdep_phi1_or_inputs_ready;
wire local_bb2_memdep_phi1_or_stall_local;
wire local_bb2_memdep_phi1_or;
wire [34:0] rci_rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_7;

assign local_bb2_memdep_phi1_or_inputs_ready = (local_bb2_memdep_phi_pop11_acl_pop_i1_0_valid_out_NO_SHIFT_REG & local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_0_NO_SHIFT_REG);
assign local_bb2_memdep_phi1_or = (local_bb2_memdep_phi_pop11_acl_pop_i1_0_NO_SHIFT_REG | local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_NO_SHIFT_REG);
assign local_bb2_memdep_phi1_or_valid_out = local_bb2_memdep_phi1_or_inputs_ready;
assign local_bb2_memdep_phi1_or_stall_local = local_bb2_memdep_phi1_or_stall_in;
assign local_bb2_memdep_phi_pop11_acl_pop_i1_0_stall_in = (local_bb2_memdep_phi1_or_stall_local | ~(local_bb2_memdep_phi1_or_inputs_ready));
assign local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_0 = (local_bb2_memdep_phi1_or_stall_local | ~(local_bb2_memdep_phi1_or_inputs_ready));
assign rci_rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_7[0] = local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_NO_SHIFT_REG;
assign rci_rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_7[32:1] = local_bb2_mul3722_pop13_mul3722_NO_SHIFT_REG;
assign rci_rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_7[33] = local_bb2_notcmp1125_pop14_notcmp1125_NO_SHIFT_REG;
assign rci_rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_7[34] = local_bb2_notexitcond1428_pop15_notexitcond1428_NO_SHIFT_REG;

// Register node:
//  * latency = 159
//  * capacity = 159
 logic rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_valid_out_NO_SHIFT_REG;
 logic rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_in_NO_SHIFT_REG;
 logic [34:0] rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_NO_SHIFT_REG;
 logic rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic [34:0] rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_NO_SHIFT_REG;
 logic rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_7),
	.data_out(rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_NO_SHIFT_REG)
);

defparam rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_fifo.DEPTH = 160;
defparam rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_fifo.DATA_WIDTH = 35;
defparam rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_fifo.IMPL = "ram";

assign rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_inputs_ready_NO_SHIFT_REG = (local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_2_NO_SHIFT_REG & local_bb2_mul3722_pop13_mul3722_valid_out_1_NO_SHIFT_REG & local_bb2_notcmp1125_pop14_notcmp1125_valid_out_1_NO_SHIFT_REG & local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_1_NO_SHIFT_REG);
assign rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_2 = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_mul3722_pop13_mul3722_stall_in_1 = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_notcmp1125_pop14_notcmp1125_stall_in_1 = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_1 = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_NO_SHIFT_REG = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_reg_166_NO_SHIFT_REG;
assign rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_in_NO_SHIFT_REG;
assign rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_valid_out_NO_SHIFT_REG = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_valid_out_reg_166_NO_SHIFT_REG;

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_5to5_bb2_mul6_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to5_bb2_mul6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to5_bb2_mul6_0_NO_SHIFT_REG;
 logic rnode_5to5_bb2_mul6_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to5_bb2_mul6_0_reg_5_NO_SHIFT_REG;
 logic rnode_5to5_bb2_mul6_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_5to5_bb2_mul6_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_5to5_bb2_mul6_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_5to5_bb2_mul6_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to5_bb2_mul6_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to5_bb2_mul6_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_5to5_bb2_mul6_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_5to5_bb2_mul6_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in((local_bb2_mul6 & 32'hFFFFFFFE)),
	.data_out(rnode_5to5_bb2_mul6_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_5to5_bb2_mul6_0_reg_5_fifo.DEPTH = 3;
defparam rnode_5to5_bb2_mul6_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_5to5_bb2_mul6_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_5to5_bb2_mul6_0_reg_5_fifo.IMPL = "zl_reg";

assign rnode_5to5_bb2_mul6_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb2_mul6_valid_out_NO_SHIFT_REG;
assign local_bb2_mul6_stall_in = rnode_5to5_bb2_mul6_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_5to5_bb2_mul6_0_NO_SHIFT_REG = rnode_5to5_bb2_mul6_0_reg_5_NO_SHIFT_REG;
assign rnode_5to5_bb2_mul6_0_stall_in_reg_5_NO_SHIFT_REG = rnode_5to5_bb2_mul6_0_stall_in_NO_SHIFT_REG;
assign rnode_5to5_bb2_mul6_0_valid_out_NO_SHIFT_REG = rnode_5to5_bb2_mul6_0_valid_out_reg_5_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp3_stall_local;
wire [32:0] cmprep_local_bb2_cmp3;
wire local_bb2_cmp3;

assign cmprep_local_bb2_cmp3 = (local_bb2_var__u9 - (input_wii_div & 32'h7FFFFFFF));
assign local_bb2_cmp3 = cmprep_local_bb2_cmp3[32];

// This section implements a staging register.
// 
wire rstag_7to7_bb2_memdep_phi1_or_valid_out_0;
wire rstag_7to7_bb2_memdep_phi1_or_stall_in_0;
wire rstag_7to7_bb2_memdep_phi1_or_valid_out_1;
wire rstag_7to7_bb2_memdep_phi1_or_stall_in_1;
wire rstag_7to7_bb2_memdep_phi1_or_inputs_ready;
wire rstag_7to7_bb2_memdep_phi1_or_stall_local;
 reg rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG;
wire rstag_7to7_bb2_memdep_phi1_or_combined_valid;
 reg rstag_7to7_bb2_memdep_phi1_or_staging_reg_NO_SHIFT_REG;
wire rstag_7to7_bb2_memdep_phi1_or;
 reg rstag_7to7_bb2_memdep_phi1_or_consumed_0_NO_SHIFT_REG;
 reg rstag_7to7_bb2_memdep_phi1_or_consumed_1_NO_SHIFT_REG;

assign rstag_7to7_bb2_memdep_phi1_or_inputs_ready = local_bb2_memdep_phi1_or_valid_out;
assign rstag_7to7_bb2_memdep_phi1_or = (rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG ? rstag_7to7_bb2_memdep_phi1_or_staging_reg_NO_SHIFT_REG : local_bb2_memdep_phi1_or);
assign rstag_7to7_bb2_memdep_phi1_or_combined_valid = (rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG | rstag_7to7_bb2_memdep_phi1_or_inputs_ready);
assign rstag_7to7_bb2_memdep_phi1_or_stall_local = ((rstag_7to7_bb2_memdep_phi1_or_stall_in_0 & ~(rstag_7to7_bb2_memdep_phi1_or_consumed_0_NO_SHIFT_REG)) | (rstag_7to7_bb2_memdep_phi1_or_stall_in_1 & ~(rstag_7to7_bb2_memdep_phi1_or_consumed_1_NO_SHIFT_REG)));
assign rstag_7to7_bb2_memdep_phi1_or_valid_out_0 = (rstag_7to7_bb2_memdep_phi1_or_combined_valid & ~(rstag_7to7_bb2_memdep_phi1_or_consumed_0_NO_SHIFT_REG));
assign rstag_7to7_bb2_memdep_phi1_or_valid_out_1 = (rstag_7to7_bb2_memdep_phi1_or_combined_valid & ~(rstag_7to7_bb2_memdep_phi1_or_consumed_1_NO_SHIFT_REG));
assign local_bb2_memdep_phi1_or_stall_in = (|rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb2_memdep_phi1_or_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_7to7_bb2_memdep_phi1_or_stall_local)
		begin
			if (~(rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG))
			begin
				rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG <= rstag_7to7_bb2_memdep_phi1_or_inputs_ready;
			end
		end
		else
		begin
			rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_7to7_bb2_memdep_phi1_or_staging_valid_NO_SHIFT_REG))
		begin
			rstag_7to7_bb2_memdep_phi1_or_staging_reg_NO_SHIFT_REG <= local_bb2_memdep_phi1_or;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb2_memdep_phi1_or_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb2_memdep_phi1_or_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_7to7_bb2_memdep_phi1_or_consumed_0_NO_SHIFT_REG <= (rstag_7to7_bb2_memdep_phi1_or_combined_valid & (rstag_7to7_bb2_memdep_phi1_or_consumed_0_NO_SHIFT_REG | ~(rstag_7to7_bb2_memdep_phi1_or_stall_in_0)) & rstag_7to7_bb2_memdep_phi1_or_stall_local);
		rstag_7to7_bb2_memdep_phi1_or_consumed_1_NO_SHIFT_REG <= (rstag_7to7_bb2_memdep_phi1_or_combined_valid & (rstag_7to7_bb2_memdep_phi1_or_consumed_1_NO_SHIFT_REG | ~(rstag_7to7_bb2_memdep_phi1_or_stall_in_1)) & rstag_7to7_bb2_memdep_phi1_or_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__u10_stall_local;
wire local_bb2_var__u10;

assign local_bb2_var__u10 = (local_bb2_cmp3 & input_wii_var__u7);

// This section implements an unregistered operation.
// 
wire local_bb2_indvars_iv_pop10_acl_pop_i64_0_valid_out_1;
wire local_bb2_indvars_iv_pop10_acl_pop_i64_0_stall_in_1;
wire local_bb2_indvars_iv_next_valid_out_1;
wire local_bb2_indvars_iv_next_stall_in_1;
wire local_bb2_var__u10_valid_out;
wire local_bb2_var__u10_stall_in;
wire local_bb2_cmp3_not_valid_out;
wire local_bb2_cmp3_not_stall_in;
wire local_bb2_cmp3_not_inputs_ready;
wire local_bb2_cmp3_not_stall_local;
wire local_bb2_cmp3_not;
wire local_bb2_cmp3_not_stall_out_local_or;
wire local_bb2_cmp3_not_stall_local_fanout;
wire local_bb2_cmp3_not_fu_valid_out_and;
 reg local_bb2_indvars_iv_pop10_acl_pop_i64_0_consumed_1_NO_SHIFT_REG;
 reg local_bb2_indvars_iv_next_consumed_1_NO_SHIFT_REG;
 reg local_bb2_var__u10_consumed_0_NO_SHIFT_REG;
 reg local_bb2_cmp3_not_consumed_0_NO_SHIFT_REG;

assign local_bb2_cmp3_not_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb2_indvars_iv_pop10_acl_pop_i64_0_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb2_cmp3_not = (local_bb2_cmp3 ^ 1'b1);
assign local_bb2_cmp3_not_stall_out_local_or = local_bb2_indvars_iv_pop10_acl_pop_i64_0_fu_stall_out;
assign local_bb2_indvars_iv_pop10_acl_pop_i64_0_stall_local = local_bb2_cmp3_not_stall_local_fanout;
assign local_bb2_cmp3_not_fu_valid_out_and = local_bb2_indvars_iv_pop10_acl_pop_i64_0_fu_valid_out;
assign local_bb2_cmp3_not_stall_local_fanout = ((local_bb2_indvars_iv_pop10_acl_pop_i64_0_stall_in_1 & ~(local_bb2_indvars_iv_pop10_acl_pop_i64_0_consumed_1_NO_SHIFT_REG)) | (local_bb2_indvars_iv_next_stall_in_1 & ~(local_bb2_indvars_iv_next_consumed_1_NO_SHIFT_REG)) | (local_bb2_var__u10_stall_in & ~(local_bb2_var__u10_consumed_0_NO_SHIFT_REG)) | (local_bb2_cmp3_not_stall_in & ~(local_bb2_cmp3_not_consumed_0_NO_SHIFT_REG)));
assign local_bb2_indvars_iv_pop10_acl_pop_i64_0_valid_out_1 = (local_bb2_cmp3_not_fu_valid_out_and & ~(local_bb2_indvars_iv_pop10_acl_pop_i64_0_consumed_1_NO_SHIFT_REG));
assign local_bb2_indvars_iv_next_valid_out_1 = (local_bb2_cmp3_not_fu_valid_out_and & ~(local_bb2_indvars_iv_next_consumed_1_NO_SHIFT_REG));
assign local_bb2_var__u10_valid_out = (local_bb2_cmp3_not_fu_valid_out_and & ~(local_bb2_var__u10_consumed_0_NO_SHIFT_REG));
assign local_bb2_cmp3_not_valid_out = (local_bb2_cmp3_not_fu_valid_out_and & ~(local_bb2_cmp3_not_consumed_0_NO_SHIFT_REG));
assign merge_node_stall_in_1 = (|local_bb2_cmp3_not_stall_out_local_or);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_indvars_iv_pop10_acl_pop_i64_0_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_indvars_iv_next_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u10_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp3_not_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_indvars_iv_pop10_acl_pop_i64_0_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp3_not_fu_valid_out_and & (local_bb2_indvars_iv_pop10_acl_pop_i64_0_consumed_1_NO_SHIFT_REG | ~(local_bb2_indvars_iv_pop10_acl_pop_i64_0_stall_in_1)) & local_bb2_cmp3_not_stall_local_fanout);
		local_bb2_indvars_iv_next_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp3_not_fu_valid_out_and & (local_bb2_indvars_iv_next_consumed_1_NO_SHIFT_REG | ~(local_bb2_indvars_iv_next_stall_in_1)) & local_bb2_cmp3_not_stall_local_fanout);
		local_bb2_var__u10_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp3_not_fu_valid_out_and & (local_bb2_var__u10_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u10_stall_in)) & local_bb2_cmp3_not_stall_local_fanout);
		local_bb2_cmp3_not_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp3_not_fu_valid_out_and & (local_bb2_cmp3_not_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp3_not_stall_in)) & local_bb2_cmp3_not_stall_local_fanout);
	end
end


// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_NO_SHIFT_REG;
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_1_NO_SHIFT_REG;
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_reg_5_NO_SHIFT_REG;
 reg rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb2_indvars_iv_pop10_acl_pop_i64_0),
	.data_out(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_fifo.DEPTH = 5;
defparam rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_fifo.DATA_WIDTH = 64;
defparam rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb2_indvars_iv_pop10_acl_pop_i64_0_valid_out_1;
assign local_bb2_indvars_iv_pop10_acl_pop_i64_0_stall_in_1 = rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_reg_5_NO_SHIFT_REG = ((rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_NO_SHIFT_REG = (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_reg_5_NO_SHIFT_REG & ~(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_1_NO_SHIFT_REG = (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_reg_5_NO_SHIFT_REG & ~(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_NO_SHIFT_REG = rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_NO_SHIFT_REG;
assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_1_NO_SHIFT_REG = rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_0_NO_SHIFT_REG <= (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_reg_5_NO_SHIFT_REG & (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_reg_5_NO_SHIFT_REG);
		rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_1_NO_SHIFT_REG <= (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_reg_5_NO_SHIFT_REG & (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_reg_5_NO_SHIFT_REG);
	end
end


// This section implements a staging register.
// 
wire rstag_1to1_bb2_var__u10_valid_out_0;
wire rstag_1to1_bb2_var__u10_stall_in_0;
wire rstag_1to1_bb2_var__u10_valid_out_1;
wire rstag_1to1_bb2_var__u10_stall_in_1;
wire rstag_1to1_bb2_var__u10_inputs_ready;
wire rstag_1to1_bb2_var__u10_stall_local;
 reg rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG;
wire rstag_1to1_bb2_var__u10_combined_valid;
 reg rstag_1to1_bb2_var__u10_staging_reg_NO_SHIFT_REG;
wire rstag_1to1_bb2_var__u10;
 reg rstag_1to1_bb2_var__u10_consumed_0_NO_SHIFT_REG;
 reg rstag_1to1_bb2_var__u10_consumed_1_NO_SHIFT_REG;

assign rstag_1to1_bb2_var__u10_inputs_ready = local_bb2_var__u10_valid_out;
assign rstag_1to1_bb2_var__u10 = (rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG ? rstag_1to1_bb2_var__u10_staging_reg_NO_SHIFT_REG : local_bb2_var__u10);
assign rstag_1to1_bb2_var__u10_combined_valid = (rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG | rstag_1to1_bb2_var__u10_inputs_ready);
assign rstag_1to1_bb2_var__u10_stall_local = ((rstag_1to1_bb2_var__u10_stall_in_0 & ~(rstag_1to1_bb2_var__u10_consumed_0_NO_SHIFT_REG)) | (rstag_1to1_bb2_var__u10_stall_in_1 & ~(rstag_1to1_bb2_var__u10_consumed_1_NO_SHIFT_REG)));
assign rstag_1to1_bb2_var__u10_valid_out_0 = (rstag_1to1_bb2_var__u10_combined_valid & ~(rstag_1to1_bb2_var__u10_consumed_0_NO_SHIFT_REG));
assign rstag_1to1_bb2_var__u10_valid_out_1 = (rstag_1to1_bb2_var__u10_combined_valid & ~(rstag_1to1_bb2_var__u10_consumed_1_NO_SHIFT_REG));
assign local_bb2_var__u10_stall_in = (|rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_1to1_bb2_var__u10_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_1to1_bb2_var__u10_stall_local)
		begin
			if (~(rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG))
			begin
				rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG <= rstag_1to1_bb2_var__u10_inputs_ready;
			end
		end
		else
		begin
			rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_1to1_bb2_var__u10_staging_valid_NO_SHIFT_REG))
		begin
			rstag_1to1_bb2_var__u10_staging_reg_NO_SHIFT_REG <= local_bb2_var__u10;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_1to1_bb2_var__u10_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_1to1_bb2_var__u10_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_1to1_bb2_var__u10_consumed_0_NO_SHIFT_REG <= (rstag_1to1_bb2_var__u10_combined_valid & (rstag_1to1_bb2_var__u10_consumed_0_NO_SHIFT_REG | ~(rstag_1to1_bb2_var__u10_stall_in_0)) & rstag_1to1_bb2_var__u10_stall_local);
		rstag_1to1_bb2_var__u10_consumed_1_NO_SHIFT_REG <= (rstag_1to1_bb2_var__u10_combined_valid & (rstag_1to1_bb2_var__u10_consumed_1_NO_SHIFT_REG | ~(rstag_1to1_bb2_var__u10_stall_in_1)) & rstag_1to1_bb2_var__u10_stall_local);
	end
end


// Register node:
//  * latency = 165
//  * capacity = 165
 logic rnode_1to166_bb2_cmp3_not_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to166_bb2_cmp3_not_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to166_bb2_cmp3_not_0_NO_SHIFT_REG;
 logic rnode_1to166_bb2_cmp3_not_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to166_bb2_cmp3_not_0_reg_166_NO_SHIFT_REG;
 logic rnode_1to166_bb2_cmp3_not_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rnode_1to166_bb2_cmp3_not_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rnode_1to166_bb2_cmp3_not_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_1to166_bb2_cmp3_not_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to166_bb2_cmp3_not_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to166_bb2_cmp3_not_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_1to166_bb2_cmp3_not_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_1to166_bb2_cmp3_not_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(local_bb2_cmp3_not),
	.data_out(rnode_1to166_bb2_cmp3_not_0_reg_166_NO_SHIFT_REG)
);

defparam rnode_1to166_bb2_cmp3_not_0_reg_166_fifo.DEPTH = 166;
defparam rnode_1to166_bb2_cmp3_not_0_reg_166_fifo.DATA_WIDTH = 1;
defparam rnode_1to166_bb2_cmp3_not_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to166_bb2_cmp3_not_0_reg_166_fifo.IMPL = "ram";

assign rnode_1to166_bb2_cmp3_not_0_reg_166_inputs_ready_NO_SHIFT_REG = local_bb2_cmp3_not_valid_out;
assign local_bb2_cmp3_not_stall_in = rnode_1to166_bb2_cmp3_not_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_1to166_bb2_cmp3_not_0_NO_SHIFT_REG = rnode_1to166_bb2_cmp3_not_0_reg_166_NO_SHIFT_REG;
assign rnode_1to166_bb2_cmp3_not_0_stall_in_reg_166_NO_SHIFT_REG = rnode_1to166_bb2_cmp3_not_0_stall_in_NO_SHIFT_REG;
assign rnode_1to166_bb2_cmp3_not_0_valid_out_NO_SHIFT_REG = rnode_1to166_bb2_cmp3_not_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u11_stall_local;
wire [63:0] local_bb2_var__u11;

assign local_bb2_var__u11 = (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_NO_SHIFT_REG << 64'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb2_var__u10_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u10_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u10_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u10_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u10_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u10_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u10_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__u10_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb2_var__u10_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb2_var__u10_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb2_var__u10_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb2_var__u10_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb2_var__u10_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(rstag_1to1_bb2_var__u10),
	.data_out(rnode_1to2_bb2_var__u10_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb2_var__u10_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb2_var__u10_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb2_var__u10_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb2_var__u10_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb2_var__u10_0_reg_2_inputs_ready_NO_SHIFT_REG = rstag_1to1_bb2_var__u10_valid_out_0;
assign rstag_1to1_bb2_var__u10_stall_in_0 = rnode_1to2_bb2_var__u10_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u10_0_NO_SHIFT_REG = rnode_1to2_bb2_var__u10_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u10_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb2_var__u10_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__u10_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb2_var__u10_0_valid_out_reg_2_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb2_indvars_iv_push10_indvars_iv_next_inputs_ready;
 reg local_bb2_indvars_iv_push10_indvars_iv_next_valid_out_NO_SHIFT_REG;
wire local_bb2_indvars_iv_push10_indvars_iv_next_stall_in;
wire local_bb2_indvars_iv_push10_indvars_iv_next_output_regs_ready;
wire [63:0] local_bb2_indvars_iv_push10_indvars_iv_next_result;
wire local_bb2_indvars_iv_push10_indvars_iv_next_fu_valid_out;
wire local_bb2_indvars_iv_push10_indvars_iv_next_fu_stall_out;
 reg [63:0] local_bb2_indvars_iv_push10_indvars_iv_next_NO_SHIFT_REG;
wire local_bb2_indvars_iv_push10_indvars_iv_next_causedstall;

acl_push local_bb2_indvars_iv_push10_indvars_iv_next_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rstag_1to1_bb2_var__u10),
	.predicate(1'b0),
	.data_in(local_bb2_indvars_iv_next),
	.stall_out(local_bb2_indvars_iv_push10_indvars_iv_next_fu_stall_out),
	.valid_in(local_bb2_indvars_iv_push10_indvars_iv_next_inputs_ready),
	.valid_out(local_bb2_indvars_iv_push10_indvars_iv_next_fu_valid_out),
	.stall_in(~(local_bb2_indvars_iv_push10_indvars_iv_next_output_regs_ready)),
	.data_out(local_bb2_indvars_iv_push10_indvars_iv_next_result),
	.feedback_out(feedback_data_out_10),
	.feedback_valid_out(feedback_valid_out_10),
	.feedback_stall_in(feedback_stall_in_10)
);

defparam local_bb2_indvars_iv_push10_indvars_iv_next_feedback.STALLFREE = 0;
defparam local_bb2_indvars_iv_push10_indvars_iv_next_feedback.DATA_WIDTH = 64;
defparam local_bb2_indvars_iv_push10_indvars_iv_next_feedback.FIFO_DEPTH = 4;
defparam local_bb2_indvars_iv_push10_indvars_iv_next_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb2_indvars_iv_push10_indvars_iv_next_feedback.STYLE = "REGULAR";

assign local_bb2_indvars_iv_push10_indvars_iv_next_inputs_ready = (local_bb2_indvars_iv_next_valid_out_1 & rstag_1to1_bb2_var__u10_valid_out_1);
assign local_bb2_indvars_iv_push10_indvars_iv_next_output_regs_ready = (&(~(local_bb2_indvars_iv_push10_indvars_iv_next_valid_out_NO_SHIFT_REG) | ~(local_bb2_indvars_iv_push10_indvars_iv_next_stall_in)));
assign local_bb2_indvars_iv_next_stall_in_1 = (local_bb2_indvars_iv_push10_indvars_iv_next_fu_stall_out | ~(local_bb2_indvars_iv_push10_indvars_iv_next_inputs_ready));
assign rstag_1to1_bb2_var__u10_stall_in_1 = (local_bb2_indvars_iv_push10_indvars_iv_next_fu_stall_out | ~(local_bb2_indvars_iv_push10_indvars_iv_next_inputs_ready));
assign local_bb2_indvars_iv_push10_indvars_iv_next_causedstall = (local_bb2_indvars_iv_push10_indvars_iv_next_inputs_ready && (local_bb2_indvars_iv_push10_indvars_iv_next_fu_stall_out && !(~(local_bb2_indvars_iv_push10_indvars_iv_next_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_indvars_iv_push10_indvars_iv_next_NO_SHIFT_REG <= 'x;
		local_bb2_indvars_iv_push10_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_indvars_iv_push10_indvars_iv_next_output_regs_ready)
		begin
			local_bb2_indvars_iv_push10_indvars_iv_next_NO_SHIFT_REG <= local_bb2_indvars_iv_push10_indvars_iv_next_result;
			local_bb2_indvars_iv_push10_indvars_iv_next_valid_out_NO_SHIFT_REG <= local_bb2_indvars_iv_push10_indvars_iv_next_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_indvars_iv_push10_indvars_iv_next_stall_in))
			begin
				local_bb2_indvars_iv_push10_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_cmp3_not_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_cmp3_not_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_cmp3_not_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_cmp3_not_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_cmp3_not_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_cmp3_not_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_cmp3_not_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_cmp3_not_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_cmp3_not_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_cmp3_not_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_cmp3_not_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_cmp3_not_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_cmp3_not_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(rnode_1to166_bb2_cmp3_not_0_NO_SHIFT_REG),
	.data_out(rnode_166to167_bb2_cmp3_not_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_cmp3_not_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_cmp3_not_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_cmp3_not_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_cmp3_not_0_reg_167_fifo.IMPL = "ll_reg";

assign rnode_166to167_bb2_cmp3_not_0_reg_167_inputs_ready_NO_SHIFT_REG = rnode_1to166_bb2_cmp3_not_0_valid_out_NO_SHIFT_REG;
assign rnode_1to166_bb2_cmp3_not_0_stall_in_NO_SHIFT_REG = rnode_166to167_bb2_cmp3_not_0_stall_out_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_cmp3_not_0_NO_SHIFT_REG = rnode_166to167_bb2_cmp3_not_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_cmp3_not_0_stall_in_reg_167_NO_SHIFT_REG = rnode_166to167_bb2_cmp3_not_0_stall_in_NO_SHIFT_REG;
assign rnode_166to167_bb2_cmp3_not_0_valid_out_NO_SHIFT_REG = rnode_166to167_bb2_cmp3_not_0_valid_out_reg_167_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_var__stall_local;
wire [31:0] local_bb2_var_;
wire [63:0] local_bb2_var_$ps;

assign local_bb2_var_$ps = (local_bb2_var__u11 & 64'hFFFFFFFFFFFFFFFE);
assign local_bb2_var_ = local_bb2_var_$ps[31:0];

// This section implements a registered operation.
// 
wire local_bb2_notexitcond9__inputs_ready;
 reg local_bb2_notexitcond9__valid_out_0_NO_SHIFT_REG;
wire local_bb2_notexitcond9__stall_in_0;
 reg local_bb2_notexitcond9__valid_out_1_NO_SHIFT_REG;
wire local_bb2_notexitcond9__stall_in_1;
wire local_bb2_notexitcond9__output_regs_ready;
wire local_bb2_notexitcond9__result;
wire local_bb2_notexitcond9__fu_valid_out;
wire local_bb2_notexitcond9__fu_stall_out;
 reg local_bb2_notexitcond9__NO_SHIFT_REG;
wire local_bb2_notexitcond9__causedstall;
wire [95:0] rci_rcnode_2to166_rc1_bb2_mul5_0_reg_2;

acl_push local_bb2_notexitcond9__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(rnode_1to2_bb2_var__u10_0_NO_SHIFT_REG),
	.stall_out(local_bb2_notexitcond9__fu_stall_out),
	.valid_in(local_bb2_notexitcond9__inputs_ready),
	.valid_out(local_bb2_notexitcond9__fu_valid_out),
	.stall_in(~(local_bb2_notexitcond9__output_regs_ready)),
	.data_out(local_bb2_notexitcond9__result),
	.feedback_out(feedback_data_out_5),
	.feedback_valid_out(feedback_valid_out_5),
	.feedback_stall_in(feedback_stall_in_5)
);

defparam local_bb2_notexitcond9__feedback.STALLFREE = 0;
defparam local_bb2_notexitcond9__feedback.DATA_WIDTH = 1;
defparam local_bb2_notexitcond9__feedback.FIFO_DEPTH = 2;
defparam local_bb2_notexitcond9__feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb2_notexitcond9__feedback.STYLE = "REGULAR";

assign local_bb2_notexitcond9__inputs_ready = rnode_1to2_bb2_var__u10_0_valid_out_NO_SHIFT_REG;
assign local_bb2_notexitcond9__output_regs_ready = ((~(local_bb2_notexitcond9__valid_out_0_NO_SHIFT_REG) | ~(local_bb2_notexitcond9__stall_in_0)) & (~(local_bb2_notexitcond9__valid_out_1_NO_SHIFT_REG) | ~(local_bb2_notexitcond9__stall_in_1)));
assign rnode_1to2_bb2_var__u10_0_stall_in_NO_SHIFT_REG = (local_bb2_notexitcond9__fu_stall_out | ~(local_bb2_notexitcond9__inputs_ready));
assign local_bb2_notexitcond9__causedstall = (local_bb2_notexitcond9__inputs_ready && (local_bb2_notexitcond9__fu_stall_out && !(~(local_bb2_notexitcond9__output_regs_ready))));
assign rci_rcnode_2to166_rc1_bb2_mul5_0_reg_2[31:0] = (local_bb2_mul5 & 32'hFFFFFFFE);
assign rci_rcnode_2to166_rc1_bb2_mul5_0_reg_2[95:32] = local_bb2_indvars_iv_push10_indvars_iv_next_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_notexitcond9__NO_SHIFT_REG <= 'x;
		local_bb2_notexitcond9__valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_notexitcond9__valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_notexitcond9__output_regs_ready)
		begin
			local_bb2_notexitcond9__NO_SHIFT_REG <= local_bb2_notexitcond9__result;
			local_bb2_notexitcond9__valid_out_0_NO_SHIFT_REG <= local_bb2_notexitcond9__fu_valid_out;
			local_bb2_notexitcond9__valid_out_1_NO_SHIFT_REG <= local_bb2_notexitcond9__fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_notexitcond9__stall_in_0))
			begin
				local_bb2_notexitcond9__valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_notexitcond9__stall_in_1))
			begin
				local_bb2_notexitcond9__valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 164
//  * capacity = 164
 logic rcnode_2to166_rc1_bb2_mul5_0_valid_out_NO_SHIFT_REG;
 logic rcnode_2to166_rc1_bb2_mul5_0_stall_in_NO_SHIFT_REG;
 logic [95:0] rcnode_2to166_rc1_bb2_mul5_0_NO_SHIFT_REG;
 logic rcnode_2to166_rc1_bb2_mul5_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic [95:0] rcnode_2to166_rc1_bb2_mul5_0_reg_166_NO_SHIFT_REG;
 logic rcnode_2to166_rc1_bb2_mul5_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_2to166_rc1_bb2_mul5_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_2to166_rc1_bb2_mul5_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_2to166_rc1_bb2_mul5_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_2to166_rc1_bb2_mul5_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_2to166_rc1_bb2_mul5_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_2to166_rc1_bb2_mul5_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_2to166_rc1_bb2_mul5_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_2to166_rc1_bb2_mul5_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_2to166_rc1_bb2_mul5_0_reg_2),
	.data_out(rcnode_2to166_rc1_bb2_mul5_0_reg_166_NO_SHIFT_REG)
);

defparam rcnode_2to166_rc1_bb2_mul5_0_reg_166_fifo.DEPTH = 165;
defparam rcnode_2to166_rc1_bb2_mul5_0_reg_166_fifo.DATA_WIDTH = 96;
defparam rcnode_2to166_rc1_bb2_mul5_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_2to166_rc1_bb2_mul5_0_reg_166_fifo.IMPL = "ram";

assign rcnode_2to166_rc1_bb2_mul5_0_reg_166_inputs_ready_NO_SHIFT_REG = (local_bb2_mul5_valid_out_1 & local_bb2_indvars_iv_push10_indvars_iv_next_valid_out_NO_SHIFT_REG);
assign rcnode_2to166_rc1_bb2_mul5_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_2to166_rc1_bb2_mul5_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_2to166_rc1_bb2_mul5_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign local_bb2_mul5_stall_in_1 = rcnode_2to166_rc1_bb2_mul5_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_indvars_iv_push10_indvars_iv_next_stall_in = rcnode_2to166_rc1_bb2_mul5_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_2to166_rc1_bb2_mul5_0_NO_SHIFT_REG = rcnode_2to166_rc1_bb2_mul5_0_reg_166_NO_SHIFT_REG;
assign rcnode_2to166_rc1_bb2_mul5_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_2to166_rc1_bb2_mul5_0_stall_in_NO_SHIFT_REG;
assign rcnode_2to166_rc1_bb2_mul5_0_valid_out_NO_SHIFT_REG = rcnode_2to166_rc1_bb2_mul5_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_notcmp_valid_out;
wire local_bb2_notcmp_stall_in;
wire local_bb2_notcmp_inputs_ready;
wire local_bb2_notcmp_stall_local;
wire local_bb2_notcmp;

assign local_bb2_notcmp_inputs_ready = rnode_166to167_bb2_cmp3_not_0_valid_out_NO_SHIFT_REG;
assign local_bb2_notcmp = (input_wii_var_ | rnode_166to167_bb2_cmp3_not_0_NO_SHIFT_REG);
assign local_bb2_notcmp_valid_out = local_bb2_notcmp_inputs_ready;
assign local_bb2_notcmp_stall_local = local_bb2_notcmp_stall_in;
assign rnode_166to167_bb2_cmp3_not_0_stall_in_NO_SHIFT_REG = (|local_bb2_notcmp_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb2_var__valid_out_1;
wire local_bb2_var__stall_in_1;
wire local_bb2_add_valid_out;
wire local_bb2_add_stall_in;
wire local_bb2_add_inputs_ready;
wire local_bb2_add_stall_local;
wire [31:0] local_bb2_add;
 reg local_bb2_var__consumed_1_NO_SHIFT_REG;
 reg local_bb2_add_consumed_0_NO_SHIFT_REG;

assign local_bb2_add_inputs_ready = (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_0_NO_SHIFT_REG & rnode_5to5_bb2_mul6_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add = ((local_bb2_var_ & 32'hFFFFFFFE) + (rnode_5to5_bb2_mul6_0_NO_SHIFT_REG & 32'hFFFFFFFE));
assign local_bb2_add_stall_local = ((local_bb2_var__stall_in_1 & ~(local_bb2_var__consumed_1_NO_SHIFT_REG)) | (local_bb2_add_stall_in & ~(local_bb2_add_consumed_0_NO_SHIFT_REG)));
assign local_bb2_var__valid_out_1 = (local_bb2_add_inputs_ready & ~(local_bb2_var__consumed_1_NO_SHIFT_REG));
assign local_bb2_add_valid_out = (local_bb2_add_inputs_ready & ~(local_bb2_add_consumed_0_NO_SHIFT_REG));
assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_0_NO_SHIFT_REG = (local_bb2_add_stall_local | ~(local_bb2_add_inputs_ready));
assign rnode_5to5_bb2_mul6_0_stall_in_NO_SHIFT_REG = (local_bb2_add_stall_local | ~(local_bb2_add_inputs_ready));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_var__consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_var__consumed_1_NO_SHIFT_REG <= (local_bb2_add_inputs_ready & (local_bb2_var__consumed_1_NO_SHIFT_REG | ~(local_bb2_var__stall_in_1)) & local_bb2_add_stall_local);
		local_bb2_add_consumed_0_NO_SHIFT_REG <= (local_bb2_add_inputs_ready & (local_bb2_add_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_stall_in)) & local_bb2_add_stall_local);
	end
end


// This section implements a registered operation.
// 
wire local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_inputs_ready;
 reg local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_valid_out_NO_SHIFT_REG;
wire local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_stall_in;
wire local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_output_regs_ready;
wire [31:0] local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_result;
wire local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_valid_out;
wire local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_stall_out;
 reg [31:0] local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_NO_SHIFT_REG;
wire local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_causedstall;

acl_push local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb2_notexitcond9__NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_NO_SHIFT_REG),
	.stall_out(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_stall_out),
	.valid_in(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_inputs_ready),
	.valid_out(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_valid_out),
	.stall_in(~(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_output_regs_ready)),
	.data_out(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_result),
	.feedback_out(feedback_data_out_12),
	.feedback_valid_out(feedback_valid_out_12),
	.feedback_stall_in(feedback_stall_in_12)
);

defparam local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_feedback.STALLFREE = 0;
defparam local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_feedback.DATA_WIDTH = 32;
defparam local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_feedback.FIFO_DEPTH = 3;
defparam local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_feedback.STYLE = "REGULAR";

assign local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_inputs_ready = (local_bb2_notexitcond9__valid_out_0_NO_SHIFT_REG & rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_output_regs_ready = (&(~(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_valid_out_NO_SHIFT_REG) | ~(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_stall_in)));
assign local_bb2_notexitcond9__stall_in_0 = (local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_stall_out | ~(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_inputs_ready));
assign rnode_2to3_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_0_NO_SHIFT_REG = (local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_stall_out | ~(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_inputs_ready));
assign local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_causedstall = (local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_inputs_ready && (local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_stall_out && !(~(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_NO_SHIFT_REG <= 'x;
		local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_output_regs_ready)
		begin
			local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_NO_SHIFT_REG <= local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_result;
			local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_valid_out_NO_SHIFT_REG <= local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_stall_in))
			begin
				local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_3to7_bb2_notexitcond9__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_stall_in_0_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_stall_in_1_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__1_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_valid_out_2_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_stall_in_2_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__2_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_valid_out_3_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_stall_in_3_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__3_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_valid_out_4_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_stall_in_4_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__4_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_reg_7_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG;
 logic rnode_3to7_bb2_notexitcond9__0_stall_out_reg_7_NO_SHIFT_REG;
 reg rnode_3to7_bb2_notexitcond9__0_consumed_0_NO_SHIFT_REG;
 reg rnode_3to7_bb2_notexitcond9__0_consumed_1_NO_SHIFT_REG;
 reg rnode_3to7_bb2_notexitcond9__0_consumed_2_NO_SHIFT_REG;
 reg rnode_3to7_bb2_notexitcond9__0_consumed_3_NO_SHIFT_REG;
 reg rnode_3to7_bb2_notexitcond9__0_consumed_4_NO_SHIFT_REG;
wire [95:0] rci_rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5;

acl_data_fifo rnode_3to7_bb2_notexitcond9__0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to7_bb2_notexitcond9__0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_3to7_bb2_notexitcond9__0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb2_notexitcond9__NO_SHIFT_REG),
	.data_out(rnode_3to7_bb2_notexitcond9__0_reg_7_NO_SHIFT_REG)
);

defparam rnode_3to7_bb2_notexitcond9__0_reg_7_fifo.DEPTH = 5;
defparam rnode_3to7_bb2_notexitcond9__0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_3to7_bb2_notexitcond9__0_reg_7_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_3to7_bb2_notexitcond9__0_reg_7_fifo.IMPL = "ll_reg";

assign rnode_3to7_bb2_notexitcond9__0_reg_7_inputs_ready_NO_SHIFT_REG = local_bb2_notexitcond9__valid_out_1_NO_SHIFT_REG;
assign local_bb2_notexitcond9__stall_in_1 = rnode_3to7_bb2_notexitcond9__0_stall_out_reg_7_NO_SHIFT_REG;
assign rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG = ((rnode_3to7_bb2_notexitcond9__0_stall_in_0_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_0_NO_SHIFT_REG)) | (rnode_3to7_bb2_notexitcond9__0_stall_in_1_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_1_NO_SHIFT_REG)) | (rnode_3to7_bb2_notexitcond9__0_stall_in_2_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_2_NO_SHIFT_REG)) | (rnode_3to7_bb2_notexitcond9__0_stall_in_3_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_3_NO_SHIFT_REG)) | (rnode_3to7_bb2_notexitcond9__0_stall_in_4_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_4_NO_SHIFT_REG)));
assign rnode_3to7_bb2_notexitcond9__0_valid_out_0_NO_SHIFT_REG = (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_0_NO_SHIFT_REG));
assign rnode_3to7_bb2_notexitcond9__0_valid_out_1_NO_SHIFT_REG = (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_1_NO_SHIFT_REG));
assign rnode_3to7_bb2_notexitcond9__0_valid_out_2_NO_SHIFT_REG = (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_2_NO_SHIFT_REG));
assign rnode_3to7_bb2_notexitcond9__0_valid_out_3_NO_SHIFT_REG = (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_3_NO_SHIFT_REG));
assign rnode_3to7_bb2_notexitcond9__0_valid_out_4_NO_SHIFT_REG = (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & ~(rnode_3to7_bb2_notexitcond9__0_consumed_4_NO_SHIFT_REG));
assign rnode_3to7_bb2_notexitcond9__0_NO_SHIFT_REG = rnode_3to7_bb2_notexitcond9__0_reg_7_NO_SHIFT_REG;
assign rnode_3to7_bb2_notexitcond9__1_NO_SHIFT_REG = rnode_3to7_bb2_notexitcond9__0_reg_7_NO_SHIFT_REG;
assign rnode_3to7_bb2_notexitcond9__2_NO_SHIFT_REG = rnode_3to7_bb2_notexitcond9__0_reg_7_NO_SHIFT_REG;
assign rnode_3to7_bb2_notexitcond9__3_NO_SHIFT_REG = rnode_3to7_bb2_notexitcond9__0_reg_7_NO_SHIFT_REG;
assign rnode_3to7_bb2_notexitcond9__4_NO_SHIFT_REG = rnode_3to7_bb2_notexitcond9__0_reg_7_NO_SHIFT_REG;
assign rci_rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5[63:0] = rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_1_NO_SHIFT_REG;
assign rci_rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5[95:64] = (local_bb2_var_ & 32'hFFFFFFFE);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_3to7_bb2_notexitcond9__0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_3to7_bb2_notexitcond9__0_consumed_1_NO_SHIFT_REG <= 1'b0;
		rnode_3to7_bb2_notexitcond9__0_consumed_2_NO_SHIFT_REG <= 1'b0;
		rnode_3to7_bb2_notexitcond9__0_consumed_3_NO_SHIFT_REG <= 1'b0;
		rnode_3to7_bb2_notexitcond9__0_consumed_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_3to7_bb2_notexitcond9__0_consumed_0_NO_SHIFT_REG <= (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & (rnode_3to7_bb2_notexitcond9__0_consumed_0_NO_SHIFT_REG | ~(rnode_3to7_bb2_notexitcond9__0_stall_in_0_NO_SHIFT_REG)) & rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG);
		rnode_3to7_bb2_notexitcond9__0_consumed_1_NO_SHIFT_REG <= (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & (rnode_3to7_bb2_notexitcond9__0_consumed_1_NO_SHIFT_REG | ~(rnode_3to7_bb2_notexitcond9__0_stall_in_1_NO_SHIFT_REG)) & rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG);
		rnode_3to7_bb2_notexitcond9__0_consumed_2_NO_SHIFT_REG <= (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & (rnode_3to7_bb2_notexitcond9__0_consumed_2_NO_SHIFT_REG | ~(rnode_3to7_bb2_notexitcond9__0_stall_in_2_NO_SHIFT_REG)) & rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG);
		rnode_3to7_bb2_notexitcond9__0_consumed_3_NO_SHIFT_REG <= (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & (rnode_3to7_bb2_notexitcond9__0_consumed_3_NO_SHIFT_REG | ~(rnode_3to7_bb2_notexitcond9__0_stall_in_3_NO_SHIFT_REG)) & rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG);
		rnode_3to7_bb2_notexitcond9__0_consumed_4_NO_SHIFT_REG <= (rnode_3to7_bb2_notexitcond9__0_valid_out_0_reg_7_NO_SHIFT_REG & (rnode_3to7_bb2_notexitcond9__0_consumed_4_NO_SHIFT_REG | ~(rnode_3to7_bb2_notexitcond9__0_stall_in_4_NO_SHIFT_REG)) & rnode_3to7_bb2_notexitcond9__0_stall_in_0_reg_7_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 161
//  * capacity = 161
 logic rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_NO_SHIFT_REG;
 logic rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_NO_SHIFT_REG;
 logic [95:0] rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_NO_SHIFT_REG;
 logic rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic [95:0] rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_NO_SHIFT_REG;
 logic rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_5),
	.data_out(rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_NO_SHIFT_REG)
);

defparam rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_fifo.DEPTH = 162;
defparam rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_fifo.DATA_WIDTH = 96;
defparam rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_fifo.IMPL = "ram";

assign rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_inputs_ready_NO_SHIFT_REG = (rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_1_NO_SHIFT_REG & local_bb2_var__valid_out_1);
assign rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign rnode_1to5_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_1_NO_SHIFT_REG = rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_var__stall_in_1 = rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_NO_SHIFT_REG = rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_reg_166_NO_SHIFT_REG;
assign rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_NO_SHIFT_REG;
assign rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_NO_SHIFT_REG = rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_reg_166_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb2_add_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb2_add_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb2_add_0_NO_SHIFT_REG;
 logic rnode_5to6_bb2_add_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb2_add_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb2_add_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb2_add_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb2_add_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb2_add_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb2_add_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb2_add_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb2_add_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb2_add_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in((local_bb2_add & 32'hFFFFFFFE)),
	.data_out(rnode_5to6_bb2_add_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb2_add_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb2_add_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb2_add_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb2_add_0_reg_6_fifo.IMPL = "ll_reg";

assign rnode_5to6_bb2_add_0_reg_6_inputs_ready_NO_SHIFT_REG = local_bb2_add_valid_out;
assign local_bb2_add_stall_in = rnode_5to6_bb2_add_0_stall_out_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb2_add_0_NO_SHIFT_REG = rnode_5to6_bb2_add_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb2_add_0_stall_in_reg_6_NO_SHIFT_REG = rnode_5to6_bb2_add_0_stall_in_NO_SHIFT_REG;
assign rnode_5to6_bb2_add_0_valid_out_NO_SHIFT_REG = rnode_5to6_bb2_add_0_valid_out_reg_6_NO_SHIFT_REG;

// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_NO_SHIFT_REG;
 logic rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_NO_SHIFT_REG;
 logic rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_NO_SHIFT_REG),
	.data_out(rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_NO_SHIFT_REG)
);

defparam rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_fifo.DEPTH = 163;
defparam rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_fifo.DATA_WIDTH = 32;
defparam rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_fifo.IMPL = "ram";

assign rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_inputs_ready_NO_SHIFT_REG = local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_valid_out_NO_SHIFT_REG;
assign local_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_stall_in = rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_NO_SHIFT_REG = rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_reg_166_NO_SHIFT_REG;
assign rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_in_reg_166_NO_SHIFT_REG = rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_in_NO_SHIFT_REG;
assign rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_valid_out_NO_SHIFT_REG = rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_inputs_ready;
 reg local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_valid_out_NO_SHIFT_REG;
wire local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_stall_in;
wire local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_output_regs_ready;
wire local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_result;
wire local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_valid_out;
wire local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_stall_out;
 reg local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_NO_SHIFT_REG;
wire local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_causedstall;

acl_push local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_3to7_bb2_notexitcond9__0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_NO_SHIFT_REG),
	.stall_out(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_stall_out),
	.valid_in(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_inputs_ready),
	.valid_out(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_valid_out),
	.stall_in(~(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_output_regs_ready)),
	.data_out(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_result),
	.feedback_out(feedback_data_out_16),
	.feedback_valid_out(feedback_valid_out_16),
	.feedback_stall_in(feedback_stall_in_16)
);

defparam local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_feedback.STALLFREE = 0;
defparam local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_feedback.DATA_WIDTH = 1;
defparam local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_feedback.FIFO_DEPTH = 3;
defparam local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_feedback.STYLE = "REGULAR";

assign local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_inputs_ready = (local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_valid_out_1_NO_SHIFT_REG & rnode_3to7_bb2_notexitcond9__0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_output_regs_ready = (&(~(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_valid_out_NO_SHIFT_REG) | ~(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_stall_in)));
assign local_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_stall_in_1 = (local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_stall_out | ~(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_inputs_ready));
assign rnode_3to7_bb2_notexitcond9__0_stall_in_0_NO_SHIFT_REG = (local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_stall_out | ~(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_inputs_ready));
assign local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_causedstall = (local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_inputs_ready && (local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_stall_out && !(~(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_NO_SHIFT_REG <= 'x;
		local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_output_regs_ready)
		begin
			local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_NO_SHIFT_REG <= local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_result;
			local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_valid_out_NO_SHIFT_REG <= local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_stall_in))
			begin
				local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul3722_push13_mul3722_pop13_inputs_ready;
 reg local_bb2_mul3722_push13_mul3722_pop13_valid_out_NO_SHIFT_REG;
wire local_bb2_mul3722_push13_mul3722_pop13_stall_in;
wire local_bb2_mul3722_push13_mul3722_pop13_output_regs_ready;
wire [31:0] local_bb2_mul3722_push13_mul3722_pop13_result;
wire local_bb2_mul3722_push13_mul3722_pop13_fu_valid_out;
wire local_bb2_mul3722_push13_mul3722_pop13_fu_stall_out;
 reg [31:0] local_bb2_mul3722_push13_mul3722_pop13_NO_SHIFT_REG;
wire local_bb2_mul3722_push13_mul3722_pop13_causedstall;

acl_push local_bb2_mul3722_push13_mul3722_pop13_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_3to7_bb2_notexitcond9__1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb2_mul3722_pop13_mul3722_NO_SHIFT_REG),
	.stall_out(local_bb2_mul3722_push13_mul3722_pop13_fu_stall_out),
	.valid_in(local_bb2_mul3722_push13_mul3722_pop13_inputs_ready),
	.valid_out(local_bb2_mul3722_push13_mul3722_pop13_fu_valid_out),
	.stall_in(~(local_bb2_mul3722_push13_mul3722_pop13_output_regs_ready)),
	.data_out(local_bb2_mul3722_push13_mul3722_pop13_result),
	.feedback_out(feedback_data_out_13),
	.feedback_valid_out(feedback_valid_out_13),
	.feedback_stall_in(feedback_stall_in_13)
);

defparam local_bb2_mul3722_push13_mul3722_pop13_feedback.STALLFREE = 0;
defparam local_bb2_mul3722_push13_mul3722_pop13_feedback.DATA_WIDTH = 32;
defparam local_bb2_mul3722_push13_mul3722_pop13_feedback.FIFO_DEPTH = 3;
defparam local_bb2_mul3722_push13_mul3722_pop13_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb2_mul3722_push13_mul3722_pop13_feedback.STYLE = "REGULAR";

assign local_bb2_mul3722_push13_mul3722_pop13_inputs_ready = (local_bb2_mul3722_pop13_mul3722_valid_out_0_NO_SHIFT_REG & rnode_3to7_bb2_notexitcond9__0_valid_out_1_NO_SHIFT_REG);
assign local_bb2_mul3722_push13_mul3722_pop13_output_regs_ready = (&(~(local_bb2_mul3722_push13_mul3722_pop13_valid_out_NO_SHIFT_REG) | ~(local_bb2_mul3722_push13_mul3722_pop13_stall_in)));
assign local_bb2_mul3722_pop13_mul3722_stall_in_0 = (local_bb2_mul3722_push13_mul3722_pop13_fu_stall_out | ~(local_bb2_mul3722_push13_mul3722_pop13_inputs_ready));
assign rnode_3to7_bb2_notexitcond9__0_stall_in_1_NO_SHIFT_REG = (local_bb2_mul3722_push13_mul3722_pop13_fu_stall_out | ~(local_bb2_mul3722_push13_mul3722_pop13_inputs_ready));
assign local_bb2_mul3722_push13_mul3722_pop13_causedstall = (local_bb2_mul3722_push13_mul3722_pop13_inputs_ready && (local_bb2_mul3722_push13_mul3722_pop13_fu_stall_out && !(~(local_bb2_mul3722_push13_mul3722_pop13_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul3722_push13_mul3722_pop13_NO_SHIFT_REG <= 'x;
		local_bb2_mul3722_push13_mul3722_pop13_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul3722_push13_mul3722_pop13_output_regs_ready)
		begin
			local_bb2_mul3722_push13_mul3722_pop13_NO_SHIFT_REG <= local_bb2_mul3722_push13_mul3722_pop13_result;
			local_bb2_mul3722_push13_mul3722_pop13_valid_out_NO_SHIFT_REG <= local_bb2_mul3722_push13_mul3722_pop13_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_mul3722_push13_mul3722_pop13_stall_in))
			begin
				local_bb2_mul3722_push13_mul3722_pop13_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_notcmp1125_push14_notcmp1125_pop14_inputs_ready;
 reg local_bb2_notcmp1125_push14_notcmp1125_pop14_valid_out_NO_SHIFT_REG;
wire local_bb2_notcmp1125_push14_notcmp1125_pop14_stall_in;
wire local_bb2_notcmp1125_push14_notcmp1125_pop14_output_regs_ready;
wire local_bb2_notcmp1125_push14_notcmp1125_pop14_result;
wire local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_valid_out;
wire local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_stall_out;
 reg local_bb2_notcmp1125_push14_notcmp1125_pop14_NO_SHIFT_REG;
wire local_bb2_notcmp1125_push14_notcmp1125_pop14_causedstall;

acl_push local_bb2_notcmp1125_push14_notcmp1125_pop14_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_3to7_bb2_notexitcond9__2_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb2_notcmp1125_pop14_notcmp1125_NO_SHIFT_REG),
	.stall_out(local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_stall_out),
	.valid_in(local_bb2_notcmp1125_push14_notcmp1125_pop14_inputs_ready),
	.valid_out(local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_valid_out),
	.stall_in(~(local_bb2_notcmp1125_push14_notcmp1125_pop14_output_regs_ready)),
	.data_out(local_bb2_notcmp1125_push14_notcmp1125_pop14_result),
	.feedback_out(feedback_data_out_14),
	.feedback_valid_out(feedback_valid_out_14),
	.feedback_stall_in(feedback_stall_in_14)
);

defparam local_bb2_notcmp1125_push14_notcmp1125_pop14_feedback.STALLFREE = 0;
defparam local_bb2_notcmp1125_push14_notcmp1125_pop14_feedback.DATA_WIDTH = 1;
defparam local_bb2_notcmp1125_push14_notcmp1125_pop14_feedback.FIFO_DEPTH = 3;
defparam local_bb2_notcmp1125_push14_notcmp1125_pop14_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb2_notcmp1125_push14_notcmp1125_pop14_feedback.STYLE = "REGULAR";

assign local_bb2_notcmp1125_push14_notcmp1125_pop14_inputs_ready = (local_bb2_notcmp1125_pop14_notcmp1125_valid_out_0_NO_SHIFT_REG & rnode_3to7_bb2_notexitcond9__0_valid_out_2_NO_SHIFT_REG);
assign local_bb2_notcmp1125_push14_notcmp1125_pop14_output_regs_ready = (&(~(local_bb2_notcmp1125_push14_notcmp1125_pop14_valid_out_NO_SHIFT_REG) | ~(local_bb2_notcmp1125_push14_notcmp1125_pop14_stall_in)));
assign local_bb2_notcmp1125_pop14_notcmp1125_stall_in_0 = (local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_stall_out | ~(local_bb2_notcmp1125_push14_notcmp1125_pop14_inputs_ready));
assign rnode_3to7_bb2_notexitcond9__0_stall_in_2_NO_SHIFT_REG = (local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_stall_out | ~(local_bb2_notcmp1125_push14_notcmp1125_pop14_inputs_ready));
assign local_bb2_notcmp1125_push14_notcmp1125_pop14_causedstall = (local_bb2_notcmp1125_push14_notcmp1125_pop14_inputs_ready && (local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_stall_out && !(~(local_bb2_notcmp1125_push14_notcmp1125_pop14_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_notcmp1125_push14_notcmp1125_pop14_NO_SHIFT_REG <= 'x;
		local_bb2_notcmp1125_push14_notcmp1125_pop14_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_notcmp1125_push14_notcmp1125_pop14_output_regs_ready)
		begin
			local_bb2_notcmp1125_push14_notcmp1125_pop14_NO_SHIFT_REG <= local_bb2_notcmp1125_push14_notcmp1125_pop14_result;
			local_bb2_notcmp1125_push14_notcmp1125_pop14_valid_out_NO_SHIFT_REG <= local_bb2_notcmp1125_push14_notcmp1125_pop14_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_notcmp1125_push14_notcmp1125_pop14_stall_in))
			begin
				local_bb2_notcmp1125_push14_notcmp1125_pop14_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_notexitcond1428_push15_notexitcond1428_pop15_inputs_ready;
 reg local_bb2_notexitcond1428_push15_notexitcond1428_pop15_valid_out_NO_SHIFT_REG;
wire local_bb2_notexitcond1428_push15_notexitcond1428_pop15_stall_in;
wire local_bb2_notexitcond1428_push15_notexitcond1428_pop15_output_regs_ready;
wire local_bb2_notexitcond1428_push15_notexitcond1428_pop15_result;
wire local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_valid_out;
wire local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_stall_out;
 reg local_bb2_notexitcond1428_push15_notexitcond1428_pop15_NO_SHIFT_REG;
wire local_bb2_notexitcond1428_push15_notexitcond1428_pop15_causedstall;
wire [1:0] rci_rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_7;

acl_push local_bb2_notexitcond1428_push15_notexitcond1428_pop15_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_3to7_bb2_notexitcond9__3_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb2_notexitcond1428_pop15_notexitcond1428_NO_SHIFT_REG),
	.stall_out(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_stall_out),
	.valid_in(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_inputs_ready),
	.valid_out(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_valid_out),
	.stall_in(~(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_output_regs_ready)),
	.data_out(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_result),
	.feedback_out(feedback_data_out_15),
	.feedback_valid_out(feedback_valid_out_15),
	.feedback_stall_in(feedback_stall_in_15)
);

defparam local_bb2_notexitcond1428_push15_notexitcond1428_pop15_feedback.STALLFREE = 0;
defparam local_bb2_notexitcond1428_push15_notexitcond1428_pop15_feedback.DATA_WIDTH = 1;
defparam local_bb2_notexitcond1428_push15_notexitcond1428_pop15_feedback.FIFO_DEPTH = 3;
defparam local_bb2_notexitcond1428_push15_notexitcond1428_pop15_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb2_notexitcond1428_push15_notexitcond1428_pop15_feedback.STYLE = "REGULAR";

assign local_bb2_notexitcond1428_push15_notexitcond1428_pop15_inputs_ready = (local_bb2_notexitcond1428_pop15_notexitcond1428_valid_out_0_NO_SHIFT_REG & rnode_3to7_bb2_notexitcond9__0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_notexitcond1428_push15_notexitcond1428_pop15_output_regs_ready = (&(~(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_valid_out_NO_SHIFT_REG) | ~(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_stall_in)));
assign local_bb2_notexitcond1428_pop15_notexitcond1428_stall_in_0 = (local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_stall_out | ~(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_inputs_ready));
assign rnode_3to7_bb2_notexitcond9__0_stall_in_3_NO_SHIFT_REG = (local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_stall_out | ~(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_inputs_ready));
assign local_bb2_notexitcond1428_push15_notexitcond1428_pop15_causedstall = (local_bb2_notexitcond1428_push15_notexitcond1428_pop15_inputs_ready && (local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_stall_out && !(~(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_output_regs_ready))));
assign rci_rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_7[0] = rstag_7to7_bb2_memdep_phi1_or;
assign rci_rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_7[1] = rnode_3to7_bb2_notexitcond9__4_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_notexitcond1428_push15_notexitcond1428_pop15_NO_SHIFT_REG <= 'x;
		local_bb2_notexitcond1428_push15_notexitcond1428_pop15_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_notexitcond1428_push15_notexitcond1428_pop15_output_regs_ready)
		begin
			local_bb2_notexitcond1428_push15_notexitcond1428_pop15_NO_SHIFT_REG <= local_bb2_notexitcond1428_push15_notexitcond1428_pop15_result;
			local_bb2_notexitcond1428_push15_notexitcond1428_pop15_valid_out_NO_SHIFT_REG <= local_bb2_notexitcond1428_push15_notexitcond1428_pop15_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_notexitcond1428_push15_notexitcond1428_pop15_stall_in))
			begin
				local_bb2_notexitcond1428_push15_notexitcond1428_pop15_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 159
//  * capacity = 159
 logic rcnode_7to166_rc4_bb2_memdep_phi1_or_0_valid_out_NO_SHIFT_REG;
 logic rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_in_NO_SHIFT_REG;
 logic [1:0] rcnode_7to166_rc4_bb2_memdep_phi1_or_0_NO_SHIFT_REG;
 logic rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic [1:0] rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_NO_SHIFT_REG;
 logic rcnode_7to166_rc4_bb2_memdep_phi1_or_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_7to166_rc4_bb2_memdep_phi1_or_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_7),
	.data_out(rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_NO_SHIFT_REG)
);

defparam rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_fifo.DEPTH = 160;
defparam rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_fifo.DATA_WIDTH = 2;
defparam rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_fifo.IMPL = "ram";

assign rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_inputs_ready_NO_SHIFT_REG = (rnode_3to7_bb2_notexitcond9__0_valid_out_4_NO_SHIFT_REG & rstag_7to7_bb2_memdep_phi1_or_valid_out_0);
assign rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign rnode_3to7_bb2_notexitcond9__0_stall_in_4_NO_SHIFT_REG = rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rstag_7to7_bb2_memdep_phi1_or_stall_in_0 = rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_7to166_rc4_bb2_memdep_phi1_or_0_NO_SHIFT_REG = rcnode_7to166_rc4_bb2_memdep_phi1_or_0_reg_166_NO_SHIFT_REG;
assign rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_in_NO_SHIFT_REG;
assign rcnode_7to166_rc4_bb2_memdep_phi1_or_0_valid_out_NO_SHIFT_REG = rcnode_7to166_rc4_bb2_memdep_phi1_or_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_idxprom_stall_local;
wire [63:0] local_bb2_idxprom;
wire [34:0] rci_rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_8;

assign local_bb2_idxprom[63:32] = 32'h0;
assign local_bb2_idxprom[31:0] = (rnode_5to6_bb2_add_0_NO_SHIFT_REG & 32'hFFFFFFFE);
assign rci_rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_8[0] = local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_NO_SHIFT_REG;
assign rci_rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_8[32:1] = local_bb2_mul3722_push13_mul3722_pop13_NO_SHIFT_REG;
assign rci_rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_8[33] = local_bb2_notcmp1125_push14_notcmp1125_pop14_NO_SHIFT_REG;
assign rci_rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_8[34] = local_bb2_notexitcond1428_push15_notexitcond1428_pop15_NO_SHIFT_REG;

// Register node:
//  * latency = 158
//  * capacity = 158
 logic rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_valid_out_NO_SHIFT_REG;
 logic rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_in_NO_SHIFT_REG;
 logic [34:0] rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_NO_SHIFT_REG;
 logic rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic [34:0] rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_NO_SHIFT_REG;
 logic rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_8),
	.data_out(rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_NO_SHIFT_REG)
);

defparam rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_fifo.DEPTH = 159;
defparam rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_fifo.DATA_WIDTH = 35;
defparam rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_fifo.IMPL = "ram";

assign rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_inputs_ready_NO_SHIFT_REG = (local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_valid_out_NO_SHIFT_REG & local_bb2_mul3722_push13_mul3722_pop13_valid_out_NO_SHIFT_REG & local_bb2_notcmp1125_push14_notcmp1125_pop14_valid_out_NO_SHIFT_REG & local_bb2_notexitcond1428_push15_notexitcond1428_pop15_valid_out_NO_SHIFT_REG);
assign rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign local_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_stall_in = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_mul3722_push13_mul3722_pop13_stall_in = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_notcmp1125_push14_notcmp1125_pop14_stall_in = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign local_bb2_notexitcond1428_push15_notexitcond1428_pop15_stall_in = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_NO_SHIFT_REG = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_reg_166_NO_SHIFT_REG;
assign rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_in_NO_SHIFT_REG;
assign rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_valid_out_NO_SHIFT_REG = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx_valid_out;
wire local_bb2_arrayidx_stall_in;
wire local_bb2_arrayidx_inputs_ready;
wire local_bb2_arrayidx_stall_local;
wire [63:0] local_bb2_arrayidx;
wire [328:0] rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166;

assign local_bb2_arrayidx_inputs_ready = rnode_5to6_bb2_add_0_valid_out_NO_SHIFT_REG;
assign local_bb2_arrayidx = ((input_in & 64'hFFFFFFFFFFFFFC00) + ((local_bb2_idxprom & 64'hFFFFFFFE) << 6'h2));
assign local_bb2_arrayidx_valid_out = local_bb2_arrayidx_inputs_ready;
assign local_bb2_arrayidx_stall_local = local_bb2_arrayidx_stall_in;
assign rnode_5to6_bb2_add_0_stall_in_NO_SHIFT_REG = (|local_bb2_arrayidx_stall_local);
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[31:0] = (rcnode_2to166_rc1_bb2_mul5_0_NO_SHIFT_REG[31:0] & 32'hFFFFFFFE);
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[63:32] = rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_NO_SHIFT_REG[31:0];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[127:64] = rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_NO_SHIFT_REG[63:0];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[128] = rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_NO_SHIFT_REG[32];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[129] = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_NO_SHIFT_REG[0];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[161:130] = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_NO_SHIFT_REG[32:1];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[162] = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_NO_SHIFT_REG[33];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[163] = rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_NO_SHIFT_REG[34];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[195:164] = rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_NO_SHIFT_REG;
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[259:196] = rcnode_2to166_rc1_bb2_mul5_0_NO_SHIFT_REG[95:32];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[260] = rcnode_7to166_rc4_bb2_memdep_phi1_or_0_NO_SHIFT_REG[0];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[261] = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_NO_SHIFT_REG[0];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[293:262] = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_NO_SHIFT_REG[32:1];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[294] = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_NO_SHIFT_REG[33];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[295] = rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_NO_SHIFT_REG[34];
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[327:296] = (rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_NO_SHIFT_REG[95:64] & 32'hFFFFFFFE);
assign rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166[328] = rcnode_7to166_rc4_bb2_memdep_phi1_or_0_NO_SHIFT_REG[1];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_166to167_rc0_bb2_mul5_0_valid_out_NO_SHIFT_REG;
 logic rcnode_166to167_rc0_bb2_mul5_0_stall_in_NO_SHIFT_REG;
 logic [328:0] rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG;
 logic rcnode_166to167_rc0_bb2_mul5_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [328:0] rcnode_166to167_rc0_bb2_mul5_0_reg_167_NO_SHIFT_REG;
 logic rcnode_166to167_rc0_bb2_mul5_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rcnode_166to167_rc0_bb2_mul5_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_IP_NO_SHIFT_REG;
 logic rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;

acl_data_fifo rcnode_166to167_rc0_bb2_mul5_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_166to167_rc0_bb2_mul5_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_166to167_rc0_bb2_mul5_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rcnode_166to167_rc0_bb2_mul5_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_166to167_rc0_bb2_mul5_0_reg_166),
	.data_out(rcnode_166to167_rc0_bb2_mul5_0_reg_167_NO_SHIFT_REG)
);

defparam rcnode_166to167_rc0_bb2_mul5_0_reg_167_fifo.DEPTH = 1;
defparam rcnode_166to167_rc0_bb2_mul5_0_reg_167_fifo.DATA_WIDTH = 329;
defparam rcnode_166to167_rc0_bb2_mul5_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_166to167_rc0_bb2_mul5_0_reg_167_fifo.IMPL = "ll_reg";

assign rcnode_166to167_rc0_bb2_mul5_0_reg_167_inputs_ready_NO_SHIFT_REG = (rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_valid_out_NO_SHIFT_REG & rcnode_2to166_rc1_bb2_mul5_0_valid_out_NO_SHIFT_REG & rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_valid_out_NO_SHIFT_REG & rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_valid_out_NO_SHIFT_REG & rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_valid_out_NO_SHIFT_REG & rcnode_7to166_rc4_bb2_memdep_phi1_or_0_valid_out_NO_SHIFT_REG & rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_valid_out_NO_SHIFT_REG);
assign rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG = (~(rcnode_166to167_rc0_bb2_mul5_0_reg_167_inputs_ready_NO_SHIFT_REG) | rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_IP_NO_SHIFT_REG);
assign rnode_4to166_bb2_pixel_y_020_pop819_push12_pixel_y_020_pop819_pop12_0_stall_in_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;
assign rcnode_2to166_rc1_bb2_mul5_0_stall_in_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;
assign rcnode_3to166_rc1_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_0_stall_in_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;
assign rcnode_5to166_rc1_bb2_indvars_iv_pop10_acl_pop_i64_0_0_stall_in_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;
assign rcnode_7to166_rc2_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_0_stall_in_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;
assign rcnode_7to166_rc4_bb2_memdep_phi1_or_0_stall_in_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;
assign rcnode_8to166_rc0_bb2_memdep_phi1_pop931_push16_memdep_phi1_pop931_pop16_0_stall_in_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_out_0_reg_167_NO_SHIFT_REG;
assign rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_reg_167_NO_SHIFT_REG;
assign rcnode_166to167_rc0_bb2_mul5_0_stall_in_reg_167_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_stall_in_NO_SHIFT_REG;
assign rcnode_166to167_rc0_bb2_mul5_0_valid_out_NO_SHIFT_REG = rcnode_166to167_rc0_bb2_mul5_0_valid_out_reg_167_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb2_arrayidx_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb2_arrayidx_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_6to7_bb2_arrayidx_0_NO_SHIFT_REG;
 logic rnode_6to7_bb2_arrayidx_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_6to7_bb2_arrayidx_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb2_arrayidx_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb2_arrayidx_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb2_arrayidx_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb2_arrayidx_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb2_arrayidx_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb2_arrayidx_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb2_arrayidx_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb2_arrayidx_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in((local_bb2_arrayidx & 64'hFFFFFFFFFFFFFFF8)),
	.data_out(rnode_6to7_bb2_arrayidx_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb2_arrayidx_0_reg_7_fifo.DEPTH = 2;
defparam rnode_6to7_bb2_arrayidx_0_reg_7_fifo.DATA_WIDTH = 64;
defparam rnode_6to7_bb2_arrayidx_0_reg_7_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_6to7_bb2_arrayidx_0_reg_7_fifo.IMPL = "ll_reg";

assign rnode_6to7_bb2_arrayidx_0_reg_7_inputs_ready_NO_SHIFT_REG = local_bb2_arrayidx_valid_out;
assign local_bb2_arrayidx_stall_in = rnode_6to7_bb2_arrayidx_0_stall_out_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb2_arrayidx_0_NO_SHIFT_REG = rnode_6to7_bb2_arrayidx_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb2_arrayidx_0_stall_in_reg_7_NO_SHIFT_REG = rnode_6to7_bb2_arrayidx_0_stall_in_NO_SHIFT_REG;
assign rnode_6to7_bb2_arrayidx_0_valid_out_NO_SHIFT_REG = rnode_6to7_bb2_arrayidx_0_valid_out_reg_7_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb2_ld__inputs_ready;
 reg local_bb2_ld__valid_out_NO_SHIFT_REG;
wire local_bb2_ld__stall_in;
wire local_bb2_ld__output_regs_ready;
wire local_bb2_ld__fu_stall_out;
wire local_bb2_ld__fu_valid_out;
wire [31:0] local_bb2_ld__lsu_dataout;
 reg [31:0] local_bb2_ld__NO_SHIFT_REG;
wire local_bb2_ld__causedstall;

lsu_top lsu_local_bb2_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld__fu_stall_out),
	.i_valid(local_bb2_ld__inputs_ready),
	.i_address((rnode_6to7_bb2_arrayidx_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFF8)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(input_wii_var_),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld__output_regs_ready)),
	.o_valid(local_bb2_ld__fu_valid_out),
	.o_readdata(local_bb2_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld__active),
	.avm_address(avm_local_bb2_ld__address),
	.avm_read(avm_local_bb2_ld__read),
	.avm_readdata(avm_local_bb2_ld__readdata),
	.avm_write(avm_local_bb2_ld__write),
	.avm_writeack(avm_local_bb2_ld__writeack),
	.avm_burstcount(avm_local_bb2_ld__burstcount),
	.avm_writedata(avm_local_bb2_ld__writedata),
	.avm_byteenable(avm_local_bb2_ld__byteenable),
	.avm_waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld_.AWIDTH = 33;
defparam lsu_local_bb2_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb2_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb2_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb2_ld_.ALIGNMENT_BYTES = 8;
defparam lsu_local_bb2_ld_.READ = 1;
defparam lsu_local_bb2_ld_.ATOMIC = 0;
defparam lsu_local_bb2_ld_.WIDTH = 32;
defparam lsu_local_bb2_ld_.MWIDTH = 512;
defparam lsu_local_bb2_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld_.MEMORY_SIDE_MEM_LATENCY = 99;
defparam lsu_local_bb2_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb2_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld_.USECACHING = 0;
defparam lsu_local_bb2_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld_.ADDRSPACE = 1;
defparam lsu_local_bb2_ld_.STYLE = "BURST-COALESCED";

assign local_bb2_ld__inputs_ready = (rnode_6to7_bb2_arrayidx_0_valid_out_NO_SHIFT_REG & rnode_1to7_var__0_valid_out_NO_SHIFT_REG & rstag_7to7_bb2_memdep_phi1_or_valid_out_1);
assign local_bb2_ld__output_regs_ready = (&(~(local_bb2_ld__valid_out_NO_SHIFT_REG) | ~(local_bb2_ld__stall_in)));
assign rnode_6to7_bb2_arrayidx_0_stall_in_NO_SHIFT_REG = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign rnode_1to7_var__0_stall_in_NO_SHIFT_REG = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign rstag_7to7_bb2_memdep_phi1_or_stall_in_1 = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign local_bb2_ld__causedstall = (local_bb2_ld__inputs_ready && (local_bb2_ld__fu_stall_out && !(~(local_bb2_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld__NO_SHIFT_REG <= 'x;
		local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld__output_regs_ready)
		begin
			local_bb2_ld__NO_SHIFT_REG <= local_bb2_ld__lsu_dataout;
			local_bb2_ld__valid_out_NO_SHIFT_REG <= local_bb2_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld__stall_in))
			begin
				local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_167to167_bb2_ld__valid_out;
wire rstag_167to167_bb2_ld__stall_in;
wire rstag_167to167_bb2_ld__inputs_ready;
wire rstag_167to167_bb2_ld__stall_local;
 reg rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG;
wire rstag_167to167_bb2_ld__combined_valid;
 reg [31:0] rstag_167to167_bb2_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_167to167_bb2_ld_;

assign rstag_167to167_bb2_ld__inputs_ready = local_bb2_ld__valid_out_NO_SHIFT_REG;
assign rstag_167to167_bb2_ld_ = (rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG ? rstag_167to167_bb2_ld__staging_reg_NO_SHIFT_REG : local_bb2_ld__NO_SHIFT_REG);
assign rstag_167to167_bb2_ld__combined_valid = (rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG | rstag_167to167_bb2_ld__inputs_ready);
assign rstag_167to167_bb2_ld__valid_out = rstag_167to167_bb2_ld__combined_valid;
assign rstag_167to167_bb2_ld__stall_local = rstag_167to167_bb2_ld__stall_in;
assign local_bb2_ld__stall_in = (|rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_167to167_bb2_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_167to167_bb2_ld__stall_local)
		begin
			if (~(rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG <= rstag_167to167_bb2_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_167to167_bb2_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_167to167_bb2_ld__staging_reg_NO_SHIFT_REG <= local_bb2_ld__NO_SHIFT_REG;
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [31:0] lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb2_mul5_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb2_indvars_iv_pop10_acl_pop_i64_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb2_var__reg_NO_SHIFT_REG;
 reg lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_reg_NO_SHIFT_REG;
 reg lvb_bb2_memdep_phi1_or_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb2_ld__reg_NO_SHIFT_REG;
 reg lvb_bb2_notcmp_reg_NO_SHIFT_REG;
 reg lvb_bb2_notexitcond9__reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb2_mul3722_pop13_mul3722_reg_NO_SHIFT_REG;
 reg lvb_bb2_notcmp1125_pop14_notcmp1125_reg_NO_SHIFT_REG;
 reg lvb_bb2_notexitcond1428_pop15_notexitcond1428_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb2_notcmp_valid_out & rcnode_166to167_rc0_bb2_mul5_0_valid_out_NO_SHIFT_REG & rstag_167to167_bb2_ld__valid_out);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb2_notcmp_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_166to167_rc0_bb2_mul5_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_167to167_bb2_ld__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819 = lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_reg_NO_SHIFT_REG;
assign lvb_bb2_mul5 = lvb_bb2_mul5_reg_NO_SHIFT_REG;
assign lvb_bb2_indvars_iv_pop10_acl_pop_i64_0 = lvb_bb2_indvars_iv_pop10_acl_pop_i64_0_reg_NO_SHIFT_REG;
assign lvb_bb2_var_ = lvb_bb2_var__reg_NO_SHIFT_REG;
assign lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931 = lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_reg_NO_SHIFT_REG;
assign lvb_bb2_memdep_phi1_or = lvb_bb2_memdep_phi1_or_reg_NO_SHIFT_REG;
assign lvb_bb2_ld_ = lvb_bb2_ld__reg_NO_SHIFT_REG;
assign lvb_bb2_notcmp = lvb_bb2_notcmp_reg_NO_SHIFT_REG;
assign lvb_bb2_notexitcond9_ = lvb_bb2_notexitcond9__reg_NO_SHIFT_REG;
assign lvb_bb2_mul3722_pop13_mul3722 = lvb_bb2_mul3722_pop13_mul3722_reg_NO_SHIFT_REG;
assign lvb_bb2_notcmp1125_pop14_notcmp1125 = lvb_bb2_notcmp1125_pop14_notcmp1125_reg_NO_SHIFT_REG;
assign lvb_bb2_notexitcond1428_pop15_notexitcond1428 = lvb_bb2_notexitcond1428_pop15_notexitcond1428_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_mul5_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_indvars_iv_pop10_acl_pop_i64_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_var__reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_memdep_phi1_or_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_ld__reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_notcmp_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_notexitcond9__reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_mul3722_pop13_mul3722_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_notcmp1125_pop14_notcmp1125_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_notexitcond1428_pop15_notexitcond1428_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819_reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[63:32];
			lvb_bb2_mul5_reg_NO_SHIFT_REG <= (rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[31:0] & 32'hFFFFFFFE);
			lvb_bb2_indvars_iv_pop10_acl_pop_i64_0_reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[127:64];
			lvb_bb2_var__reg_NO_SHIFT_REG <= (rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[327:296] & 32'hFFFFFFFE);
			lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931_reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[129];
			lvb_bb2_memdep_phi1_or_reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[260];
			lvb_bb2_ld__reg_NO_SHIFT_REG <= rstag_167to167_bb2_ld_;
			lvb_bb2_notcmp_reg_NO_SHIFT_REG <= local_bb2_notcmp;
			lvb_bb2_notexitcond9__reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[328];
			lvb_bb2_mul3722_pop13_mul3722_reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[161:130];
			lvb_bb2_notcmp1125_pop14_notcmp1125_reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[162];
			lvb_bb2_notexitcond1428_pop15_notexitcond1428_reg_NO_SHIFT_REG <= rcnode_166to167_rc0_bb2_mul5_0_NO_SHIFT_REG[163];
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_3
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_inSize_x,
		input [31:0] 		input_r,
		input [31:0] 		input_wii_div,
		input [31:0] 		input_wii_div1,
		input 		input_wii_cmp19,
		input [31:0] 		input_wii_add7,
		input [31:0] 		input_wii_sub20,
		input [31:0] 		input_wii_sub22,
		input 		input_wii_var_,
		input 		input_wii_var__u12,
		input 		input_wii_var__u13,
		input 		input_wii_var__u14,
		input 		valid_in_0,
		output 		stall_out_0,
		input 		input_forked16_0,
		input [31:0] 		input_pixel_y_020_pop820_0,
		input [31:0] 		input_mul3723_0,
		input 		input_notcmp1126_0,
		input 		input_notexitcond1429_0,
		input 		input_memdep_phi1_pop932_0,
		input [31:0] 		input_mul534_0,
		input [63:0] 		input_indvars_iv_pop1036_0,
		input [31:0] 		input_var__u15_0,
		input 		input_memdep_phi1_or38_0,
		input [31:0] 		input_var__u16_0,
		input 		input_notcmp40_0,
		input 		input_notexitcond942_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input 		input_forked16_1,
		input [31:0] 		input_pixel_y_020_pop820_1,
		input [31:0] 		input_mul3723_1,
		input 		input_notcmp1126_1,
		input 		input_notexitcond1429_1,
		input 		input_memdep_phi1_pop932_1,
		input [31:0] 		input_mul534_1,
		input [63:0] 		input_indvars_iv_pop1036_1,
		input [31:0] 		input_var__u15_1,
		input 		input_memdep_phi1_or38_1,
		input [31:0] 		input_var__u16_1,
		input 		input_notcmp40_1,
		input 		input_notexitcond942_1,
		output 		valid_out,
		input 		stall_in,
		output 		lvb_forked16,
		output [31:0] 		lvb_bb3_c0_exe1,
		output [31:0] 		lvb_bb3_c0_exe2,
		output 		lvb_bb3_c0_exe3,
		output 		lvb_bb3_c0_exe4,
		output [31:0] 		lvb_bb3_c0_exe5,
		output [31:0] 		lvb_bb3_c0_exe6,
		output 		lvb_bb3_c0_exe7,
		output 		lvb_bb3_c0_exe8,
		output 		lvb_bb3_c0_exe9,
		output [63:0] 		lvb_bb3_c0_exe10,
		output [31:0] 		lvb_bb3_c0_exe11,
		output 		lvb_bb3_c0_exe12,
		output [31:0] 		lvb_bb3_c0_exe13,
		output 		lvb_bb3_c0_exe14,
		output 		lvb_bb3_c0_exe15,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		feedback_valid_in_17,
		output 		feedback_stall_out_17,
		input [31:0] 		feedback_data_in_17,
		input 		feedback_valid_in_23,
		output 		feedback_stall_out_23,
		input [31:0] 		feedback_data_in_23,
		output 		feedback_stall_out_2,
		input 		feedback_valid_in_3,
		output 		feedback_stall_out_3,
		input 		feedback_data_in_3,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		input 		feedback_valid_in_18,
		output 		feedback_stall_out_18,
		input [31:0] 		feedback_data_in_18,
		input 		feedback_valid_in_19,
		output 		feedback_stall_out_19,
		input [31:0] 		feedback_data_in_19,
		input 		feedback_valid_in_20,
		output 		feedback_stall_out_20,
		input 		feedback_data_in_20,
		input 		feedback_valid_in_21,
		output 		feedback_stall_out_21,
		input 		feedback_data_in_21,
		input 		feedback_valid_in_22,
		output 		feedback_stall_out_22,
		input 		feedback_data_in_22,
		input 		feedback_valid_in_24,
		output 		feedback_stall_out_24,
		input [63:0] 		feedback_data_in_24,
		input 		feedback_valid_in_25,
		output 		feedback_stall_out_25,
		input [31:0] 		feedback_data_in_25,
		input 		feedback_valid_in_26,
		output 		feedback_stall_out_26,
		input 		feedback_data_in_26,
		input 		feedback_valid_in_27,
		output 		feedback_stall_out_27,
		input [31:0] 		feedback_data_in_27,
		input 		feedback_valid_in_28,
		output 		feedback_stall_out_28,
		input 		feedback_data_in_28,
		input 		feedback_valid_in_29,
		output 		feedback_stall_out_29,
		input 		feedback_data_in_29,
		output 		feedback_valid_out_3,
		input 		feedback_stall_in_3,
		output 		feedback_data_out_3,
		output 		feedback_valid_out_17,
		input 		feedback_stall_in_17,
		output [31:0] 		feedback_data_out_17,
		output 		feedback_valid_out_23,
		input 		feedback_stall_in_23,
		output [31:0] 		feedback_data_out_23,
		output 		feedback_valid_out_18,
		input 		feedback_stall_in_18,
		output [31:0] 		feedback_data_out_18,
		output 		feedback_valid_out_19,
		input 		feedback_stall_in_19,
		output [31:0] 		feedback_data_out_19,
		output 		feedback_valid_out_20,
		input 		feedback_stall_in_20,
		output 		feedback_data_out_20,
		output 		feedback_valid_out_21,
		input 		feedback_stall_in_21,
		output 		feedback_data_out_21,
		output 		feedback_valid_out_22,
		input 		feedback_stall_in_22,
		output 		feedback_data_out_22,
		output 		feedback_valid_out_24,
		input 		feedback_stall_in_24,
		output [63:0] 		feedback_data_out_24,
		output 		feedback_valid_out_25,
		input 		feedback_stall_in_25,
		output [31:0] 		feedback_data_out_25,
		output 		feedback_valid_out_26,
		input 		feedback_stall_in_26,
		output 		feedback_data_out_26,
		output 		feedback_valid_out_27,
		input 		feedback_stall_in_27,
		output [31:0] 		feedback_data_out_27,
		output 		feedback_valid_out_28,
		input 		feedback_stall_in_28,
		output 		feedback_data_out_28,
		output 		feedback_valid_out_29,
		input 		feedback_stall_in_29,
		output 		feedback_data_out_29
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_node_stall_in_8;
 reg merge_node_valid_out_8_NO_SHIFT_REG;
wire merge_node_stall_in_9;
 reg merge_node_valid_out_9_NO_SHIFT_REG;
wire merge_node_stall_in_10;
 reg merge_node_valid_out_10_NO_SHIFT_REG;
wire merge_node_stall_in_11;
 reg merge_node_valid_out_11_NO_SHIFT_REG;
wire merge_node_stall_in_12;
 reg merge_node_valid_out_12_NO_SHIFT_REG;
wire merge_node_stall_in_13;
 reg merge_node_valid_out_13_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg input_forked16_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pixel_y_020_pop820_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul3723_0_staging_reg_NO_SHIFT_REG;
 reg input_notcmp1126_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1429_0_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_pop932_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul534_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_pop1036_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u15_0_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_or38_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u16_0_staging_reg_NO_SHIFT_REG;
 reg input_notcmp40_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond942_0_staging_reg_NO_SHIFT_REG;
 reg local_lvm_forked16_NO_SHIFT_REG;
 reg [31:0] local_lvm_pixel_y_020_pop820_NO_SHIFT_REG;
 reg [31:0] local_lvm_mul3723_NO_SHIFT_REG;
 reg local_lvm_notcmp1126_NO_SHIFT_REG;
 reg local_lvm_notexitcond1429_NO_SHIFT_REG;
 reg local_lvm_memdep_phi1_pop932_NO_SHIFT_REG;
 reg [31:0] local_lvm_mul534_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv_pop1036_NO_SHIFT_REG;
 reg [31:0] local_lvm_var__u15_NO_SHIFT_REG;
 reg local_lvm_memdep_phi1_or38_NO_SHIFT_REG;
 reg [31:0] local_lvm_var__u16_NO_SHIFT_REG;
 reg local_lvm_notcmp40_NO_SHIFT_REG;
 reg local_lvm_notexitcond942_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg input_forked16_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pixel_y_020_pop820_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul3723_1_staging_reg_NO_SHIFT_REG;
 reg input_notcmp1126_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1429_1_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_pop932_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul534_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_pop1036_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u15_1_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_or38_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u16_1_staging_reg_NO_SHIFT_REG;
 reg input_notcmp40_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond942_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG) | (merge_node_stall_in_8 & merge_node_valid_out_8_NO_SHIFT_REG) | (merge_node_stall_in_9 & merge_node_valid_out_9_NO_SHIFT_REG) | (merge_node_stall_in_10 & merge_node_valid_out_10_NO_SHIFT_REG) | (merge_node_stall_in_11 & merge_node_valid_out_11_NO_SHIFT_REG) | (merge_node_stall_in_12 & merge_node_valid_out_12_NO_SHIFT_REG) | (merge_node_stall_in_13 & merge_node_valid_out_13_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_forked16_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_pixel_y_020_pop820_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul3723_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp1126_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1429_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_pop932_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul534_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_pop1036_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u15_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_or38_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u16_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp40_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond942_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_forked16_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_pixel_y_020_pop820_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul3723_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp1126_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1429_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_pop932_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul534_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_pop1036_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u15_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_or38_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u16_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp40_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond942_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_forked16_0_staging_reg_NO_SHIFT_REG <= input_forked16_0;
				input_pixel_y_020_pop820_0_staging_reg_NO_SHIFT_REG <= input_pixel_y_020_pop820_0;
				input_mul3723_0_staging_reg_NO_SHIFT_REG <= input_mul3723_0;
				input_notcmp1126_0_staging_reg_NO_SHIFT_REG <= input_notcmp1126_0;
				input_notexitcond1429_0_staging_reg_NO_SHIFT_REG <= input_notexitcond1429_0;
				input_memdep_phi1_pop932_0_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_pop932_0;
				input_mul534_0_staging_reg_NO_SHIFT_REG <= input_mul534_0;
				input_indvars_iv_pop1036_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv_pop1036_0;
				input_var__u15_0_staging_reg_NO_SHIFT_REG <= input_var__u15_0;
				input_memdep_phi1_or38_0_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_or38_0;
				input_var__u16_0_staging_reg_NO_SHIFT_REG <= input_var__u16_0;
				input_notcmp40_0_staging_reg_NO_SHIFT_REG <= input_notcmp40_0;
				input_notexitcond942_0_staging_reg_NO_SHIFT_REG <= input_notexitcond942_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_forked16_1_staging_reg_NO_SHIFT_REG <= input_forked16_1;
				input_pixel_y_020_pop820_1_staging_reg_NO_SHIFT_REG <= input_pixel_y_020_pop820_1;
				input_mul3723_1_staging_reg_NO_SHIFT_REG <= input_mul3723_1;
				input_notcmp1126_1_staging_reg_NO_SHIFT_REG <= input_notcmp1126_1;
				input_notexitcond1429_1_staging_reg_NO_SHIFT_REG <= input_notexitcond1429_1;
				input_memdep_phi1_pop932_1_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_pop932_1;
				input_mul534_1_staging_reg_NO_SHIFT_REG <= input_mul534_1;
				input_indvars_iv_pop1036_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv_pop1036_1;
				input_var__u15_1_staging_reg_NO_SHIFT_REG <= input_var__u15_1;
				input_memdep_phi1_or38_1_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_or38_1;
				input_var__u16_1_staging_reg_NO_SHIFT_REG <= input_var__u16_1;
				input_notcmp40_1_staging_reg_NO_SHIFT_REG <= input_notcmp40_1;
				input_notexitcond942_1_staging_reg_NO_SHIFT_REG <= input_notexitcond942_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked16_NO_SHIFT_REG <= input_forked16_0_staging_reg_NO_SHIFT_REG;
					local_lvm_pixel_y_020_pop820_NO_SHIFT_REG <= input_pixel_y_020_pop820_0_staging_reg_NO_SHIFT_REG;
					local_lvm_mul3723_NO_SHIFT_REG <= input_mul3723_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp1126_NO_SHIFT_REG <= input_notcmp1126_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1429_NO_SHIFT_REG <= input_notexitcond1429_0_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_pop932_NO_SHIFT_REG <= input_memdep_phi1_pop932_0_staging_reg_NO_SHIFT_REG;
					local_lvm_mul534_NO_SHIFT_REG <= input_mul534_0_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_pop1036_NO_SHIFT_REG <= input_indvars_iv_pop1036_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u15_NO_SHIFT_REG <= input_var__u15_0_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_or38_NO_SHIFT_REG <= input_memdep_phi1_or38_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp40_NO_SHIFT_REG <= input_notcmp40_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond942_NO_SHIFT_REG <= input_notexitcond942_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked16_NO_SHIFT_REG <= input_forked16_0;
					local_lvm_pixel_y_020_pop820_NO_SHIFT_REG <= input_pixel_y_020_pop820_0;
					local_lvm_mul3723_NO_SHIFT_REG <= input_mul3723_0;
					local_lvm_notcmp1126_NO_SHIFT_REG <= input_notcmp1126_0;
					local_lvm_notexitcond1429_NO_SHIFT_REG <= input_notexitcond1429_0;
					local_lvm_memdep_phi1_pop932_NO_SHIFT_REG <= input_memdep_phi1_pop932_0;
					local_lvm_mul534_NO_SHIFT_REG <= input_mul534_0;
					local_lvm_indvars_iv_pop1036_NO_SHIFT_REG <= input_indvars_iv_pop1036_0;
					local_lvm_var__u15_NO_SHIFT_REG <= input_var__u15_0;
					local_lvm_memdep_phi1_or38_NO_SHIFT_REG <= input_memdep_phi1_or38_0;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_0;
					local_lvm_notcmp40_NO_SHIFT_REG <= input_notcmp40_0;
					local_lvm_notexitcond942_NO_SHIFT_REG <= input_notexitcond942_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked16_NO_SHIFT_REG <= input_forked16_1_staging_reg_NO_SHIFT_REG;
					local_lvm_pixel_y_020_pop820_NO_SHIFT_REG <= input_pixel_y_020_pop820_1_staging_reg_NO_SHIFT_REG;
					local_lvm_mul3723_NO_SHIFT_REG <= input_mul3723_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp1126_NO_SHIFT_REG <= input_notcmp1126_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1429_NO_SHIFT_REG <= input_notexitcond1429_1_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_pop932_NO_SHIFT_REG <= input_memdep_phi1_pop932_1_staging_reg_NO_SHIFT_REG;
					local_lvm_mul534_NO_SHIFT_REG <= input_mul534_1_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_pop1036_NO_SHIFT_REG <= input_indvars_iv_pop1036_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u15_NO_SHIFT_REG <= input_var__u15_1_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_or38_NO_SHIFT_REG <= input_memdep_phi1_or38_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp40_NO_SHIFT_REG <= input_notcmp40_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond942_NO_SHIFT_REG <= input_notexitcond942_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked16_NO_SHIFT_REG <= input_forked16_1;
					local_lvm_pixel_y_020_pop820_NO_SHIFT_REG <= input_pixel_y_020_pop820_1;
					local_lvm_mul3723_NO_SHIFT_REG <= input_mul3723_1;
					local_lvm_notcmp1126_NO_SHIFT_REG <= input_notcmp1126_1;
					local_lvm_notexitcond1429_NO_SHIFT_REG <= input_notexitcond1429_1;
					local_lvm_memdep_phi1_pop932_NO_SHIFT_REG <= input_memdep_phi1_pop932_1;
					local_lvm_mul534_NO_SHIFT_REG <= input_mul534_1;
					local_lvm_indvars_iv_pop1036_NO_SHIFT_REG <= input_indvars_iv_pop1036_1;
					local_lvm_var__u15_NO_SHIFT_REG <= input_var__u15_1;
					local_lvm_memdep_phi1_or38_NO_SHIFT_REG <= input_memdep_phi1_or38_1;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_1;
					local_lvm_notcmp40_NO_SHIFT_REG <= input_notcmp40_1;
					local_lvm_notexitcond942_NO_SHIFT_REG <= input_notexitcond942_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_9_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_10_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_11_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_12_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_13_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_8_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_9_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_10_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_11_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_12_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_13_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_8))
			begin
				merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_9))
			begin
				merge_node_valid_out_9_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_10))
			begin
				merge_node_valid_out_10_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_11))
			begin
				merge_node_valid_out_11_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_12))
			begin
				merge_node_valid_out_12_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_13))
			begin
				merge_node_valid_out_13_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni1_stall_local;
wire [383:0] local_bb3_c0_eni1;

assign local_bb3_c0_eni1[7:0] = 8'bx;
assign local_bb3_c0_eni1[8] = local_lvm_forked16_NO_SHIFT_REG;
assign local_bb3_c0_eni1[383:9] = 375'bx;

// Register node:
//  * latency = 9
//  * capacity = 9
 logic rnode_1to10_forked16_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to10_forked16_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to10_forked16_0_NO_SHIFT_REG;
 logic rnode_1to10_forked16_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to10_forked16_0_reg_10_NO_SHIFT_REG;
 logic rnode_1to10_forked16_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_1to10_forked16_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_1to10_forked16_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_1to10_forked16_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to10_forked16_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to10_forked16_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_1to10_forked16_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_1to10_forked16_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(local_lvm_forked16_NO_SHIFT_REG),
	.data_out(rnode_1to10_forked16_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_1to10_forked16_0_reg_10_fifo.DEPTH = 10;
defparam rnode_1to10_forked16_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_1to10_forked16_0_reg_10_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to10_forked16_0_reg_10_fifo.IMPL = "ram";

assign rnode_1to10_forked16_0_reg_10_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_13_NO_SHIFT_REG;
assign merge_node_stall_in_13 = rnode_1to10_forked16_0_stall_out_reg_10_NO_SHIFT_REG;
assign rnode_1to10_forked16_0_NO_SHIFT_REG = rnode_1to10_forked16_0_reg_10_NO_SHIFT_REG;
assign rnode_1to10_forked16_0_stall_in_reg_10_NO_SHIFT_REG = rnode_1to10_forked16_0_stall_in_NO_SHIFT_REG;
assign rnode_1to10_forked16_0_valid_out_NO_SHIFT_REG = rnode_1to10_forked16_0_valid_out_reg_10_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni2_stall_local;
wire [383:0] local_bb3_c0_eni2;

assign local_bb3_c0_eni2[31:0] = local_bb3_c0_eni1[31:0];
assign local_bb3_c0_eni2[63:32] = local_lvm_mul534_NO_SHIFT_REG;
assign local_bb3_c0_eni2[383:64] = local_bb3_c0_eni1[383:64];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_forked16_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_forked16_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_forked16_0_NO_SHIFT_REG;
 logic rnode_10to11_forked16_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_forked16_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_forked16_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_forked16_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_forked16_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_forked16_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_forked16_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_forked16_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_forked16_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_forked16_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(rnode_1to10_forked16_0_NO_SHIFT_REG),
	.data_out(rnode_10to11_forked16_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_forked16_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_forked16_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_forked16_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_forked16_0_reg_11_fifo.IMPL = "ll_reg";

assign rnode_10to11_forked16_0_reg_11_inputs_ready_NO_SHIFT_REG = rnode_1to10_forked16_0_valid_out_NO_SHIFT_REG;
assign rnode_1to10_forked16_0_stall_in_NO_SHIFT_REG = rnode_10to11_forked16_0_stall_out_reg_11_NO_SHIFT_REG;
assign rnode_10to11_forked16_0_NO_SHIFT_REG = rnode_10to11_forked16_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_forked16_0_stall_in_reg_11_NO_SHIFT_REG = rnode_10to11_forked16_0_stall_in_NO_SHIFT_REG;
assign rnode_10to11_forked16_0_valid_out_NO_SHIFT_REG = rnode_10to11_forked16_0_valid_out_reg_11_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni3_stall_local;
wire [383:0] local_bb3_c0_eni3;

assign local_bb3_c0_eni3[63:0] = local_bb3_c0_eni2[63:0];
assign local_bb3_c0_eni3[95:64] = local_lvm_pixel_y_020_pop820_NO_SHIFT_REG;
assign local_bb3_c0_eni3[383:96] = local_bb3_c0_eni2[383:96];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni4_stall_local;
wire [383:0] local_bb3_c0_eni4;

assign local_bb3_c0_eni4[95:0] = local_bb3_c0_eni3[95:0];
assign local_bb3_c0_eni4[127:96] = local_lvm_mul3723_NO_SHIFT_REG;
assign local_bb3_c0_eni4[383:128] = local_bb3_c0_eni3[383:128];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni5_stall_local;
wire [383:0] local_bb3_c0_eni5;

assign local_bb3_c0_eni5[127:0] = local_bb3_c0_eni4[127:0];
assign local_bb3_c0_eni5[128] = local_lvm_notcmp1126_NO_SHIFT_REG;
assign local_bb3_c0_eni5[383:129] = local_bb3_c0_eni4[383:129];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni6_stall_local;
wire [383:0] local_bb3_c0_eni6;

assign local_bb3_c0_eni6[135:0] = local_bb3_c0_eni5[135:0];
assign local_bb3_c0_eni6[136] = local_lvm_notexitcond1429_NO_SHIFT_REG;
assign local_bb3_c0_eni6[383:137] = local_bb3_c0_eni5[383:137];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni7_stall_local;
wire [383:0] local_bb3_c0_eni7;

assign local_bb3_c0_eni7[143:0] = local_bb3_c0_eni6[143:0];
assign local_bb3_c0_eni7[144] = local_lvm_memdep_phi1_pop932_NO_SHIFT_REG;
assign local_bb3_c0_eni7[383:145] = local_bb3_c0_eni6[383:145];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni8_stall_local;
wire [383:0] local_bb3_c0_eni8;

assign local_bb3_c0_eni8[191:0] = local_bb3_c0_eni7[191:0];
assign local_bb3_c0_eni8[255:192] = local_lvm_indvars_iv_pop1036_NO_SHIFT_REG;
assign local_bb3_c0_eni8[383:256] = local_bb3_c0_eni7[383:256];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni9_stall_local;
wire [383:0] local_bb3_c0_eni9;

assign local_bb3_c0_eni9[255:0] = local_bb3_c0_eni8[255:0];
assign local_bb3_c0_eni9[287:256] = local_lvm_var__u15_NO_SHIFT_REG;
assign local_bb3_c0_eni9[383:288] = local_bb3_c0_eni8[383:288];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni10_stall_local;
wire [383:0] local_bb3_c0_eni10;

assign local_bb3_c0_eni10[287:0] = local_bb3_c0_eni9[287:0];
assign local_bb3_c0_eni10[288] = local_lvm_memdep_phi1_or38_NO_SHIFT_REG;
assign local_bb3_c0_eni10[383:289] = local_bb3_c0_eni9[383:289];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni11_stall_local;
wire [383:0] local_bb3_c0_eni11;

assign local_bb3_c0_eni11[319:0] = local_bb3_c0_eni10[319:0];
assign local_bb3_c0_eni11[351:320] = local_lvm_var__u16_NO_SHIFT_REG;
assign local_bb3_c0_eni11[383:352] = local_bb3_c0_eni10[383:352];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni12_stall_local;
wire [383:0] local_bb3_c0_eni12;

assign local_bb3_c0_eni12[351:0] = local_bb3_c0_eni11[351:0];
assign local_bb3_c0_eni12[352] = local_lvm_notcmp40_NO_SHIFT_REG;
assign local_bb3_c0_eni12[383:353] = local_bb3_c0_eni11[383:353];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni13_stall_local;
wire [383:0] local_bb3_c0_eni13;

assign local_bb3_c0_eni13[359:0] = local_bb3_c0_eni12[359:0];
assign local_bb3_c0_eni13[360] = local_lvm_notexitcond942_NO_SHIFT_REG;
assign local_bb3_c0_eni13[383:361] = local_bb3_c0_eni12[383:361];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_valid_out_2;
wire local_bb3_c0_ene1_stall_in_2;
wire local_bb3_c0_ene3_valid_out;
wire local_bb3_c0_ene3_stall_in;
wire local_bb3_c0_ene4_valid_out;
wire local_bb3_c0_ene4_stall_in;
wire local_bb3_c0_ene5_valid_out;
wire local_bb3_c0_ene5_stall_in;
wire local_bb3_c0_ene6_valid_out;
wire local_bb3_c0_ene6_stall_in;
wire local_bb3_c0_ene7_valid_out;
wire local_bb3_c0_ene7_stall_in;
wire local_bb3_c0_ene8_valid_out;
wire local_bb3_c0_ene8_stall_in;
wire local_bb3_c0_ene9_valid_out;
wire local_bb3_c0_ene9_stall_in;
wire local_bb3_c0_ene10_valid_out;
wire local_bb3_c0_ene10_stall_in;
wire local_bb3_c0_ene11_valid_out;
wire local_bb3_c0_ene11_stall_in;
wire local_bb3_c0_ene12_valid_out;
wire local_bb3_c0_ene12_stall_in;
wire local_bb3_c0_ene13_valid_out;
wire local_bb3_c0_ene13_stall_in;
wire SFC_1_VALID_1_1_0_valid_out_0;
wire SFC_1_VALID_1_1_0_stall_in_0;
wire local_bb3_i_211_pop17_add7_valid_out_1;
wire local_bb3_i_211_pop17_add7_stall_in_1;
wire local_bb3_mul534_pop23_c0_ene2_valid_out_1;
wire local_bb3_mul534_pop23_c0_ene2_stall_in_1;
wire local_bb3_add17_valid_out;
wire local_bb3_add17_stall_in;
wire local_bb3_c0_enter_c0_eni13_inputs_ready;
wire local_bb3_c0_enter_c0_eni13_stall_local;
wire local_bb3_c0_enter_c0_eni13_input_accepted;
wire [383:0] local_bb3_c0_enter_c0_eni13;
wire local_bb3_c0_exit_c0_exi15_entry_stall;
wire local_bb3_c0_enter_c0_eni13_valid_bit;
wire local_bb3_c0_exit_c0_exi15_output_regs_ready;
wire local_bb3_c0_exit_c0_exi15_valid_in;
wire local_bb3_c0_exit_c0_exi15_phases;
wire local_bb3_c0_enter_c0_eni13_inc_pipelined_thread;
wire local_bb3_c0_enter_c0_eni13_dec_pipelined_thread;
wire local_bb3_c0_enter_c0_eni13_fu_stall_out;

assign local_bb3_c0_enter_c0_eni13_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_3_NO_SHIFT_REG & merge_node_valid_out_4_NO_SHIFT_REG & merge_node_valid_out_5_NO_SHIFT_REG & merge_node_valid_out_6_NO_SHIFT_REG & merge_node_valid_out_7_NO_SHIFT_REG & merge_node_valid_out_8_NO_SHIFT_REG & merge_node_valid_out_9_NO_SHIFT_REG & merge_node_valid_out_10_NO_SHIFT_REG & merge_node_valid_out_11_NO_SHIFT_REG & merge_node_valid_out_12_NO_SHIFT_REG);
assign local_bb3_c0_enter_c0_eni13 = local_bb3_c0_eni13;
assign local_bb3_c0_enter_c0_eni13_input_accepted = (local_bb3_c0_enter_c0_eni13_inputs_ready && !(local_bb3_c0_exit_c0_exi15_entry_stall));
assign local_bb3_c0_enter_c0_eni13_valid_bit = local_bb3_c0_enter_c0_eni13_input_accepted;
assign local_bb3_c0_enter_c0_eni13_inc_pipelined_thread = 1'b1;
assign local_bb3_c0_enter_c0_eni13_dec_pipelined_thread = ~(1'b0);
assign local_bb3_c0_enter_c0_eni13_fu_stall_out = (~(local_bb3_c0_enter_c0_eni13_inputs_ready) | local_bb3_c0_exit_c0_exi15_entry_stall);
assign local_bb3_c0_enter_c0_eni13_stall_local = (local_bb3_c0_ene1_stall_in_2 | local_bb3_c0_ene3_stall_in | local_bb3_c0_ene4_stall_in | local_bb3_c0_ene5_stall_in | local_bb3_c0_ene6_stall_in | local_bb3_c0_ene7_stall_in | local_bb3_c0_ene8_stall_in | local_bb3_c0_ene9_stall_in | local_bb3_c0_ene10_stall_in | local_bb3_c0_ene11_stall_in | local_bb3_c0_ene12_stall_in | local_bb3_c0_ene13_stall_in | SFC_1_VALID_1_1_0_stall_in_0 | local_bb3_i_211_pop17_add7_stall_in_1 | local_bb3_mul534_pop23_c0_ene2_stall_in_1 | local_bb3_add17_stall_in);
assign local_bb3_c0_ene1_valid_out_2 = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene3_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene4_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene5_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene6_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene7_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene8_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene9_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene10_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene11_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene12_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_c0_ene13_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign SFC_1_VALID_1_1_0_valid_out_0 = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_i_211_pop17_add7_valid_out_1 = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_mul534_pop23_c0_ene2_valid_out_1 = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign local_bb3_add17_valid_out = local_bb3_c0_enter_c0_eni13_inputs_ready;
assign merge_node_stall_in_0 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_1 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_2 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_3 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_4 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_5 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_6 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_7 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_8 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_9 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_10 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_11 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));
assign merge_node_stall_in_12 = (local_bb3_c0_enter_c0_eni13_fu_stall_out | ~(local_bb3_c0_enter_c0_eni13_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_stall_local;
wire local_bb3_c0_ene1;

assign local_bb3_c0_ene1 = local_bb3_c0_enter_c0_eni13[8];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene2_stall_local;
wire [31:0] local_bb3_c0_ene2;

assign local_bb3_c0_ene2 = local_bb3_c0_enter_c0_eni13[63:32];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene3_stall_local;
wire [31:0] local_bb3_c0_ene3;

assign local_bb3_c0_ene3 = local_bb3_c0_enter_c0_eni13[95:64];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene4_stall_local;
wire [31:0] local_bb3_c0_ene4;

assign local_bb3_c0_ene4 = local_bb3_c0_enter_c0_eni13[127:96];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene5_stall_local;
wire local_bb3_c0_ene5;

assign local_bb3_c0_ene5 = local_bb3_c0_enter_c0_eni13[128];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene6_stall_local;
wire local_bb3_c0_ene6;

assign local_bb3_c0_ene6 = local_bb3_c0_enter_c0_eni13[136];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene7_stall_local;
wire local_bb3_c0_ene7;

assign local_bb3_c0_ene7 = local_bb3_c0_enter_c0_eni13[144];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene8_stall_local;
wire [63:0] local_bb3_c0_ene8;

assign local_bb3_c0_ene8 = local_bb3_c0_enter_c0_eni13[255:192];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene9_stall_local;
wire [31:0] local_bb3_c0_ene9;

assign local_bb3_c0_ene9 = local_bb3_c0_enter_c0_eni13[287:256];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene10_stall_local;
wire local_bb3_c0_ene10;

assign local_bb3_c0_ene10 = local_bb3_c0_enter_c0_eni13[288];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene11_stall_local;
wire [31:0] local_bb3_c0_ene11;

assign local_bb3_c0_ene11 = local_bb3_c0_enter_c0_eni13[351:320];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene12_stall_local;
wire local_bb3_c0_ene12;

assign local_bb3_c0_ene12 = local_bb3_c0_enter_c0_eni13[352];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene13_stall_local;
wire local_bb3_c0_ene13;

assign local_bb3_c0_ene13 = local_bb3_c0_enter_c0_eni13[360];

// This section implements an unregistered operation.
// 
wire SFC_1_VALID_1_1_0_stall_local;
wire SFC_1_VALID_1_1_0;

assign SFC_1_VALID_1_1_0 = local_bb3_c0_enter_c0_eni13_valid_bit;

// This section implements an unregistered operation.
// 
wire local_bb3_i_211_pop17_add7_stall_local;
wire [31:0] local_bb3_i_211_pop17_add7;
wire local_bb3_i_211_pop17_add7_fu_valid_out;
wire local_bb3_i_211_pop17_add7_fu_stall_out;

acl_pop local_bb3_i_211_pop17_add7_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_c0_ene1),
	.predicate(1'b0),
	.data_in(input_wii_add7),
	.stall_out(local_bb3_i_211_pop17_add7_fu_stall_out),
	.valid_in(SFC_1_VALID_1_1_0),
	.valid_out(local_bb3_i_211_pop17_add7_fu_valid_out),
	.stall_in(local_bb3_i_211_pop17_add7_stall_local),
	.data_out(local_bb3_i_211_pop17_add7),
	.feedback_in(feedback_data_in_17),
	.feedback_valid_in(feedback_valid_in_17),
	.feedback_stall_out(feedback_stall_out_17)
);

defparam local_bb3_i_211_pop17_add7_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_i_211_pop17_add7_feedback.DATA_WIDTH = 32;
defparam local_bb3_i_211_pop17_add7_feedback.STYLE = "REGULAR";

assign local_bb3_i_211_pop17_add7_stall_local = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_mul534_pop23_c0_ene2_stall_local;
wire [31:0] local_bb3_mul534_pop23_c0_ene2;
wire local_bb3_mul534_pop23_c0_ene2_fu_valid_out;
wire local_bb3_mul534_pop23_c0_ene2_fu_stall_out;

acl_pop local_bb3_mul534_pop23_c0_ene2_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_c0_ene1),
	.predicate(1'b0),
	.data_in(local_bb3_c0_ene2),
	.stall_out(local_bb3_mul534_pop23_c0_ene2_fu_stall_out),
	.valid_in(SFC_1_VALID_1_1_0),
	.valid_out(local_bb3_mul534_pop23_c0_ene2_fu_valid_out),
	.stall_in(local_bb3_mul534_pop23_c0_ene2_stall_local),
	.data_out(local_bb3_mul534_pop23_c0_ene2),
	.feedback_in(feedback_data_in_23),
	.feedback_valid_in(feedback_valid_in_23),
	.feedback_stall_out(feedback_stall_out_23)
);

defparam local_bb3_mul534_pop23_c0_ene2_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_mul534_pop23_c0_ene2_feedback.DATA_WIDTH = 32;
defparam local_bb3_mul534_pop23_c0_ene2_feedback.STYLE = "REGULAR";

assign local_bb3_mul534_pop23_c0_ene2_stall_local = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_add17_stall_local;
wire [31:0] local_bb3_add17;

assign local_bb3_add17 = (local_bb3_i_211_pop17_add7 + local_bb3_mul534_pop23_c0_ene2);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_c0_ene1_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_c0_ene1_0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_c0_ene1_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene1),
	.data_out(rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene1_stall_in_2 = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_1_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene3_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene3_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene3_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene3_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene3_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene3_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene3_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene3_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene3_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene3_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene3),
	.data_out(rnode_1to3_bb3_c0_ene3_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene3_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene3_0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_1to3_bb3_c0_ene3_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene3_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene3_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene3_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene3_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene3_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene3_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene4_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene4_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene4_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene4_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene4_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene4_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene4_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene4_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene4_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene4_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene4),
	.data_out(rnode_1to3_bb3_c0_ene4_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene4_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene4_0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_1to3_bb3_c0_ene4_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene4_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene4_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene4_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene4_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene4_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene4_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene5_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene5_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene5_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene5_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene5_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene5_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene5_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene5_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene5_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene5_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene5),
	.data_out(rnode_1to3_bb3_c0_ene5_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene5_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene5_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb3_c0_ene5_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene5_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene5_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene5_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene5_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene5_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene5_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene6_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene6_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene6_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene6_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene6_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene6_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene6_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene6_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene6_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene6_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene6),
	.data_out(rnode_1to3_bb3_c0_ene6_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene6_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene6_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb3_c0_ene6_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene6_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene6_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene6_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene6_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene6_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene6_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene7_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene7_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene7_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene7_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene7_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene7_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene7_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene7_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene7_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene7_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene7),
	.data_out(rnode_1to3_bb3_c0_ene7_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene7_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene7_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb3_c0_ene7_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene7_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene7_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene7_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene7_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene7_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene7_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene8_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_1to3_bb3_c0_ene8_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene8_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to3_bb3_c0_ene8_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene8_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene8_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene8_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene8_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene8_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene8_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene8_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene8_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene8),
	.data_out(rnode_1to3_bb3_c0_ene8_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene8_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene8_0_reg_3_fifo.DATA_WIDTH = 64;
defparam rnode_1to3_bb3_c0_ene8_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene8_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene8_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene8_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene8_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene8_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene8_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene9_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene9_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene9_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene9_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene9_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene9_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene9_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene9_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene9_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene9_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene9_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene9_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene9_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene9),
	.data_out(rnode_1to3_bb3_c0_ene9_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene9_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene9_0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_1to3_bb3_c0_ene9_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene9_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene9_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene9_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene9_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene9_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene9_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene9_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene10_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene10_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene10_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene10_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene10_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene10_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene10_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene10_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene10_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene10_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene10_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene10_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene10_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene10),
	.data_out(rnode_1to3_bb3_c0_ene10_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene10_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene10_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb3_c0_ene10_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene10_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene10_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene10_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene10_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene10_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene10_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene10_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene11_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene11_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene11_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene11_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_c0_ene11_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene11_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene11_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene11_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene11_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene11_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene11_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene11_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene11_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene11),
	.data_out(rnode_1to3_bb3_c0_ene11_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene11_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene11_0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_1to3_bb3_c0_ene11_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene11_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene11_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene11_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene11_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene11_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene11_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene11_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene12_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene12_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene12_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene12_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene12_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene12_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene12_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene12_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene12_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene12_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene12_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene12_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene12_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene12),
	.data_out(rnode_1to3_bb3_c0_ene12_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene12_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene12_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb3_c0_ene12_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene12_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene12_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene12_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene12_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene12_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene12_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene12_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_c0_ene13_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene13_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene13_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene13_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene13_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene13_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene13_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_c0_ene13_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_c0_ene13_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_c0_ene13_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_c0_ene13_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_c0_ene13_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_c0_ene13_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene13),
	.data_out(rnode_1to3_bb3_c0_ene13_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_c0_ene13_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_c0_ene13_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb3_c0_ene13_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_c0_ene13_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_c0_ene13_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene13_stall_in = 1'b0;
assign rnode_1to3_bb3_c0_ene13_0_NO_SHIFT_REG = rnode_1to3_bb3_c0_ene13_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_c0_ene13_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_c0_ene13_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_1_2_0_inputs_ready;
 reg SFC_1_VALID_1_2_0_valid_out_0_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_0;
 reg SFC_1_VALID_1_2_0_valid_out_1_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_1;
 reg SFC_1_VALID_1_2_0_valid_out_2_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_2;
 reg SFC_1_VALID_1_2_0_valid_out_3_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_3;
wire SFC_1_VALID_1_2_0_output_regs_ready;
 reg SFC_1_VALID_1_2_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_1_2_0_causedstall;

assign SFC_1_VALID_1_2_0_inputs_ready = 1'b1;
assign SFC_1_VALID_1_2_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_1_1_0_stall_in_0 = 1'b0;
assign SFC_1_VALID_1_2_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_1_2_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_1_2_0_output_regs_ready)
		begin
			SFC_1_VALID_1_2_0_NO_SHIFT_REG <= SFC_1_VALID_1_1_0;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_i_211_pop17_add7_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb3_i_211_pop17_add7_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_i_211_pop17_add7_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_i_211_pop17_add7_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_i_211_pop17_add7_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_i_211_pop17_add7_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_i_211_pop17_add7_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_i_211_pop17_add7_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_i_211_pop17_add7_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_i_211_pop17_add7),
	.data_out(rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_i_211_pop17_add7_stall_in_1 = 1'b0;
assign rnode_1to2_bb3_i_211_pop17_add7_0_NO_SHIFT_REG = rnode_1to2_bb3_i_211_pop17_add7_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_i_211_pop17_add7_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_i_211_pop17_add7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_mul534_pop23_c0_ene2_1_NO_SHIFT_REG;
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_valid_out_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_in_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_in_0_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb3_mul534_pop23_c0_ene2_0_valid_out_0_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_mul534_pop23_c0_ene2),
	.data_out(rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_mul534_pop23_c0_ene2_stall_in_1 = 1'b0;
assign rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_in_0_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb3_mul534_pop23_c0_ene2_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to3_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG = rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb3_mul534_pop23_c0_ene2_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to3_bb3_mul534_pop23_c0_ene2_1_NO_SHIFT_REG = rnode_1to3_bb3_mul534_pop23_c0_ene2_0_reg_3_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_add17_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_add17_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_add17_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_add17_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb3_add17_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_add17_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_add17_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_add17_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_add17_0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_add17_0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_add17_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_add17),
	.data_out(rnode_1to2_bb3_add17_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_add17_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_add17_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb3_add17_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_add17_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb3_add17_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add17_stall_in = 1'b0;
assign rnode_1to2_bb3_add17_0_stall_in_0_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_add17_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_add17_0_NO_SHIFT_REG = rnode_1to2_bb3_add17_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_add17_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_add17_1_NO_SHIFT_REG = rnode_1to2_bb3_add17_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_add17_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_add17_2_NO_SHIFT_REG = rnode_1to2_bb3_add17_0_reg_2_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_1_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_2_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_4_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_4_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_5_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_5_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_5_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_6_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_6_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_6_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_7_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_7_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_7_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_8_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_8_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_8_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_9_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_9_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_9_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_10_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_10_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_10_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_c0_ene1_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_c0_ene1_0_stall_in_0_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_c0_ene1_0_valid_out_0_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_c0_ene1_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb3_c0_ene1_1_NO_SHIFT_REG),
	.data_out(rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_0_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_1_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_2_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_3_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_4_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_5_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_5_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_6_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_6_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_7_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_7_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_8_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_8_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_9_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_9_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_10_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_c0_ene1_10_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_1_VALID_2_3_0_inputs_ready;
 reg SFC_1_VALID_2_3_0_valid_out_0_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_0;
 reg SFC_1_VALID_2_3_0_valid_out_1_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_1;
 reg SFC_1_VALID_2_3_0_valid_out_2_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_2;
 reg SFC_1_VALID_2_3_0_valid_out_3_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_3;
 reg SFC_1_VALID_2_3_0_valid_out_4_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_4;
 reg SFC_1_VALID_2_3_0_valid_out_5_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_5;
 reg SFC_1_VALID_2_3_0_valid_out_6_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_6;
 reg SFC_1_VALID_2_3_0_valid_out_7_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_7;
 reg SFC_1_VALID_2_3_0_valid_out_8_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_8;
 reg SFC_1_VALID_2_3_0_valid_out_9_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_9;
 reg SFC_1_VALID_2_3_0_valid_out_10_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_10;
 reg SFC_1_VALID_2_3_0_valid_out_11_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_11;
 reg SFC_1_VALID_2_3_0_valid_out_12_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_12;
 reg SFC_1_VALID_2_3_0_valid_out_13_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_13;
 reg SFC_1_VALID_2_3_0_valid_out_14_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_14;
 reg SFC_1_VALID_2_3_0_valid_out_15_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_15;
 reg SFC_1_VALID_2_3_0_valid_out_16_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_16;
 reg SFC_1_VALID_2_3_0_valid_out_17_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_17;
 reg SFC_1_VALID_2_3_0_valid_out_18_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_18;
 reg SFC_1_VALID_2_3_0_valid_out_19_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_19;
 reg SFC_1_VALID_2_3_0_valid_out_20_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_20;
 reg SFC_1_VALID_2_3_0_valid_out_21_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_21;
 reg SFC_1_VALID_2_3_0_valid_out_22_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_22;
 reg SFC_1_VALID_2_3_0_valid_out_23_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in_23;
wire SFC_1_VALID_2_3_0_output_regs_ready;
 reg SFC_1_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_2_3_0_causedstall;

assign SFC_1_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_1_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_1_2_0_stall_in_0 = 1'b0;
assign SFC_1_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_2_3_0_output_regs_ready)
		begin
			SFC_1_VALID_2_3_0_NO_SHIFT_REG <= SFC_1_VALID_1_2_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_keep_going4_acl_pipeline_1_inputs_ready;
 reg local_bb3_keep_going4_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb3_keep_going4_acl_pipeline_1_stall_in;
wire local_bb3_keep_going4_acl_pipeline_1_output_regs_ready;
wire local_bb3_keep_going4_acl_pipeline_1_keep_going;
wire local_bb3_keep_going4_acl_pipeline_1_fu_valid_out;
wire local_bb3_keep_going4_acl_pipeline_1_fu_stall_out;
 reg local_bb3_keep_going4_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb3_keep_going4_acl_pipeline_1_feedback_pipelined;
wire local_bb3_keep_going4_acl_pipeline_1_causedstall;

acl_pipeline local_bb3_keep_going4_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb3_keep_going4_acl_pipeline_1_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_keep_going4_acl_pipeline_1_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_keep_going4_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_2),
	.not_exitcond_in(feedback_data_in_3),
	.not_exitcond_valid_in(feedback_valid_in_3),
	.not_exitcond_stall_out(feedback_stall_out_3),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb3_keep_going4_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb3_keep_going4_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb3_keep_going4_acl_pipeline_1_inputs_ready = 1'b1;
assign local_bb3_keep_going4_acl_pipeline_1_output_regs_ready = 1'b1;
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign SFC_1_VALID_1_2_0_stall_in_1 = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb3_keep_going4_acl_pipeline_1_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_keep_going4_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb3_keep_going4_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_keep_going4_acl_pipeline_1_output_regs_ready)
		begin
			local_bb3_keep_going4_acl_pipeline_1_NO_SHIFT_REG <= local_bb3_keep_going4_acl_pipeline_1_keep_going;
			local_bb3_keep_going4_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_keep_going4_acl_pipeline_1_stall_in))
			begin
				local_bb3_keep_going4_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_inc34_stall_local;
wire [31:0] local_bb3_inc34;

assign local_bb3_inc34 = (rnode_1to2_bb3_i_211_pop17_add7_0_NO_SHIFT_REG + 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_mul534_pop23_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul534_pop23_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul534_pop23_c0_ene2_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_mul534_pop23_c0_ene2_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(rnode_1to3_bb3_mul534_pop23_c0_ene2_1_NO_SHIFT_REG),
	.data_out(rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG = rnode_3to4_bb3_mul534_pop23_c0_ene2_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_mul534_pop23_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i1_i_valid_out;
wire local_bb3_cmp_i1_i_stall_in;
wire local_bb3_cmp_i1_i_inputs_ready;
wire local_bb3_cmp_i1_i_stall_local;
wire local_bb3_cmp_i1_i;

assign local_bb3_cmp_i1_i_inputs_ready = rnode_1to2_bb3_add17_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_cmp_i1_i = ($signed(rnode_1to2_bb3_add17_0_NO_SHIFT_REG) < $signed(32'h0));
assign local_bb3_cmp_i1_i_valid_out = 1'b1;
assign rnode_1to2_bb3_add17_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp1_i3_i_valid_out;
wire local_bb3_cmp1_i3_i_stall_in;
wire local_bb3_cmp1_i3_i_inputs_ready;
wire local_bb3_cmp1_i3_i_stall_local;
wire local_bb3_cmp1_i3_i;

assign local_bb3_cmp1_i3_i_inputs_ready = rnode_1to2_bb3_add17_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_cmp1_i3_i = ($signed(rnode_1to2_bb3_add17_1_NO_SHIFT_REG) > $signed(input_wii_sub22));
assign local_bb3_cmp1_i3_i_valid_out = 1'b1;
assign rnode_1to2_bb3_add17_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_add17_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_add17_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to3_bb3_add17_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_add17_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to3_bb3_add17_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_add17_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_add17_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_add17_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_add17_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_add17_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_add17_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_add17_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_add17_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb3_add17_2_NO_SHIFT_REG),
	.data_out(rnode_2to3_bb3_add17_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_add17_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_add17_0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_2to3_bb3_add17_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_add17_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_add17_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_add17_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_add17_0_NO_SHIFT_REG = rnode_2to3_bb3_add17_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_add17_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_add17_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_3_4_0_inputs_ready;
 reg SFC_1_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_3_4_0_stall_in;
wire SFC_1_VALID_3_4_0_output_regs_ready;
 reg SFC_1_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_3_4_0_causedstall;

assign SFC_1_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_1_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_0 = 1'b0;
assign SFC_1_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_3_4_0_output_regs_ready)
		begin
			SFC_1_VALID_3_4_0_NO_SHIFT_REG <= SFC_1_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_valid_out_0;
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_stall_in_0;
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_valid_out_1;
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_stall_in_1;
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_inputs_ready;
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_stall_local;
wire [31:0] local_bb3_pixel_y_020_pop820_pop18_c0_ene3;
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_fu_valid_out;
wire local_bb3_pixel_y_020_pop820_pop18_c0_ene3_fu_stall_out;

acl_pop local_bb3_pixel_y_020_pop820_pop18_c0_ene3_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene3_0_NO_SHIFT_REG),
	.stall_out(local_bb3_pixel_y_020_pop820_pop18_c0_ene3_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_pixel_y_020_pop820_pop18_c0_ene3_fu_valid_out),
	.stall_in(local_bb3_pixel_y_020_pop820_pop18_c0_ene3_stall_local),
	.data_out(local_bb3_pixel_y_020_pop820_pop18_c0_ene3),
	.feedback_in(feedback_data_in_18),
	.feedback_valid_in(feedback_valid_in_18),
	.feedback_stall_out(feedback_stall_out_18)
);

defparam local_bb3_pixel_y_020_pop820_pop18_c0_ene3_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_pixel_y_020_pop820_pop18_c0_ene3_feedback.DATA_WIDTH = 32;
defparam local_bb3_pixel_y_020_pop820_pop18_c0_ene3_feedback.STYLE = "REGULAR";

assign local_bb3_pixel_y_020_pop820_pop18_c0_ene3_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_1_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene3_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG);
assign local_bb3_pixel_y_020_pop820_pop18_c0_ene3_stall_local = 1'b0;
assign local_bb3_pixel_y_020_pop820_pop18_c0_ene3_valid_out_0 = 1'b1;
assign local_bb3_pixel_y_020_pop820_pop18_c0_ene3_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_1 = 1'b0;
assign rnode_1to3_bb3_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_mul3723_pop19_c0_ene4_valid_out_0;
wire local_bb3_mul3723_pop19_c0_ene4_stall_in_0;
wire local_bb3_mul3723_pop19_c0_ene4_valid_out_1;
wire local_bb3_mul3723_pop19_c0_ene4_stall_in_1;
wire local_bb3_mul3723_pop19_c0_ene4_inputs_ready;
wire local_bb3_mul3723_pop19_c0_ene4_stall_local;
wire [31:0] local_bb3_mul3723_pop19_c0_ene4;
wire local_bb3_mul3723_pop19_c0_ene4_fu_valid_out;
wire local_bb3_mul3723_pop19_c0_ene4_fu_stall_out;

acl_pop local_bb3_mul3723_pop19_c0_ene4_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene4_0_NO_SHIFT_REG),
	.stall_out(local_bb3_mul3723_pop19_c0_ene4_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_mul3723_pop19_c0_ene4_fu_valid_out),
	.stall_in(local_bb3_mul3723_pop19_c0_ene4_stall_local),
	.data_out(local_bb3_mul3723_pop19_c0_ene4),
	.feedback_in(feedback_data_in_19),
	.feedback_valid_in(feedback_valid_in_19),
	.feedback_stall_out(feedback_stall_out_19)
);

defparam local_bb3_mul3723_pop19_c0_ene4_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_mul3723_pop19_c0_ene4_feedback.DATA_WIDTH = 32;
defparam local_bb3_mul3723_pop19_c0_ene4_feedback.STYLE = "REGULAR";

assign local_bb3_mul3723_pop19_c0_ene4_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_2_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene4_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG);
assign local_bb3_mul3723_pop19_c0_ene4_stall_local = 1'b0;
assign local_bb3_mul3723_pop19_c0_ene4_valid_out_0 = 1'b1;
assign local_bb3_mul3723_pop19_c0_ene4_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_2 = 1'b0;
assign rnode_1to3_bb3_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_notcmp1126_pop20_c0_ene5_valid_out_0;
wire local_bb3_notcmp1126_pop20_c0_ene5_stall_in_0;
wire local_bb3_notcmp1126_pop20_c0_ene5_valid_out_1;
wire local_bb3_notcmp1126_pop20_c0_ene5_stall_in_1;
wire local_bb3_notcmp1126_pop20_c0_ene5_inputs_ready;
wire local_bb3_notcmp1126_pop20_c0_ene5_stall_local;
wire local_bb3_notcmp1126_pop20_c0_ene5;
wire local_bb3_notcmp1126_pop20_c0_ene5_fu_valid_out;
wire local_bb3_notcmp1126_pop20_c0_ene5_fu_stall_out;

acl_pop local_bb3_notcmp1126_pop20_c0_ene5_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_2_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene5_0_NO_SHIFT_REG),
	.stall_out(local_bb3_notcmp1126_pop20_c0_ene5_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notcmp1126_pop20_c0_ene5_fu_valid_out),
	.stall_in(local_bb3_notcmp1126_pop20_c0_ene5_stall_local),
	.data_out(local_bb3_notcmp1126_pop20_c0_ene5),
	.feedback_in(feedback_data_in_20),
	.feedback_valid_in(feedback_valid_in_20),
	.feedback_stall_out(feedback_stall_out_20)
);

defparam local_bb3_notcmp1126_pop20_c0_ene5_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_notcmp1126_pop20_c0_ene5_feedback.DATA_WIDTH = 1;
defparam local_bb3_notcmp1126_pop20_c0_ene5_feedback.STYLE = "REGULAR";

assign local_bb3_notcmp1126_pop20_c0_ene5_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_3_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene5_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_2_NO_SHIFT_REG);
assign local_bb3_notcmp1126_pop20_c0_ene5_stall_local = 1'b0;
assign local_bb3_notcmp1126_pop20_c0_ene5_valid_out_0 = 1'b1;
assign local_bb3_notcmp1126_pop20_c0_ene5_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_3 = 1'b0;
assign rnode_1to3_bb3_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_notexitcond1429_pop21_c0_ene6_valid_out_0;
wire local_bb3_notexitcond1429_pop21_c0_ene6_stall_in_0;
wire local_bb3_notexitcond1429_pop21_c0_ene6_valid_out_1;
wire local_bb3_notexitcond1429_pop21_c0_ene6_stall_in_1;
wire local_bb3_notexitcond1429_pop21_c0_ene6_inputs_ready;
wire local_bb3_notexitcond1429_pop21_c0_ene6_stall_local;
wire local_bb3_notexitcond1429_pop21_c0_ene6;
wire local_bb3_notexitcond1429_pop21_c0_ene6_fu_valid_out;
wire local_bb3_notexitcond1429_pop21_c0_ene6_fu_stall_out;

acl_pop local_bb3_notexitcond1429_pop21_c0_ene6_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_3_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene6_0_NO_SHIFT_REG),
	.stall_out(local_bb3_notexitcond1429_pop21_c0_ene6_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notexitcond1429_pop21_c0_ene6_fu_valid_out),
	.stall_in(local_bb3_notexitcond1429_pop21_c0_ene6_stall_local),
	.data_out(local_bb3_notexitcond1429_pop21_c0_ene6),
	.feedback_in(feedback_data_in_21),
	.feedback_valid_in(feedback_valid_in_21),
	.feedback_stall_out(feedback_stall_out_21)
);

defparam local_bb3_notexitcond1429_pop21_c0_ene6_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_notexitcond1429_pop21_c0_ene6_feedback.DATA_WIDTH = 1;
defparam local_bb3_notexitcond1429_pop21_c0_ene6_feedback.STYLE = "REGULAR";

assign local_bb3_notexitcond1429_pop21_c0_ene6_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_4_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene6_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_3_NO_SHIFT_REG);
assign local_bb3_notexitcond1429_pop21_c0_ene6_stall_local = 1'b0;
assign local_bb3_notexitcond1429_pop21_c0_ene6_valid_out_0 = 1'b1;
assign local_bb3_notexitcond1429_pop21_c0_ene6_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_4 = 1'b0;
assign rnode_1to3_bb3_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_valid_out_0;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_stall_in_0;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_valid_out_1;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_stall_in_1;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_inputs_ready;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_stall_local;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_fu_valid_out;
wire local_bb3_memdep_phi1_pop932_pop22_c0_ene7_fu_stall_out;

acl_pop local_bb3_memdep_phi1_pop932_pop22_c0_ene7_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_4_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene7_0_NO_SHIFT_REG),
	.stall_out(local_bb3_memdep_phi1_pop932_pop22_c0_ene7_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_memdep_phi1_pop932_pop22_c0_ene7_fu_valid_out),
	.stall_in(local_bb3_memdep_phi1_pop932_pop22_c0_ene7_stall_local),
	.data_out(local_bb3_memdep_phi1_pop932_pop22_c0_ene7),
	.feedback_in(feedback_data_in_22),
	.feedback_valid_in(feedback_valid_in_22),
	.feedback_stall_out(feedback_stall_out_22)
);

defparam local_bb3_memdep_phi1_pop932_pop22_c0_ene7_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_memdep_phi1_pop932_pop22_c0_ene7_feedback.DATA_WIDTH = 1;
defparam local_bb3_memdep_phi1_pop932_pop22_c0_ene7_feedback.STYLE = "REGULAR";

assign local_bb3_memdep_phi1_pop932_pop22_c0_ene7_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_5_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene7_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_4_NO_SHIFT_REG);
assign local_bb3_memdep_phi1_pop932_pop22_c0_ene7_stall_local = 1'b0;
assign local_bb3_memdep_phi1_pop932_pop22_c0_ene7_valid_out_0 = 1'b1;
assign local_bb3_memdep_phi1_pop932_pop22_c0_ene7_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_5 = 1'b0;
assign rnode_1to3_bb3_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_4_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_valid_out_0;
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_stall_in_0;
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_valid_out_1;
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_stall_in_1;
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_inputs_ready;
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_stall_local;
wire [63:0] local_bb3_indvars_iv_pop1036_pop24_c0_ene8;
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_fu_valid_out;
wire local_bb3_indvars_iv_pop1036_pop24_c0_ene8_fu_stall_out;

acl_pop local_bb3_indvars_iv_pop1036_pop24_c0_ene8_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_5_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene8_0_NO_SHIFT_REG),
	.stall_out(local_bb3_indvars_iv_pop1036_pop24_c0_ene8_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_indvars_iv_pop1036_pop24_c0_ene8_fu_valid_out),
	.stall_in(local_bb3_indvars_iv_pop1036_pop24_c0_ene8_stall_local),
	.data_out(local_bb3_indvars_iv_pop1036_pop24_c0_ene8),
	.feedback_in(feedback_data_in_24),
	.feedback_valid_in(feedback_valid_in_24),
	.feedback_stall_out(feedback_stall_out_24)
);

defparam local_bb3_indvars_iv_pop1036_pop24_c0_ene8_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_indvars_iv_pop1036_pop24_c0_ene8_feedback.DATA_WIDTH = 64;
defparam local_bb3_indvars_iv_pop1036_pop24_c0_ene8_feedback.STYLE = "REGULAR";

assign local_bb3_indvars_iv_pop1036_pop24_c0_ene8_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_6_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene8_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_5_NO_SHIFT_REG);
assign local_bb3_indvars_iv_pop1036_pop24_c0_ene8_stall_local = 1'b0;
assign local_bb3_indvars_iv_pop1036_pop24_c0_ene8_valid_out_0 = 1'b1;
assign local_bb3_indvars_iv_pop1036_pop24_c0_ene8_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_6 = 1'b0;
assign rnode_1to3_bb3_c0_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_5_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__pop25_c0_ene9_valid_out_0;
wire local_bb3__pop25_c0_ene9_stall_in_0;
wire local_bb3__pop25_c0_ene9_valid_out_1;
wire local_bb3__pop25_c0_ene9_stall_in_1;
wire local_bb3__pop25_c0_ene9_inputs_ready;
wire local_bb3__pop25_c0_ene9_stall_local;
wire [31:0] local_bb3__pop25_c0_ene9;
wire local_bb3__pop25_c0_ene9_fu_valid_out;
wire local_bb3__pop25_c0_ene9_fu_stall_out;

acl_pop local_bb3__pop25_c0_ene9_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene9_0_NO_SHIFT_REG),
	.stall_out(local_bb3__pop25_c0_ene9_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3__pop25_c0_ene9_fu_valid_out),
	.stall_in(local_bb3__pop25_c0_ene9_stall_local),
	.data_out(local_bb3__pop25_c0_ene9),
	.feedback_in(feedback_data_in_25),
	.feedback_valid_in(feedback_valid_in_25),
	.feedback_stall_out(feedback_stall_out_25)
);

defparam local_bb3__pop25_c0_ene9_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3__pop25_c0_ene9_feedback.DATA_WIDTH = 32;
defparam local_bb3__pop25_c0_ene9_feedback.STYLE = "REGULAR";

assign local_bb3__pop25_c0_ene9_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_7_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene9_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_6_NO_SHIFT_REG);
assign local_bb3__pop25_c0_ene9_stall_local = 1'b0;
assign local_bb3__pop25_c0_ene9_valid_out_0 = 1'b1;
assign local_bb3__pop25_c0_ene9_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_7 = 1'b0;
assign rnode_1to3_bb3_c0_ene9_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_6_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_valid_out_0;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_stall_in_0;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_valid_out_1;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_stall_in_1;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_inputs_ready;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_stall_local;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_fu_valid_out;
wire local_bb3_memdep_phi1_or38_pop26_c0_ene10_fu_stall_out;

acl_pop local_bb3_memdep_phi1_or38_pop26_c0_ene10_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_7_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene10_0_NO_SHIFT_REG),
	.stall_out(local_bb3_memdep_phi1_or38_pop26_c0_ene10_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_memdep_phi1_or38_pop26_c0_ene10_fu_valid_out),
	.stall_in(local_bb3_memdep_phi1_or38_pop26_c0_ene10_stall_local),
	.data_out(local_bb3_memdep_phi1_or38_pop26_c0_ene10),
	.feedback_in(feedback_data_in_26),
	.feedback_valid_in(feedback_valid_in_26),
	.feedback_stall_out(feedback_stall_out_26)
);

defparam local_bb3_memdep_phi1_or38_pop26_c0_ene10_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_memdep_phi1_or38_pop26_c0_ene10_feedback.DATA_WIDTH = 1;
defparam local_bb3_memdep_phi1_or38_pop26_c0_ene10_feedback.STYLE = "REGULAR";

assign local_bb3_memdep_phi1_or38_pop26_c0_ene10_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_8_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene10_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_7_NO_SHIFT_REG);
assign local_bb3_memdep_phi1_or38_pop26_c0_ene10_stall_local = 1'b0;
assign local_bb3_memdep_phi1_or38_pop26_c0_ene10_valid_out_0 = 1'b1;
assign local_bb3_memdep_phi1_or38_pop26_c0_ene10_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_8 = 1'b0;
assign rnode_1to3_bb3_c0_ene10_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_7_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3__pop27_c0_ene11_valid_out_0;
wire local_bb3__pop27_c0_ene11_stall_in_0;
wire local_bb3__pop27_c0_ene11_valid_out_1;
wire local_bb3__pop27_c0_ene11_stall_in_1;
wire local_bb3__pop27_c0_ene11_inputs_ready;
wire local_bb3__pop27_c0_ene11_stall_local;
wire [31:0] local_bb3__pop27_c0_ene11;
wire local_bb3__pop27_c0_ene11_fu_valid_out;
wire local_bb3__pop27_c0_ene11_fu_stall_out;

acl_pop local_bb3__pop27_c0_ene11_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_8_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene11_0_NO_SHIFT_REG),
	.stall_out(local_bb3__pop27_c0_ene11_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3__pop27_c0_ene11_fu_valid_out),
	.stall_in(local_bb3__pop27_c0_ene11_stall_local),
	.data_out(local_bb3__pop27_c0_ene11),
	.feedback_in(feedback_data_in_27),
	.feedback_valid_in(feedback_valid_in_27),
	.feedback_stall_out(feedback_stall_out_27)
);

defparam local_bb3__pop27_c0_ene11_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3__pop27_c0_ene11_feedback.DATA_WIDTH = 32;
defparam local_bb3__pop27_c0_ene11_feedback.STYLE = "REGULAR";

assign local_bb3__pop27_c0_ene11_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_9_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene11_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_8_NO_SHIFT_REG);
assign local_bb3__pop27_c0_ene11_stall_local = 1'b0;
assign local_bb3__pop27_c0_ene11_valid_out_0 = 1'b1;
assign local_bb3__pop27_c0_ene11_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_9 = 1'b0;
assign rnode_1to3_bb3_c0_ene11_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_8_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_notcmp40_pop28_c0_ene12_valid_out_0;
wire local_bb3_notcmp40_pop28_c0_ene12_stall_in_0;
wire local_bb3_notcmp40_pop28_c0_ene12_valid_out_1;
wire local_bb3_notcmp40_pop28_c0_ene12_stall_in_1;
wire local_bb3_notcmp40_pop28_c0_ene12_inputs_ready;
wire local_bb3_notcmp40_pop28_c0_ene12_stall_local;
wire local_bb3_notcmp40_pop28_c0_ene12;
wire local_bb3_notcmp40_pop28_c0_ene12_fu_valid_out;
wire local_bb3_notcmp40_pop28_c0_ene12_fu_stall_out;

acl_pop local_bb3_notcmp40_pop28_c0_ene12_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_9_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene12_0_NO_SHIFT_REG),
	.stall_out(local_bb3_notcmp40_pop28_c0_ene12_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notcmp40_pop28_c0_ene12_fu_valid_out),
	.stall_in(local_bb3_notcmp40_pop28_c0_ene12_stall_local),
	.data_out(local_bb3_notcmp40_pop28_c0_ene12),
	.feedback_in(feedback_data_in_28),
	.feedback_valid_in(feedback_valid_in_28),
	.feedback_stall_out(feedback_stall_out_28)
);

defparam local_bb3_notcmp40_pop28_c0_ene12_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_notcmp40_pop28_c0_ene12_feedback.DATA_WIDTH = 1;
defparam local_bb3_notcmp40_pop28_c0_ene12_feedback.STYLE = "REGULAR";

assign local_bb3_notcmp40_pop28_c0_ene12_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_10_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene12_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_9_NO_SHIFT_REG);
assign local_bb3_notcmp40_pop28_c0_ene12_stall_local = 1'b0;
assign local_bb3_notcmp40_pop28_c0_ene12_valid_out_0 = 1'b1;
assign local_bb3_notcmp40_pop28_c0_ene12_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_10 = 1'b0;
assign rnode_1to3_bb3_c0_ene12_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_9_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_notexitcond942_pop29_c0_ene13_valid_out_0;
wire local_bb3_notexitcond942_pop29_c0_ene13_stall_in_0;
wire local_bb3_notexitcond942_pop29_c0_ene13_valid_out_1;
wire local_bb3_notexitcond942_pop29_c0_ene13_stall_in_1;
wire local_bb3_notexitcond942_pop29_c0_ene13_inputs_ready;
wire local_bb3_notexitcond942_pop29_c0_ene13_stall_local;
wire local_bb3_notexitcond942_pop29_c0_ene13;
wire local_bb3_notexitcond942_pop29_c0_ene13_fu_valid_out;
wire local_bb3_notexitcond942_pop29_c0_ene13_fu_stall_out;

acl_pop local_bb3_notexitcond942_pop29_c0_ene13_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_2to3_bb3_c0_ene1_10_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_c0_ene13_0_NO_SHIFT_REG),
	.stall_out(local_bb3_notexitcond942_pop29_c0_ene13_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notexitcond942_pop29_c0_ene13_fu_valid_out),
	.stall_in(local_bb3_notexitcond942_pop29_c0_ene13_stall_local),
	.data_out(local_bb3_notexitcond942_pop29_c0_ene13),
	.feedback_in(feedback_data_in_29),
	.feedback_valid_in(feedback_valid_in_29),
	.feedback_stall_out(feedback_stall_out_29)
);

defparam local_bb3_notexitcond942_pop29_c0_ene13_feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_notexitcond942_pop29_c0_ene13_feedback.DATA_WIDTH = 1;
defparam local_bb3_notexitcond942_pop29_c0_ene13_feedback.STYLE = "REGULAR";

assign local_bb3_notexitcond942_pop29_c0_ene13_inputs_ready = (SFC_1_VALID_2_3_0_valid_out_11_NO_SHIFT_REG & rnode_1to3_bb3_c0_ene13_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_c0_ene1_0_valid_out_10_NO_SHIFT_REG);
assign local_bb3_notexitcond942_pop29_c0_ene13_stall_local = 1'b0;
assign local_bb3_notexitcond942_pop29_c0_ene13_valid_out_0 = 1'b1;
assign local_bb3_notexitcond942_pop29_c0_ene13_valid_out_1 = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in_11 = 1'b0;
assign rnode_1to3_bb3_c0_ene13_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_10_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_keep_going4_acl_pipeline_1_NO_SHIFT_REG),
	.data_out(rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_keep_going4_acl_pipeline_1_stall_in = 1'b0;
assign rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG = rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp9_stall_local;
wire local_bb3_cmp9;

assign local_bb3_cmp9 = ($signed(local_bb3_inc34) > $signed(input_r));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_mul534_pop23_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul534_pop23_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul534_pop23_c0_ene2_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_mul534_pop23_c0_ene2_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_mul534_pop23_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG = rnode_4to5_bb3_mul534_pop23_c0_ene2_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_mul534_pop23_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_cmp_i1_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp_i1_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp_i1_i_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp_i1_i_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp_i1_i_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp_i1_i_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp_i1_i_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp_i1_i_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_cmp_i1_i_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_cmp_i1_i_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_cmp_i1_i_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_cmp_i1_i_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_cmp_i1_i_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_cmp_i1_i),
	.data_out(rnode_2to3_bb3_cmp_i1_i_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_cmp_i1_i_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_cmp_i1_i_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_cmp_i1_i_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_cmp_i1_i_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_cmp_i1_i_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp_i1_i_stall_in = 1'b0;
assign rnode_2to3_bb3_cmp_i1_i_0_NO_SHIFT_REG = rnode_2to3_bb3_cmp_i1_i_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_cmp_i1_i_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_cmp_i1_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_cmp1_i3_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp1_i3_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp1_i3_i_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp1_i3_i_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp1_i3_i_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp1_i3_i_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp1_i3_i_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_cmp1_i3_i_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_cmp1_i3_i_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_cmp1_i3_i_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_cmp1_i3_i_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_cmp1_i3_i_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_cmp1_i3_i_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_cmp1_i3_i),
	.data_out(rnode_2to3_bb3_cmp1_i3_i_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_cmp1_i3_i_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_cmp1_i3_i_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_cmp1_i3_i_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_cmp1_i3_i_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_cmp1_i3_i_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp1_i3_i_stall_in = 1'b0;
assign rnode_2to3_bb3_cmp1_i3_i_0_NO_SHIFT_REG = rnode_2to3_bb3_cmp1_i3_i_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_cmp1_i3_i_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_cmp1_i3_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_4_5_0_inputs_ready;
 reg SFC_1_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_4_5_0_stall_in;
wire SFC_1_VALID_4_5_0_output_regs_ready;
 reg SFC_1_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_4_5_0_causedstall;

assign SFC_1_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_1_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_3_4_0_stall_in = 1'b0;
assign SFC_1_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_4_5_0_output_regs_ready)
		begin
			SFC_1_VALID_4_5_0_NO_SHIFT_REG <= SFC_1_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_pixel_y_020_pop820_pop18_c0_ene3),
	.data_out(rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_pixel_y_020_pop820_pop18_c0_ene3_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG = rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_mul3723_pop19_c0_ene4),
	.data_out(rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_mul3723_pop19_c0_ene4_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG = rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_notcmp1126_pop20_c0_ene5),
	.data_out(rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notcmp1126_pop20_c0_ene5_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG = rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_notexitcond1429_pop21_c0_ene6),
	.data_out(rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notexitcond1429_pop21_c0_ene6_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG = rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_memdep_phi1_pop932_pop22_c0_ene7),
	.data_out(rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_memdep_phi1_pop932_pop22_c0_ene7_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG = rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_indvars_iv_pop1036_pop24_c0_ene8),
	.data_out(rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_fifo.DATA_WIDTH = 64;
defparam rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_indvars_iv_pop1036_pop24_c0_ene8_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG = rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3__pop25_c0_ene9_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop25_c0_ene9_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3__pop25_c0_ene9_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop25_c0_ene9_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop25_c0_ene9_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop25_c0_ene9_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3__pop25_c0_ene9_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3__pop25_c0_ene9_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3__pop25_c0_ene9_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3__pop25_c0_ene9),
	.data_out(rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__pop25_c0_ene9_stall_in_1 = 1'b0;
assign rnode_3to4_bb3__pop25_c0_ene9_0_NO_SHIFT_REG = rnode_3to4_bb3__pop25_c0_ene9_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3__pop25_c0_ene9_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3__pop25_c0_ene9_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_memdep_phi1_or38_pop26_c0_ene10),
	.data_out(rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_memdep_phi1_or38_pop26_c0_ene10_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG = rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3__pop27_c0_ene11_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop27_c0_ene11_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3__pop27_c0_ene11_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop27_c0_ene11_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop27_c0_ene11_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3__pop27_c0_ene11_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3__pop27_c0_ene11_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3__pop27_c0_ene11_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3__pop27_c0_ene11_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3__pop27_c0_ene11),
	.data_out(rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__pop27_c0_ene11_stall_in_1 = 1'b0;
assign rnode_3to4_bb3__pop27_c0_ene11_0_NO_SHIFT_REG = rnode_3to4_bb3__pop27_c0_ene11_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3__pop27_c0_ene11_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3__pop27_c0_ene11_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_notcmp40_pop28_c0_ene12),
	.data_out(rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notcmp40_pop28_c0_ene12_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG = rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_notexitcond942_pop29_c0_ene13),
	.data_out(rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notexitcond942_pop29_c0_ene13_stall_in_1 = 1'b0;
assign rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG = rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_keep_going4_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG = rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__stall_local;
wire local_bb3_var_;

assign local_bb3_var_ = (input_wii_var__u12 | local_bb3_cmp9);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_mul534_pop23_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul534_pop23_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul534_pop23_c0_ene2_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_mul534_pop23_c0_ene2_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_mul534_pop23_c0_ene2_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_mul534_pop23_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG = rnode_5to6_bb3_mul534_pop23_c0_ene2_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_mul534_pop23_c0_ene2_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_mul534_pop23_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3__1_stall_local;
wire [31:0] local_bb3__1;

assign local_bb3__1 = (rnode_2to3_bb3_cmp1_i3_i_0_NO_SHIFT_REG ? input_wii_sub22 : rnode_2to3_bb3_add17_0_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_1_VALID_5_6_0_inputs_ready;
 reg SFC_1_VALID_5_6_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_5_6_0_stall_in;
wire SFC_1_VALID_5_6_0_output_regs_ready;
 reg SFC_1_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_5_6_0_causedstall;

assign SFC_1_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_1_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_4_5_0_stall_in = 1'b0;
assign SFC_1_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_5_6_0_output_regs_ready)
		begin
			SFC_1_VALID_5_6_0_NO_SHIFT_REG <= SFC_1_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG = rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_mul3723_pop19_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG = rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG = rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG = rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG = rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_fifo.DATA_WIDTH = 64;
defparam rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG = rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3__pop25_c0_ene9_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop25_c0_ene9_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3__pop25_c0_ene9_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop25_c0_ene9_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop25_c0_ene9_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop25_c0_ene9_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3__pop25_c0_ene9_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3__pop25_c0_ene9_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3__pop25_c0_ene9_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3__pop25_c0_ene9_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3__pop25_c0_ene9_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3__pop25_c0_ene9_0_NO_SHIFT_REG = rnode_4to5_bb3__pop25_c0_ene9_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3__pop25_c0_ene9_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3__pop25_c0_ene9_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG = rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3__pop27_c0_ene11_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop27_c0_ene11_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3__pop27_c0_ene11_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop27_c0_ene11_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop27_c0_ene11_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3__pop27_c0_ene11_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3__pop27_c0_ene11_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3__pop27_c0_ene11_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3__pop27_c0_ene11_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3__pop27_c0_ene11_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3__pop27_c0_ene11_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3__pop27_c0_ene11_0_NO_SHIFT_REG = rnode_4to5_bb3__pop27_c0_ene11_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3__pop27_c0_ene11_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3__pop27_c0_ene11_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_notcmp40_pop28_c0_ene12_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG = rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG = rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_keep_going4_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_NO_SHIFT_REG = rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_inc34_valid_out_1;
wire local_bb3_inc34_stall_in_1;
wire local_bb3_var__valid_out_1;
wire local_bb3_var__stall_in_1;
wire local_bb3_notexit6_valid_out_0;
wire local_bb3_notexit6_stall_in_0;
wire local_bb3_notexit6_valid_out_1;
wire local_bb3_notexit6_stall_in_1;
wire local_bb3_notexit6_inputs_ready;
wire local_bb3_notexit6_stall_local;
wire local_bb3_notexit6;

assign local_bb3_notexit6_inputs_ready = rnode_1to2_bb3_i_211_pop17_add7_0_valid_out_NO_SHIFT_REG;
assign local_bb3_notexit6 = (local_bb3_var_ ^ 1'b1);
assign local_bb3_inc34_valid_out_1 = 1'b1;
assign local_bb3_var__valid_out_1 = 1'b1;
assign local_bb3_notexit6_valid_out_0 = 1'b1;
assign local_bb3_notexit6_valid_out_1 = 1'b1;
assign rnode_1to2_bb3_i_211_pop17_add7_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi1_stall_local;
wire [447:0] local_bb3_c0_exi1;

assign local_bb3_c0_exi1[31:0] = 32'bx;
assign local_bb3_c0_exi1[63:32] = rnode_5to6_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG;
assign local_bb3_c0_exi1[447:64] = 384'bx;

// This section implements an unregistered operation.
// 
wire local_bb3_cond5_i9_i_valid_out;
wire local_bb3_cond5_i9_i_stall_in;
wire local_bb3_cond5_i9_i_inputs_ready;
wire local_bb3_cond5_i9_i_stall_local;
wire [31:0] local_bb3_cond5_i9_i;

assign local_bb3_cond5_i9_i_inputs_ready = (rnode_2to3_bb3_cmp1_i3_i_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_add17_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_cmp_i1_i_0_valid_out_NO_SHIFT_REG);
assign local_bb3_cond5_i9_i = (rnode_2to3_bb3_cmp_i1_i_0_NO_SHIFT_REG ? 32'h0 : local_bb3__1);
assign local_bb3_cond5_i9_i_valid_out = 1'b1;
assign rnode_2to3_bb3_cmp1_i3_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_add17_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_cmp_i1_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG = rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_mul3723_pop19_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG = rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG = rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG = rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG = rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_fifo.DATA_WIDTH = 64;
defparam rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG = rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3__pop25_c0_ene9_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop25_c0_ene9_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3__pop25_c0_ene9_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop25_c0_ene9_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop25_c0_ene9_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop25_c0_ene9_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3__pop25_c0_ene9_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3__pop25_c0_ene9_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3__pop25_c0_ene9_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3__pop25_c0_ene9_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3__pop25_c0_ene9_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3__pop25_c0_ene9_0_NO_SHIFT_REG = rnode_5to6_bb3__pop25_c0_ene9_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3__pop25_c0_ene9_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3__pop25_c0_ene9_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG = rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3__pop27_c0_ene11_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop27_c0_ene11_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3__pop27_c0_ene11_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop27_c0_ene11_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop27_c0_ene11_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3__pop27_c0_ene11_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3__pop27_c0_ene11_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3__pop27_c0_ene11_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3__pop27_c0_ene11_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3__pop27_c0_ene11_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3__pop27_c0_ene11_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3__pop27_c0_ene11_0_NO_SHIFT_REG = rnode_5to6_bb3__pop27_c0_ene11_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3__pop27_c0_ene11_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3__pop27_c0_ene11_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_notcmp40_pop28_c0_ene12_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG = rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG = rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_var__0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_var__0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_var__0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_var__0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_var__0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_var_),
	.data_out(rnode_2to3_bb3_var__0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_var__0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_var__0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_var__0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_var__0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_var__0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__stall_in_1 = 1'b0;
assign rnode_2to3_bb3_var__0_NO_SHIFT_REG = rnode_2to3_bb3_var__0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_var__0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_var__0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb3_notexitcond5_notexit6_inputs_ready;
 reg local_bb3_notexitcond5_notexit6_valid_out_0_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_0;
 reg local_bb3_notexitcond5_notexit6_valid_out_1_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_1;
 reg local_bb3_notexitcond5_notexit6_valid_out_2_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_2;
 reg local_bb3_notexitcond5_notexit6_valid_out_3_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_3;
 reg local_bb3_notexitcond5_notexit6_valid_out_4_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_4;
 reg local_bb3_notexitcond5_notexit6_valid_out_5_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_5;
 reg local_bb3_notexitcond5_notexit6_valid_out_6_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_6;
 reg local_bb3_notexitcond5_notexit6_valid_out_7_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_7;
 reg local_bb3_notexitcond5_notexit6_valid_out_8_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_8;
 reg local_bb3_notexitcond5_notexit6_valid_out_9_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_9;
 reg local_bb3_notexitcond5_notexit6_valid_out_10_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_10;
 reg local_bb3_notexitcond5_notexit6_valid_out_11_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_11;
 reg local_bb3_notexitcond5_notexit6_valid_out_12_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_stall_in_12;
wire local_bb3_notexitcond5_notexit6_output_regs_ready;
wire local_bb3_notexitcond5_notexit6_result;
wire local_bb3_notexitcond5_notexit6_fu_valid_out;
wire local_bb3_notexitcond5_notexit6_fu_stall_out;
 reg local_bb3_notexitcond5_notexit6_NO_SHIFT_REG;
wire local_bb3_notexitcond5_notexit6_causedstall;

acl_push local_bb3_notexitcond5_notexit6_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(local_bb3_notexit6),
	.stall_out(local_bb3_notexitcond5_notexit6_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notexitcond5_notexit6_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_notexitcond5_notexit6_result),
	.feedback_out(feedback_data_out_3),
	.feedback_valid_out(feedback_valid_out_3),
	.feedback_stall_in(feedback_stall_in_3)
);

defparam local_bb3_notexitcond5_notexit6_feedback.STALLFREE = 1;
defparam local_bb3_notexitcond5_notexit6_feedback.DATA_WIDTH = 1;
defparam local_bb3_notexitcond5_notexit6_feedback.FIFO_DEPTH = 1;
defparam local_bb3_notexitcond5_notexit6_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb3_notexitcond5_notexit6_feedback.STYLE = "REGULAR";

assign local_bb3_notexitcond5_notexit6_inputs_ready = 1'b1;
assign local_bb3_notexitcond5_notexit6_output_regs_ready = 1'b1;
assign local_bb3_notexit6_stall_in_0 = 1'b0;
assign SFC_1_VALID_1_2_0_stall_in_2 = 1'b0;
assign local_bb3_notexitcond5_notexit6_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_notexitcond5_notexit6_NO_SHIFT_REG <= 'x;
		local_bb3_notexitcond5_notexit6_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_7_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_8_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_9_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_10_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_11_NO_SHIFT_REG <= 1'b0;
		local_bb3_notexitcond5_notexit6_valid_out_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_notexitcond5_notexit6_output_regs_ready)
		begin
			local_bb3_notexitcond5_notexit6_NO_SHIFT_REG <= local_bb3_notexitcond5_notexit6_result;
			local_bb3_notexitcond5_notexit6_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_6_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_7_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_8_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_9_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_10_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_11_NO_SHIFT_REG <= 1'b1;
			local_bb3_notexitcond5_notexit6_valid_out_12_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_notexitcond5_notexit6_stall_in_0))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_1))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_2))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_3))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_4))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_5))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_6))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_7))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_8))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_9))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_9_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_10))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_10_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_11))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_11_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_notexitcond5_notexit6_stall_in_12))
			begin
				local_bb3_notexitcond5_notexit6_valid_out_12_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_i_211_push17_inc34_inputs_ready;
 reg local_bb3_i_211_push17_inc34_valid_out_NO_SHIFT_REG;
wire local_bb3_i_211_push17_inc34_stall_in;
wire local_bb3_i_211_push17_inc34_output_regs_ready;
wire [31:0] local_bb3_i_211_push17_inc34_result;
wire local_bb3_i_211_push17_inc34_fu_valid_out;
wire local_bb3_i_211_push17_inc34_fu_stall_out;
 reg [31:0] local_bb3_i_211_push17_inc34_NO_SHIFT_REG;
wire local_bb3_i_211_push17_inc34_causedstall;

acl_push local_bb3_i_211_push17_inc34_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexit6),
	.predicate(1'b0),
	.data_in(local_bb3_inc34),
	.stall_out(local_bb3_i_211_push17_inc34_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_i_211_push17_inc34_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_i_211_push17_inc34_result),
	.feedback_out(feedback_data_out_17),
	.feedback_valid_out(feedback_valid_out_17),
	.feedback_stall_in(feedback_stall_in_17)
);

defparam local_bb3_i_211_push17_inc34_feedback.STALLFREE = 1;
defparam local_bb3_i_211_push17_inc34_feedback.DATA_WIDTH = 32;
defparam local_bb3_i_211_push17_inc34_feedback.FIFO_DEPTH = 2;
defparam local_bb3_i_211_push17_inc34_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb3_i_211_push17_inc34_feedback.STYLE = "REGULAR";

assign local_bb3_i_211_push17_inc34_inputs_ready = 1'b1;
assign local_bb3_i_211_push17_inc34_output_regs_ready = 1'b1;
assign local_bb3_inc34_stall_in_1 = 1'b0;
assign local_bb3_notexit6_stall_in_1 = 1'b0;
assign SFC_1_VALID_1_2_0_stall_in_3 = 1'b0;
assign local_bb3_i_211_push17_inc34_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_i_211_push17_inc34_NO_SHIFT_REG <= 'x;
		local_bb3_i_211_push17_inc34_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_i_211_push17_inc34_output_regs_ready)
		begin
			local_bb3_i_211_push17_inc34_NO_SHIFT_REG <= local_bb3_i_211_push17_inc34_result;
			local_bb3_i_211_push17_inc34_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_i_211_push17_inc34_stall_in))
			begin
				local_bb3_i_211_push17_inc34_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_mul24_inputs_ready;
 reg local_bb3_mul24_valid_out_NO_SHIFT_REG;
wire local_bb3_mul24_stall_in;
wire local_bb3_mul24_output_regs_ready;
wire [31:0] local_bb3_mul24;
 reg local_bb3_mul24_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_mul24_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_mul24_causedstall;

acl_int_mult int_module_local_bb3_mul24 (
	.clock(clock),
	.dataa(local_bb3_cond5_i9_i),
	.datab(input_inSize_x),
	.enable(local_bb3_mul24_output_regs_ready),
	.result(local_bb3_mul24)
);

defparam int_module_local_bb3_mul24.INPUT1_WIDTH = 32;
defparam int_module_local_bb3_mul24.INPUT2_WIDTH = 32;
defparam int_module_local_bb3_mul24.OUTPUT_WIDTH = 32;
defparam int_module_local_bb3_mul24.LATENCY = 3;
defparam int_module_local_bb3_mul24.SIGNED = 0;

assign local_bb3_mul24_inputs_ready = 1'b1;
assign local_bb3_mul24_output_regs_ready = 1'b1;
assign local_bb3_cond5_i9_i_stall_in = 1'b0;
assign local_bb3_mul24_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul24_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul24_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul24_output_regs_ready)
		begin
			local_bb3_mul24_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb3_mul24_valid_pipe_1_NO_SHIFT_REG <= local_bb3_mul24_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul24_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul24_output_regs_ready)
		begin
			local_bb3_mul24_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_mul24_stall_in))
			begin
				local_bb3_mul24_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb3_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb3_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_3to5_bb3_var__0_NO_SHIFT_REG;
 logic rnode_3to5_bb3_var__0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to5_bb3_var__0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_var__0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_var__0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_var__0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb3_var__0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb3_var__0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb3_var__0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb3_var__0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb3_var__0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_2to3_bb3_var__0_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb3_var__0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb3_var__0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb3_var__0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_3to5_bb3_var__0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb3_var__0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb3_var__0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_var__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_var__0_NO_SHIFT_REG = rnode_3to5_bb3_var__0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb3_var__0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_var__0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb3_mul534_push23_mul534_pop23_inputs_ready;
 reg local_bb3_mul534_push23_mul534_pop23_valid_out_NO_SHIFT_REG;
wire local_bb3_mul534_push23_mul534_pop23_stall_in;
wire local_bb3_mul534_push23_mul534_pop23_output_regs_ready;
wire [31:0] local_bb3_mul534_push23_mul534_pop23_result;
wire local_bb3_mul534_push23_mul534_pop23_fu_valid_out;
wire local_bb3_mul534_push23_mul534_pop23_fu_stall_out;
 reg [31:0] local_bb3_mul534_push23_mul534_pop23_NO_SHIFT_REG;
wire local_bb3_mul534_push23_mul534_pop23_causedstall;

acl_push local_bb3_mul534_push23_mul534_pop23_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_1to3_bb3_mul534_pop23_c0_ene2_0_NO_SHIFT_REG),
	.stall_out(local_bb3_mul534_push23_mul534_pop23_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_mul534_push23_mul534_pop23_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_mul534_push23_mul534_pop23_result),
	.feedback_out(feedback_data_out_23),
	.feedback_valid_out(feedback_valid_out_23),
	.feedback_stall_in(feedback_stall_in_23)
);

defparam local_bb3_mul534_push23_mul534_pop23_feedback.STALLFREE = 1;
defparam local_bb3_mul534_push23_mul534_pop23_feedback.DATA_WIDTH = 32;
defparam local_bb3_mul534_push23_mul534_pop23_feedback.FIFO_DEPTH = 2;
defparam local_bb3_mul534_push23_mul534_pop23_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb3_mul534_push23_mul534_pop23_feedback.STYLE = "REGULAR";

assign local_bb3_mul534_push23_mul534_pop23_inputs_ready = 1'b1;
assign local_bb3_mul534_push23_mul534_pop23_output_regs_ready = 1'b1;
assign local_bb3_notexitcond5_notexit6_stall_in_0 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_12 = 1'b0;
assign rnode_1to3_bb3_mul534_pop23_c0_ene2_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb3_mul534_push23_mul534_pop23_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul534_push23_mul534_pop23_NO_SHIFT_REG <= 'x;
		local_bb3_mul534_push23_mul534_pop23_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul534_push23_mul534_pop23_output_regs_ready)
		begin
			local_bb3_mul534_push23_mul534_pop23_NO_SHIFT_REG <= local_bb3_mul534_push23_mul534_pop23_result;
			local_bb3_mul534_push23_mul534_pop23_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_mul534_push23_mul534_pop23_stall_in))
			begin
				local_bb3_mul534_push23_mul534_pop23_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_inputs_ready;
 reg local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_valid_out_NO_SHIFT_REG;
wire local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_stall_in;
wire local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_output_regs_ready;
wire [31:0] local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_result;
wire local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_fu_valid_out;
wire local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_fu_stall_out;
 reg [31:0] local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_NO_SHIFT_REG;
wire local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_causedstall;

acl_push local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_pixel_y_020_pop820_pop18_c0_ene3),
	.stall_out(local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_result),
	.feedback_out(feedback_data_out_18),
	.feedback_valid_out(feedback_valid_out_18),
	.feedback_stall_in(feedback_stall_in_18)
);

defparam local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_feedback.STALLFREE = 1;
defparam local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_feedback.DATA_WIDTH = 32;
defparam local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_feedback.FIFO_DEPTH = 2;
defparam local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_feedback.STYLE = "REGULAR";

assign local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_inputs_ready = 1'b1;
assign local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_output_regs_ready = 1'b1;
assign local_bb3_pixel_y_020_pop820_pop18_c0_ene3_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_1 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_13 = 1'b0;
assign local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_NO_SHIFT_REG <= 'x;
		local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_output_regs_ready)
		begin
			local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_NO_SHIFT_REG <= local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_result;
			local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_stall_in))
			begin
				local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_mul3723_push19_mul3723_pop19_inputs_ready;
 reg local_bb3_mul3723_push19_mul3723_pop19_valid_out_NO_SHIFT_REG;
wire local_bb3_mul3723_push19_mul3723_pop19_stall_in;
wire local_bb3_mul3723_push19_mul3723_pop19_output_regs_ready;
wire [31:0] local_bb3_mul3723_push19_mul3723_pop19_result;
wire local_bb3_mul3723_push19_mul3723_pop19_fu_valid_out;
wire local_bb3_mul3723_push19_mul3723_pop19_fu_stall_out;
 reg [31:0] local_bb3_mul3723_push19_mul3723_pop19_NO_SHIFT_REG;
wire local_bb3_mul3723_push19_mul3723_pop19_causedstall;

acl_push local_bb3_mul3723_push19_mul3723_pop19_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_mul3723_pop19_c0_ene4),
	.stall_out(local_bb3_mul3723_push19_mul3723_pop19_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_mul3723_push19_mul3723_pop19_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_mul3723_push19_mul3723_pop19_result),
	.feedback_out(feedback_data_out_19),
	.feedback_valid_out(feedback_valid_out_19),
	.feedback_stall_in(feedback_stall_in_19)
);

defparam local_bb3_mul3723_push19_mul3723_pop19_feedback.STALLFREE = 1;
defparam local_bb3_mul3723_push19_mul3723_pop19_feedback.DATA_WIDTH = 32;
defparam local_bb3_mul3723_push19_mul3723_pop19_feedback.FIFO_DEPTH = 2;
defparam local_bb3_mul3723_push19_mul3723_pop19_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_mul3723_push19_mul3723_pop19_feedback.STYLE = "REGULAR";

assign local_bb3_mul3723_push19_mul3723_pop19_inputs_ready = 1'b1;
assign local_bb3_mul3723_push19_mul3723_pop19_output_regs_ready = 1'b1;
assign local_bb3_mul3723_pop19_c0_ene4_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_2 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_14 = 1'b0;
assign local_bb3_mul3723_push19_mul3723_pop19_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul3723_push19_mul3723_pop19_NO_SHIFT_REG <= 'x;
		local_bb3_mul3723_push19_mul3723_pop19_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul3723_push19_mul3723_pop19_output_regs_ready)
		begin
			local_bb3_mul3723_push19_mul3723_pop19_NO_SHIFT_REG <= local_bb3_mul3723_push19_mul3723_pop19_result;
			local_bb3_mul3723_push19_mul3723_pop19_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_mul3723_push19_mul3723_pop19_stall_in))
			begin
				local_bb3_mul3723_push19_mul3723_pop19_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_notcmp1126_push20_notcmp1126_pop20_inputs_ready;
 reg local_bb3_notcmp1126_push20_notcmp1126_pop20_valid_out_NO_SHIFT_REG;
wire local_bb3_notcmp1126_push20_notcmp1126_pop20_stall_in;
wire local_bb3_notcmp1126_push20_notcmp1126_pop20_output_regs_ready;
wire local_bb3_notcmp1126_push20_notcmp1126_pop20_result;
wire local_bb3_notcmp1126_push20_notcmp1126_pop20_fu_valid_out;
wire local_bb3_notcmp1126_push20_notcmp1126_pop20_fu_stall_out;
 reg local_bb3_notcmp1126_push20_notcmp1126_pop20_NO_SHIFT_REG;
wire local_bb3_notcmp1126_push20_notcmp1126_pop20_causedstall;

acl_push local_bb3_notcmp1126_push20_notcmp1126_pop20_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_notcmp1126_pop20_c0_ene5),
	.stall_out(local_bb3_notcmp1126_push20_notcmp1126_pop20_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notcmp1126_push20_notcmp1126_pop20_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_notcmp1126_push20_notcmp1126_pop20_result),
	.feedback_out(feedback_data_out_20),
	.feedback_valid_out(feedback_valid_out_20),
	.feedback_stall_in(feedback_stall_in_20)
);

defparam local_bb3_notcmp1126_push20_notcmp1126_pop20_feedback.STALLFREE = 1;
defparam local_bb3_notcmp1126_push20_notcmp1126_pop20_feedback.DATA_WIDTH = 1;
defparam local_bb3_notcmp1126_push20_notcmp1126_pop20_feedback.FIFO_DEPTH = 2;
defparam local_bb3_notcmp1126_push20_notcmp1126_pop20_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_notcmp1126_push20_notcmp1126_pop20_feedback.STYLE = "REGULAR";

assign local_bb3_notcmp1126_push20_notcmp1126_pop20_inputs_ready = 1'b1;
assign local_bb3_notcmp1126_push20_notcmp1126_pop20_output_regs_ready = 1'b1;
assign local_bb3_notcmp1126_pop20_c0_ene5_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_3 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_15 = 1'b0;
assign local_bb3_notcmp1126_push20_notcmp1126_pop20_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_notcmp1126_push20_notcmp1126_pop20_NO_SHIFT_REG <= 'x;
		local_bb3_notcmp1126_push20_notcmp1126_pop20_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_notcmp1126_push20_notcmp1126_pop20_output_regs_ready)
		begin
			local_bb3_notcmp1126_push20_notcmp1126_pop20_NO_SHIFT_REG <= local_bb3_notcmp1126_push20_notcmp1126_pop20_result;
			local_bb3_notcmp1126_push20_notcmp1126_pop20_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_notcmp1126_push20_notcmp1126_pop20_stall_in))
			begin
				local_bb3_notcmp1126_push20_notcmp1126_pop20_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_notexitcond1429_push21_notexitcond1429_pop21_inputs_ready;
 reg local_bb3_notexitcond1429_push21_notexitcond1429_pop21_valid_out_NO_SHIFT_REG;
wire local_bb3_notexitcond1429_push21_notexitcond1429_pop21_stall_in;
wire local_bb3_notexitcond1429_push21_notexitcond1429_pop21_output_regs_ready;
wire local_bb3_notexitcond1429_push21_notexitcond1429_pop21_result;
wire local_bb3_notexitcond1429_push21_notexitcond1429_pop21_fu_valid_out;
wire local_bb3_notexitcond1429_push21_notexitcond1429_pop21_fu_stall_out;
 reg local_bb3_notexitcond1429_push21_notexitcond1429_pop21_NO_SHIFT_REG;
wire local_bb3_notexitcond1429_push21_notexitcond1429_pop21_causedstall;

acl_push local_bb3_notexitcond1429_push21_notexitcond1429_pop21_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_notexitcond1429_pop21_c0_ene6),
	.stall_out(local_bb3_notexitcond1429_push21_notexitcond1429_pop21_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notexitcond1429_push21_notexitcond1429_pop21_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_notexitcond1429_push21_notexitcond1429_pop21_result),
	.feedback_out(feedback_data_out_21),
	.feedback_valid_out(feedback_valid_out_21),
	.feedback_stall_in(feedback_stall_in_21)
);

defparam local_bb3_notexitcond1429_push21_notexitcond1429_pop21_feedback.STALLFREE = 1;
defparam local_bb3_notexitcond1429_push21_notexitcond1429_pop21_feedback.DATA_WIDTH = 1;
defparam local_bb3_notexitcond1429_push21_notexitcond1429_pop21_feedback.FIFO_DEPTH = 2;
defparam local_bb3_notexitcond1429_push21_notexitcond1429_pop21_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_notexitcond1429_push21_notexitcond1429_pop21_feedback.STYLE = "REGULAR";

assign local_bb3_notexitcond1429_push21_notexitcond1429_pop21_inputs_ready = 1'b1;
assign local_bb3_notexitcond1429_push21_notexitcond1429_pop21_output_regs_ready = 1'b1;
assign local_bb3_notexitcond1429_pop21_c0_ene6_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_4 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_16 = 1'b0;
assign local_bb3_notexitcond1429_push21_notexitcond1429_pop21_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_notexitcond1429_push21_notexitcond1429_pop21_NO_SHIFT_REG <= 'x;
		local_bb3_notexitcond1429_push21_notexitcond1429_pop21_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_notexitcond1429_push21_notexitcond1429_pop21_output_regs_ready)
		begin
			local_bb3_notexitcond1429_push21_notexitcond1429_pop21_NO_SHIFT_REG <= local_bb3_notexitcond1429_push21_notexitcond1429_pop21_result;
			local_bb3_notexitcond1429_push21_notexitcond1429_pop21_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_notexitcond1429_push21_notexitcond1429_pop21_stall_in))
			begin
				local_bb3_notexitcond1429_push21_notexitcond1429_pop21_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_inputs_ready;
 reg local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_valid_out_NO_SHIFT_REG;
wire local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_stall_in;
wire local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_output_regs_ready;
wire local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_result;
wire local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_fu_valid_out;
wire local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_fu_stall_out;
 reg local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_NO_SHIFT_REG;
wire local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_causedstall;

acl_push local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_memdep_phi1_pop932_pop22_c0_ene7),
	.stall_out(local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_result),
	.feedback_out(feedback_data_out_22),
	.feedback_valid_out(feedback_valid_out_22),
	.feedback_stall_in(feedback_stall_in_22)
);

defparam local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_feedback.STALLFREE = 1;
defparam local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_feedback.DATA_WIDTH = 1;
defparam local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_feedback.FIFO_DEPTH = 2;
defparam local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_feedback.STYLE = "REGULAR";

assign local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_inputs_ready = 1'b1;
assign local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_output_regs_ready = 1'b1;
assign local_bb3_memdep_phi1_pop932_pop22_c0_ene7_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_5 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_17 = 1'b0;
assign local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_NO_SHIFT_REG <= 'x;
		local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_output_regs_ready)
		begin
			local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_NO_SHIFT_REG <= local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_result;
			local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_stall_in))
			begin
				local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_inputs_ready;
 reg local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_valid_out_NO_SHIFT_REG;
wire local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_stall_in;
wire local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_output_regs_ready;
wire [63:0] local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_result;
wire local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_fu_valid_out;
wire local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_fu_stall_out;
 reg [63:0] local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_NO_SHIFT_REG;
wire local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_causedstall;

acl_push local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_indvars_iv_pop1036_pop24_c0_ene8),
	.stall_out(local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_result),
	.feedback_out(feedback_data_out_24),
	.feedback_valid_out(feedback_valid_out_24),
	.feedback_stall_in(feedback_stall_in_24)
);

defparam local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_feedback.STALLFREE = 1;
defparam local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_feedback.DATA_WIDTH = 64;
defparam local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_feedback.FIFO_DEPTH = 2;
defparam local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_feedback.STYLE = "REGULAR";

assign local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_inputs_ready = 1'b1;
assign local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_output_regs_ready = 1'b1;
assign local_bb3_indvars_iv_pop1036_pop24_c0_ene8_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_6 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_18 = 1'b0;
assign local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_NO_SHIFT_REG <= 'x;
		local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_output_regs_ready)
		begin
			local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_NO_SHIFT_REG <= local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_result;
			local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_stall_in))
			begin
				local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3__push25__pop25_inputs_ready;
 reg local_bb3__push25__pop25_valid_out_NO_SHIFT_REG;
wire local_bb3__push25__pop25_stall_in;
wire local_bb3__push25__pop25_output_regs_ready;
wire [31:0] local_bb3__push25__pop25_result;
wire local_bb3__push25__pop25_fu_valid_out;
wire local_bb3__push25__pop25_fu_stall_out;
 reg [31:0] local_bb3__push25__pop25_NO_SHIFT_REG;
wire local_bb3__push25__pop25_causedstall;

acl_push local_bb3__push25__pop25_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3__pop25_c0_ene9),
	.stall_out(local_bb3__push25__pop25_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3__push25__pop25_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3__push25__pop25_result),
	.feedback_out(feedback_data_out_25),
	.feedback_valid_out(feedback_valid_out_25),
	.feedback_stall_in(feedback_stall_in_25)
);

defparam local_bb3__push25__pop25_feedback.STALLFREE = 1;
defparam local_bb3__push25__pop25_feedback.DATA_WIDTH = 32;
defparam local_bb3__push25__pop25_feedback.FIFO_DEPTH = 2;
defparam local_bb3__push25__pop25_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3__push25__pop25_feedback.STYLE = "REGULAR";

assign local_bb3__push25__pop25_inputs_ready = 1'b1;
assign local_bb3__push25__pop25_output_regs_ready = 1'b1;
assign local_bb3__pop25_c0_ene9_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_7 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_19 = 1'b0;
assign local_bb3__push25__pop25_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3__push25__pop25_NO_SHIFT_REG <= 'x;
		local_bb3__push25__pop25_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3__push25__pop25_output_regs_ready)
		begin
			local_bb3__push25__pop25_NO_SHIFT_REG <= local_bb3__push25__pop25_result;
			local_bb3__push25__pop25_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3__push25__pop25_stall_in))
			begin
				local_bb3__push25__pop25_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_inputs_ready;
 reg local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_valid_out_NO_SHIFT_REG;
wire local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_stall_in;
wire local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_output_regs_ready;
wire local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_result;
wire local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_fu_valid_out;
wire local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_fu_stall_out;
 reg local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_NO_SHIFT_REG;
wire local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_causedstall;

acl_push local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_memdep_phi1_or38_pop26_c0_ene10),
	.stall_out(local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_result),
	.feedback_out(feedback_data_out_26),
	.feedback_valid_out(feedback_valid_out_26),
	.feedback_stall_in(feedback_stall_in_26)
);

defparam local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_feedback.STALLFREE = 1;
defparam local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_feedback.DATA_WIDTH = 1;
defparam local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_feedback.FIFO_DEPTH = 2;
defparam local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_feedback.STYLE = "REGULAR";

assign local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_inputs_ready = 1'b1;
assign local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_output_regs_ready = 1'b1;
assign local_bb3_memdep_phi1_or38_pop26_c0_ene10_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_8 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_20 = 1'b0;
assign local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_NO_SHIFT_REG <= 'x;
		local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_output_regs_ready)
		begin
			local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_NO_SHIFT_REG <= local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_result;
			local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_stall_in))
			begin
				local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3__push27__pop27_inputs_ready;
 reg local_bb3__push27__pop27_valid_out_NO_SHIFT_REG;
wire local_bb3__push27__pop27_stall_in;
wire local_bb3__push27__pop27_output_regs_ready;
wire [31:0] local_bb3__push27__pop27_result;
wire local_bb3__push27__pop27_fu_valid_out;
wire local_bb3__push27__pop27_fu_stall_out;
 reg [31:0] local_bb3__push27__pop27_NO_SHIFT_REG;
wire local_bb3__push27__pop27_causedstall;

acl_push local_bb3__push27__pop27_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3__pop27_c0_ene11),
	.stall_out(local_bb3__push27__pop27_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3__push27__pop27_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3__push27__pop27_result),
	.feedback_out(feedback_data_out_27),
	.feedback_valid_out(feedback_valid_out_27),
	.feedback_stall_in(feedback_stall_in_27)
);

defparam local_bb3__push27__pop27_feedback.STALLFREE = 1;
defparam local_bb3__push27__pop27_feedback.DATA_WIDTH = 32;
defparam local_bb3__push27__pop27_feedback.FIFO_DEPTH = 2;
defparam local_bb3__push27__pop27_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3__push27__pop27_feedback.STYLE = "REGULAR";

assign local_bb3__push27__pop27_inputs_ready = 1'b1;
assign local_bb3__push27__pop27_output_regs_ready = 1'b1;
assign local_bb3__pop27_c0_ene11_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_9 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_21 = 1'b0;
assign local_bb3__push27__pop27_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3__push27__pop27_NO_SHIFT_REG <= 'x;
		local_bb3__push27__pop27_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3__push27__pop27_output_regs_ready)
		begin
			local_bb3__push27__pop27_NO_SHIFT_REG <= local_bb3__push27__pop27_result;
			local_bb3__push27__pop27_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3__push27__pop27_stall_in))
			begin
				local_bb3__push27__pop27_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_notcmp40_push28_notcmp40_pop28_inputs_ready;
 reg local_bb3_notcmp40_push28_notcmp40_pop28_valid_out_NO_SHIFT_REG;
wire local_bb3_notcmp40_push28_notcmp40_pop28_stall_in;
wire local_bb3_notcmp40_push28_notcmp40_pop28_output_regs_ready;
wire local_bb3_notcmp40_push28_notcmp40_pop28_result;
wire local_bb3_notcmp40_push28_notcmp40_pop28_fu_valid_out;
wire local_bb3_notcmp40_push28_notcmp40_pop28_fu_stall_out;
 reg local_bb3_notcmp40_push28_notcmp40_pop28_NO_SHIFT_REG;
wire local_bb3_notcmp40_push28_notcmp40_pop28_causedstall;

acl_push local_bb3_notcmp40_push28_notcmp40_pop28_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_notcmp40_pop28_c0_ene12),
	.stall_out(local_bb3_notcmp40_push28_notcmp40_pop28_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notcmp40_push28_notcmp40_pop28_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_notcmp40_push28_notcmp40_pop28_result),
	.feedback_out(feedback_data_out_28),
	.feedback_valid_out(feedback_valid_out_28),
	.feedback_stall_in(feedback_stall_in_28)
);

defparam local_bb3_notcmp40_push28_notcmp40_pop28_feedback.STALLFREE = 1;
defparam local_bb3_notcmp40_push28_notcmp40_pop28_feedback.DATA_WIDTH = 1;
defparam local_bb3_notcmp40_push28_notcmp40_pop28_feedback.FIFO_DEPTH = 2;
defparam local_bb3_notcmp40_push28_notcmp40_pop28_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_notcmp40_push28_notcmp40_pop28_feedback.STYLE = "REGULAR";

assign local_bb3_notcmp40_push28_notcmp40_pop28_inputs_ready = 1'b1;
assign local_bb3_notcmp40_push28_notcmp40_pop28_output_regs_ready = 1'b1;
assign local_bb3_notcmp40_pop28_c0_ene12_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_10 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_22 = 1'b0;
assign local_bb3_notcmp40_push28_notcmp40_pop28_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_notcmp40_push28_notcmp40_pop28_NO_SHIFT_REG <= 'x;
		local_bb3_notcmp40_push28_notcmp40_pop28_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_notcmp40_push28_notcmp40_pop28_output_regs_ready)
		begin
			local_bb3_notcmp40_push28_notcmp40_pop28_NO_SHIFT_REG <= local_bb3_notcmp40_push28_notcmp40_pop28_result;
			local_bb3_notcmp40_push28_notcmp40_pop28_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_notcmp40_push28_notcmp40_pop28_stall_in))
			begin
				local_bb3_notcmp40_push28_notcmp40_pop28_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_notexitcond942_push29_notexitcond942_pop29_inputs_ready;
 reg local_bb3_notexitcond942_push29_notexitcond942_pop29_valid_out_NO_SHIFT_REG;
wire local_bb3_notexitcond942_push29_notexitcond942_pop29_stall_in;
wire local_bb3_notexitcond942_push29_notexitcond942_pop29_output_regs_ready;
wire local_bb3_notexitcond942_push29_notexitcond942_pop29_result;
wire local_bb3_notexitcond942_push29_notexitcond942_pop29_fu_valid_out;
wire local_bb3_notexitcond942_push29_notexitcond942_pop29_fu_stall_out;
 reg local_bb3_notexitcond942_push29_notexitcond942_pop29_NO_SHIFT_REG;
wire local_bb3_notexitcond942_push29_notexitcond942_pop29_causedstall;

acl_push local_bb3_notexitcond942_push29_notexitcond942_pop29_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb3_notexitcond942_pop29_c0_ene13),
	.stall_out(local_bb3_notexitcond942_push29_notexitcond942_pop29_fu_stall_out),
	.valid_in(SFC_1_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notexitcond942_push29_notexitcond942_pop29_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_notexitcond942_push29_notexitcond942_pop29_result),
	.feedback_out(feedback_data_out_29),
	.feedback_valid_out(feedback_valid_out_29),
	.feedback_stall_in(feedback_stall_in_29)
);

defparam local_bb3_notexitcond942_push29_notexitcond942_pop29_feedback.STALLFREE = 1;
defparam local_bb3_notexitcond942_push29_notexitcond942_pop29_feedback.DATA_WIDTH = 1;
defparam local_bb3_notexitcond942_push29_notexitcond942_pop29_feedback.FIFO_DEPTH = 2;
defparam local_bb3_notexitcond942_push29_notexitcond942_pop29_feedback.MIN_FIFO_LATENCY = 2;
defparam local_bb3_notexitcond942_push29_notexitcond942_pop29_feedback.STYLE = "REGULAR";

assign local_bb3_notexitcond942_push29_notexitcond942_pop29_inputs_ready = 1'b1;
assign local_bb3_notexitcond942_push29_notexitcond942_pop29_output_regs_ready = 1'b1;
assign local_bb3_notexitcond942_pop29_c0_ene13_stall_in_0 = 1'b0;
assign local_bb3_notexitcond5_notexit6_stall_in_11 = 1'b0;
assign SFC_1_VALID_2_3_0_stall_in_23 = 1'b0;
assign local_bb3_notexitcond942_push29_notexitcond942_pop29_causedstall = (SFC_1_VALID_2_3_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_notexitcond942_push29_notexitcond942_pop29_NO_SHIFT_REG <= 'x;
		local_bb3_notexitcond942_push29_notexitcond942_pop29_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_notexitcond942_push29_notexitcond942_pop29_output_regs_ready)
		begin
			local_bb3_notexitcond942_push29_notexitcond942_pop29_NO_SHIFT_REG <= local_bb3_notexitcond942_push29_notexitcond942_pop29_result;
			local_bb3_notexitcond942_push29_notexitcond942_pop29_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_notexitcond942_push29_notexitcond942_pop29_stall_in))
			begin
				local_bb3_notexitcond942_push29_notexitcond942_pop29_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_notexitcond5_notexit6_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_notexitcond5_notexit6_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_notexitcond5_notexit6_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_notexitcond5_notexit6_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_notexitcond5_notexit6_NO_SHIFT_REG),
	.data_out(rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notexitcond5_notexit6_stall_in_12 = 1'b0;
assign rnode_3to4_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG = rnode_3to4_bb3_notexitcond5_notexit6_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_notexitcond5_notexit6_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_notexitcond5_notexit6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_i_211_push17_inc34_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_i_211_push17_inc34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_i_211_push17_inc34_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_i_211_push17_inc34_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_i_211_push17_inc34_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_i_211_push17_inc34_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_i_211_push17_inc34_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_i_211_push17_inc34_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_i_211_push17_inc34_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_i_211_push17_inc34_NO_SHIFT_REG),
	.data_out(rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_i_211_push17_inc34_stall_in = 1'b0;
assign rnode_3to4_bb3_i_211_push17_inc34_0_NO_SHIFT_REG = rnode_3to4_bb3_i_211_push17_inc34_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_i_211_push17_inc34_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_i_211_push17_inc34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi2_stall_local;
wire [447:0] local_bb3_c0_exi2;

assign local_bb3_c0_exi2[63:0] = local_bb3_c0_exi1[63:0];
assign local_bb3_c0_exi2[95:64] = local_bb3_mul24;
assign local_bb3_c0_exi2[447:96] = local_bb3_c0_exi1[447:96];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_var__0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_var__0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_var__0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_var__0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_var__0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_var__0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_var__0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_var__0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_var__0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_var__0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_var__0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_3to5_bb3_var__0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_var__0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_var__0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_var__0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_var__0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_var__0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_var__0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to5_bb3_var__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_var__0_NO_SHIFT_REG = rnode_5to6_bb3_var__0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_var__0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_var__0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_mul534_push23_mul534_pop23_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul534_push23_mul534_pop23_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3_mul534_push23_mul534_pop23_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul534_push23_mul534_pop23_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul534_push23_mul534_pop23_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul534_push23_mul534_pop23_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_mul534_push23_mul534_pop23_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_mul534_push23_mul534_pop23_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_mul534_push23_mul534_pop23_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_mul534_push23_mul534_pop23_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_mul534_push23_mul534_pop23_stall_in = 1'b0;
assign rnode_4to6_bb3_mul534_push23_mul534_pop23_0_NO_SHIFT_REG = rnode_4to6_bb3_mul534_push23_mul534_pop23_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_mul534_push23_mul534_pop23_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_mul534_push23_mul534_pop23_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_stall_in = 1'b0;
assign rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_NO_SHIFT_REG = rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_mul3723_push19_mul3723_pop19_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_mul3723_push19_mul3723_pop19_stall_in = 1'b0;
assign rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_NO_SHIFT_REG = rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_notcmp1126_push20_notcmp1126_pop20_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notcmp1126_push20_notcmp1126_pop20_stall_in = 1'b0;
assign rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_NO_SHIFT_REG = rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_notexitcond1429_push21_notexitcond1429_pop21_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notexitcond1429_push21_notexitcond1429_pop21_stall_in = 1'b0;
assign rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_NO_SHIFT_REG = rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_stall_in = 1'b0;
assign rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_NO_SHIFT_REG = rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_fifo.DATA_WIDTH = 64;
defparam rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_stall_in = 1'b0;
assign rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_NO_SHIFT_REG = rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3__push25__pop25_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push25__pop25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3__push25__pop25_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push25__pop25_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3__push25__pop25_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push25__pop25_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push25__pop25_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push25__pop25_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3__push25__pop25_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3__push25__pop25_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3__push25__pop25_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3__push25__pop25_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3__push25__pop25_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3__push25__pop25_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3__push25__pop25_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3__push25__pop25_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3__push25__pop25_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_4to6_bb3__push25__pop25_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3__push25__pop25_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3__push25__pop25_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__push25__pop25_stall_in = 1'b0;
assign rnode_4to6_bb3__push25__pop25_0_NO_SHIFT_REG = rnode_4to6_bb3__push25__pop25_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3__push25__pop25_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3__push25__pop25_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_stall_in = 1'b0;
assign rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_NO_SHIFT_REG = rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3__push27__pop27_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push27__pop27_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3__push27__pop27_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push27__pop27_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to6_bb3__push27__pop27_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push27__pop27_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push27__pop27_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3__push27__pop27_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3__push27__pop27_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3__push27__pop27_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3__push27__pop27_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3__push27__pop27_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3__push27__pop27_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3__push27__pop27_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3__push27__pop27_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3__push27__pop27_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3__push27__pop27_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_4to6_bb3__push27__pop27_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3__push27__pop27_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3__push27__pop27_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3__push27__pop27_stall_in = 1'b0;
assign rnode_4to6_bb3__push27__pop27_0_NO_SHIFT_REG = rnode_4to6_bb3__push27__pop27_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3__push27__pop27_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3__push27__pop27_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_notcmp40_push28_notcmp40_pop28_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notcmp40_push28_notcmp40_pop28_stall_in = 1'b0;
assign rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_NO_SHIFT_REG = rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb3_notexitcond942_push29_notexitcond942_pop29_NO_SHIFT_REG),
	.data_out(rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_fifo.DEPTH = 2;
defparam rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notexitcond942_push29_notexitcond942_pop29_stall_in = 1'b0;
assign rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_NO_SHIFT_REG = rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_reg_6_NO_SHIFT_REG;
assign rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_notexitcond5_notexit6_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_notexitcond5_notexit6_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_notexitcond5_notexit6_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_notexitcond5_notexit6_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_notexitcond5_notexit6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG = rnode_4to5_bb3_notexitcond5_notexit6_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_notexitcond5_notexit6_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_notexitcond5_notexit6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_i_211_push17_inc34_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_i_211_push17_inc34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_i_211_push17_inc34_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_i_211_push17_inc34_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_i_211_push17_inc34_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_i_211_push17_inc34_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_i_211_push17_inc34_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_i_211_push17_inc34_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_i_211_push17_inc34_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_i_211_push17_inc34_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_i_211_push17_inc34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_i_211_push17_inc34_0_NO_SHIFT_REG = rnode_4to5_bb3_i_211_push17_inc34_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_i_211_push17_inc34_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_i_211_push17_inc34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi3_stall_local;
wire [447:0] local_bb3_c0_exi3;

assign local_bb3_c0_exi3[95:0] = local_bb3_c0_exi2[95:0];
assign local_bb3_c0_exi3[96] = rnode_5to6_bb3_var__0_NO_SHIFT_REG;
assign local_bb3_c0_exi3[447:97] = local_bb3_c0_exi2[447:97];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_notexitcond5_notexit6_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_notexitcond5_notexit6_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_notexitcond5_notexit6_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_notexitcond5_notexit6_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_notexitcond5_notexit6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG = rnode_5to6_bb3_notexitcond5_notexit6_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_notexitcond5_notexit6_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond5_notexit6_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb3_i_211_push17_inc34_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb3_i_211_push17_inc34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_i_211_push17_inc34_0_NO_SHIFT_REG;
 logic rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_i_211_push17_inc34_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_i_211_push17_inc34_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb3_i_211_push17_inc34_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb3_i_211_push17_inc34_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb3_i_211_push17_inc34_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb3_i_211_push17_inc34_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_4to5_bb3_i_211_push17_inc34_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_4to5_bb3_i_211_push17_inc34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_i_211_push17_inc34_0_NO_SHIFT_REG = rnode_5to6_bb3_i_211_push17_inc34_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb3_i_211_push17_inc34_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_i_211_push17_inc34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi4_stall_local;
wire [447:0] local_bb3_c0_exi4;

assign local_bb3_c0_exi4[103:0] = local_bb3_c0_exi3[103:0];
assign local_bb3_c0_exi4[104] = rnode_5to6_bb3_notexitcond5_notexit6_0_NO_SHIFT_REG;
assign local_bb3_c0_exi4[447:105] = local_bb3_c0_exi3[447:105];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi5_stall_local;
wire [447:0] local_bb3_c0_exi5;

assign local_bb3_c0_exi5[127:0] = local_bb3_c0_exi4[127:0];
assign local_bb3_c0_exi5[159:128] = rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_NO_SHIFT_REG;
assign local_bb3_c0_exi5[447:160] = local_bb3_c0_exi4[447:160];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi6_stall_local;
wire [447:0] local_bb3_c0_exi6;

assign local_bb3_c0_exi6[159:0] = local_bb3_c0_exi5[159:0];
assign local_bb3_c0_exi6[191:160] = rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_NO_SHIFT_REG;
assign local_bb3_c0_exi6[447:192] = local_bb3_c0_exi5[447:192];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi7_stall_local;
wire [447:0] local_bb3_c0_exi7;

assign local_bb3_c0_exi7[191:0] = local_bb3_c0_exi6[191:0];
assign local_bb3_c0_exi7[192] = rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_NO_SHIFT_REG;
assign local_bb3_c0_exi7[447:193] = local_bb3_c0_exi6[447:193];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi8_stall_local;
wire [447:0] local_bb3_c0_exi8;

assign local_bb3_c0_exi8[199:0] = local_bb3_c0_exi7[199:0];
assign local_bb3_c0_exi8[200] = rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_NO_SHIFT_REG;
assign local_bb3_c0_exi8[447:201] = local_bb3_c0_exi7[447:201];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi9_stall_local;
wire [447:0] local_bb3_c0_exi9;

assign local_bb3_c0_exi9[207:0] = local_bb3_c0_exi8[207:0];
assign local_bb3_c0_exi9[208] = rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_NO_SHIFT_REG;
assign local_bb3_c0_exi9[447:209] = local_bb3_c0_exi8[447:209];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi10_stall_local;
wire [447:0] local_bb3_c0_exi10;

assign local_bb3_c0_exi10[255:0] = local_bb3_c0_exi9[255:0];
assign local_bb3_c0_exi10[319:256] = rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_NO_SHIFT_REG;
assign local_bb3_c0_exi10[447:320] = local_bb3_c0_exi9[447:320];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi11_stall_local;
wire [447:0] local_bb3_c0_exi11;

assign local_bb3_c0_exi11[319:0] = local_bb3_c0_exi10[319:0];
assign local_bb3_c0_exi11[351:320] = rnode_5to6_bb3__pop25_c0_ene9_0_NO_SHIFT_REG;
assign local_bb3_c0_exi11[447:352] = local_bb3_c0_exi10[447:352];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi12_stall_local;
wire [447:0] local_bb3_c0_exi12;

assign local_bb3_c0_exi12[351:0] = local_bb3_c0_exi11[351:0];
assign local_bb3_c0_exi12[352] = rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_NO_SHIFT_REG;
assign local_bb3_c0_exi12[447:353] = local_bb3_c0_exi11[447:353];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi13_stall_local;
wire [447:0] local_bb3_c0_exi13;

assign local_bb3_c0_exi13[383:0] = local_bb3_c0_exi12[383:0];
assign local_bb3_c0_exi13[415:384] = rnode_5to6_bb3__pop27_c0_ene11_0_NO_SHIFT_REG;
assign local_bb3_c0_exi13[447:416] = local_bb3_c0_exi12[447:416];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi14_stall_local;
wire [447:0] local_bb3_c0_exi14;

assign local_bb3_c0_exi14[415:0] = local_bb3_c0_exi13[415:0];
assign local_bb3_c0_exi14[416] = rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_NO_SHIFT_REG;
assign local_bb3_c0_exi14[447:417] = local_bb3_c0_exi13[447:417];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi15_valid_out;
wire local_bb3_c0_exi15_stall_in;
wire local_bb3_c0_exi15_inputs_ready;
wire local_bb3_c0_exi15_stall_local;
wire [447:0] local_bb3_c0_exi15;

assign local_bb3_c0_exi15_inputs_ready = (rnode_5to6_bb3_mul534_pop23_c0_ene2_0_valid_out_NO_SHIFT_REG & local_bb3_mul24_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_var__0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3__pop25_c0_ene9_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3__pop27_c0_ene11_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb3_notexitcond5_notexit6_0_valid_out_NO_SHIFT_REG);
assign local_bb3_c0_exi15[423:0] = local_bb3_c0_exi14[423:0];
assign local_bb3_c0_exi15[424] = rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_NO_SHIFT_REG;
assign local_bb3_c0_exi15[447:425] = local_bb3_c0_exi14[447:425];
assign local_bb3_c0_exi15_valid_out = 1'b1;
assign rnode_5to6_bb3_mul534_pop23_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb3_mul24_stall_in = 1'b0;
assign rnode_5to6_bb3_var__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_pixel_y_020_pop820_pop18_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_mul3723_pop19_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notcmp1126_pop20_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond1429_pop21_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_memdep_phi1_pop932_pop22_c0_ene7_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_indvars_iv_pop1036_pop24_c0_ene8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3__pop25_c0_ene9_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_memdep_phi1_or38_pop26_c0_ene10_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3__pop27_c0_ene11_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notcmp40_pop28_c0_ene12_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond942_pop29_c0_ene13_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_notexitcond5_notexit6_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb3_c0_exit_c0_exi15_inputs_ready;
 reg local_bb3_c0_exit_c0_exi15_valid_out_0_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_0;
 reg local_bb3_c0_exit_c0_exi15_valid_out_1_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_1;
 reg local_bb3_c0_exit_c0_exi15_valid_out_2_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_2;
 reg local_bb3_c0_exit_c0_exi15_valid_out_3_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_3;
 reg local_bb3_c0_exit_c0_exi15_valid_out_4_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_4;
 reg local_bb3_c0_exit_c0_exi15_valid_out_5_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_5;
 reg local_bb3_c0_exit_c0_exi15_valid_out_6_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_6;
 reg local_bb3_c0_exit_c0_exi15_valid_out_7_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_7;
 reg local_bb3_c0_exit_c0_exi15_valid_out_8_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_8;
 reg local_bb3_c0_exit_c0_exi15_valid_out_9_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_9;
 reg local_bb3_c0_exit_c0_exi15_valid_out_10_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_10;
 reg local_bb3_c0_exit_c0_exi15_valid_out_11_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_11;
 reg local_bb3_c0_exit_c0_exi15_valid_out_12_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_12;
 reg local_bb3_c0_exit_c0_exi15_valid_out_13_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_13;
 reg local_bb3_c0_exit_c0_exi15_valid_out_14_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi15_stall_in_14;
 reg [447:0] local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG;
wire [447:0] local_bb3_c0_exit_c0_exi15_in;
wire local_bb3_c0_exit_c0_exi15_valid;
wire local_bb3_c0_exit_c0_exi15_causedstall;

acl_stall_free_sink local_bb3_c0_exit_c0_exi15_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb3_c0_exi15),
	.data_out(local_bb3_c0_exit_c0_exi15_in),
	.input_accepted(local_bb3_c0_enter_c0_eni13_input_accepted),
	.valid_out(local_bb3_c0_exit_c0_exi15_valid),
	.stall_in(~(local_bb3_c0_exit_c0_exi15_output_regs_ready)),
	.stall_entry(local_bb3_c0_exit_c0_exi15_entry_stall),
	.valid_in(local_bb3_c0_exit_c0_exi15_valid_in),
	.IIphases(local_bb3_c0_exit_c0_exi15_phases),
	.inc_pipelined_thread(local_bb3_c0_enter_c0_eni13_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb3_c0_enter_c0_eni13_dec_pipelined_thread)
);

defparam local_bb3_c0_exit_c0_exi15_instance.DATA_WIDTH = 448;
defparam local_bb3_c0_exit_c0_exi15_instance.PIPELINE_DEPTH = 10;
defparam local_bb3_c0_exit_c0_exi15_instance.SHARINGII = 1;
defparam local_bb3_c0_exit_c0_exi15_instance.SCHEDULEII = 1;
defparam local_bb3_c0_exit_c0_exi15_instance.ALWAYS_THROTTLE = 0;

assign local_bb3_c0_exit_c0_exi15_inputs_ready = 1'b1;
assign local_bb3_c0_exit_c0_exi15_output_regs_ready = ((~(local_bb3_c0_exit_c0_exi15_valid_out_0_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_0)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_1_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_1)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_2_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_2)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_3_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_3)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_4_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_4)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_5_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_5)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_6_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_6)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_7_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_7)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_8_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_8)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_9_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_9)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_10_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_10)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_11_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_11)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_12_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_12)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_13_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_13)) & (~(local_bb3_c0_exit_c0_exi15_valid_out_14_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi15_stall_in_14)));
assign local_bb3_c0_exit_c0_exi15_valid_in = SFC_1_VALID_5_6_0_NO_SHIFT_REG;
assign local_bb3_c0_exi15_stall_in = 1'b0;
assign SFC_1_VALID_5_6_0_stall_in = 1'b0;
assign rnode_4to6_bb3_mul534_push23_mul534_pop23_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_pixel_y_020_pop820_push18_pixel_y_020_pop820_pop18_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_mul3723_push19_mul3723_pop19_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notcmp1126_push20_notcmp1126_pop20_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notexitcond1429_push21_notexitcond1429_pop21_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_memdep_phi1_pop932_push22_memdep_phi1_pop932_pop22_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_indvars_iv_pop1036_push24_indvars_iv_pop1036_pop24_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3__push25__pop25_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_memdep_phi1_or38_push26_memdep_phi1_or38_pop26_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3__push27__pop27_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notcmp40_push28_notcmp40_pop28_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to6_bb3_notexitcond942_push29_notexitcond942_pop29_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_keep_going4_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb3_i_211_push17_inc34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb3_c0_exit_c0_exi15_causedstall = (1'b1 && (1'b0 && !(~(local_bb3_c0_exit_c0_exi15_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG <= 'x;
		local_bb3_c0_exit_c0_exi15_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_7_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_8_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_9_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_10_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_11_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_12_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_13_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi15_valid_out_14_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_c0_exit_c0_exi15_output_regs_ready)
		begin
			local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_in;
			local_bb3_c0_exit_c0_exi15_valid_out_0_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_1_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_2_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_3_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_4_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_5_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_6_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_7_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_8_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_9_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_10_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_11_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_12_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_13_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
			local_bb3_c0_exit_c0_exi15_valid_out_14_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi15_valid;
		end
		else
		begin
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_0))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_1))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_2))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_3))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_4))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_5))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_6))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_7))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_8))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_9))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_9_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_10))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_10_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_11))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_11_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_12))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_12_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_13))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_13_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi15_stall_in_14))
			begin
				local_bb3_c0_exit_c0_exi15_valid_out_14_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe1_stall_local;
wire [31:0] local_bb3_c0_exe1;

assign local_bb3_c0_exe1 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe2_stall_local;
wire [31:0] local_bb3_c0_exe2;

assign local_bb3_c0_exe2 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[95:64];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe3_stall_local;
wire local_bb3_c0_exe3;

assign local_bb3_c0_exe3 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[96];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe4_stall_local;
wire local_bb3_c0_exe4;

assign local_bb3_c0_exe4 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[104];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe5_stall_local;
wire [31:0] local_bb3_c0_exe5;

assign local_bb3_c0_exe5 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[159:128];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe6_stall_local;
wire [31:0] local_bb3_c0_exe6;

assign local_bb3_c0_exe6 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[191:160];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe7_stall_local;
wire local_bb3_c0_exe7;

assign local_bb3_c0_exe7 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[192];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe8_stall_local;
wire local_bb3_c0_exe8;

assign local_bb3_c0_exe8 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[200];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe9_stall_local;
wire local_bb3_c0_exe9;

assign local_bb3_c0_exe9 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[208];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe10_stall_local;
wire [63:0] local_bb3_c0_exe10;

assign local_bb3_c0_exe10 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[319:256];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe11_stall_local;
wire [31:0] local_bb3_c0_exe11;

assign local_bb3_c0_exe11 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[351:320];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe12_stall_local;
wire local_bb3_c0_exe12;

assign local_bb3_c0_exe12 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[352];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe13_stall_local;
wire [31:0] local_bb3_c0_exe13;

assign local_bb3_c0_exe13 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[415:384];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe14_stall_local;
wire local_bb3_c0_exe14;

assign local_bb3_c0_exe14 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[416];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe15_valid_out;
wire local_bb3_c0_exe15_stall_in;
wire local_bb3_c0_exe14_valid_out;
wire local_bb3_c0_exe14_stall_in;
wire local_bb3_c0_exe13_valid_out;
wire local_bb3_c0_exe13_stall_in;
wire local_bb3_c0_exe12_valid_out;
wire local_bb3_c0_exe12_stall_in;
wire local_bb3_c0_exe11_valid_out;
wire local_bb3_c0_exe11_stall_in;
wire local_bb3_c0_exe10_valid_out;
wire local_bb3_c0_exe10_stall_in;
wire local_bb3_c0_exe9_valid_out;
wire local_bb3_c0_exe9_stall_in;
wire local_bb3_c0_exe8_valid_out;
wire local_bb3_c0_exe8_stall_in;
wire local_bb3_c0_exe7_valid_out;
wire local_bb3_c0_exe7_stall_in;
wire local_bb3_c0_exe6_valid_out;
wire local_bb3_c0_exe6_stall_in;
wire local_bb3_c0_exe5_valid_out;
wire local_bb3_c0_exe5_stall_in;
wire local_bb3_c0_exe4_valid_out;
wire local_bb3_c0_exe4_stall_in;
wire local_bb3_c0_exe3_valid_out;
wire local_bb3_c0_exe3_stall_in;
wire local_bb3_c0_exe2_valid_out;
wire local_bb3_c0_exe2_stall_in;
wire local_bb3_c0_exe1_valid_out;
wire local_bb3_c0_exe1_stall_in;
wire local_bb3_c0_exe15_inputs_ready;
wire local_bb3_c0_exe15_stall_local;
wire local_bb3_c0_exe15;

assign local_bb3_c0_exe15_inputs_ready = (local_bb3_c0_exit_c0_exi15_valid_out_14_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_13_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_12_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_11_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_10_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_9_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_8_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_7_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_6_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_5_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_4_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_3_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_2_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_1_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi15_valid_out_0_NO_SHIFT_REG);
assign local_bb3_c0_exe15 = local_bb3_c0_exit_c0_exi15_NO_SHIFT_REG[424];
assign local_bb3_c0_exe15_stall_local = (local_bb3_c0_exe15_stall_in | local_bb3_c0_exe14_stall_in | local_bb3_c0_exe13_stall_in | local_bb3_c0_exe12_stall_in | local_bb3_c0_exe11_stall_in | local_bb3_c0_exe10_stall_in | local_bb3_c0_exe9_stall_in | local_bb3_c0_exe8_stall_in | local_bb3_c0_exe7_stall_in | local_bb3_c0_exe6_stall_in | local_bb3_c0_exe5_stall_in | local_bb3_c0_exe4_stall_in | local_bb3_c0_exe3_stall_in | local_bb3_c0_exe2_stall_in | local_bb3_c0_exe1_stall_in);
assign local_bb3_c0_exe15_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe14_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe13_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe12_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe11_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe10_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe9_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe8_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe7_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe6_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe5_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe4_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe3_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe2_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exe1_valid_out = local_bb3_c0_exe15_inputs_ready;
assign local_bb3_c0_exit_c0_exi15_stall_in_14 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_13 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_12 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_11 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_10 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_9 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_8 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_7 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_6 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_5 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_4 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_3 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_2 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_1 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));
assign local_bb3_c0_exit_c0_exi15_stall_in_0 = (local_bb3_c0_exe15_stall_local | ~(local_bb3_c0_exe15_inputs_ready));

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg lvb_forked16_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe1_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe2_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe3_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe4_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe5_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe6_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe7_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe8_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe9_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb3_c0_exe10_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe11_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe12_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe13_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe14_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe15_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb3_c0_exe15_valid_out & local_bb3_c0_exe14_valid_out & local_bb3_c0_exe13_valid_out & local_bb3_c0_exe12_valid_out & local_bb3_c0_exe11_valid_out & local_bb3_c0_exe10_valid_out & local_bb3_c0_exe9_valid_out & local_bb3_c0_exe8_valid_out & local_bb3_c0_exe7_valid_out & local_bb3_c0_exe6_valid_out & local_bb3_c0_exe5_valid_out & local_bb3_c0_exe4_valid_out & local_bb3_c0_exe3_valid_out & local_bb3_c0_exe2_valid_out & local_bb3_c0_exe1_valid_out & rnode_10to11_forked16_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb3_c0_exe15_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe14_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe13_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe12_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe11_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe10_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe9_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe8_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe7_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe6_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe5_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe4_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe3_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_10to11_forked16_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_forked16 = lvb_forked16_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe1 = lvb_bb3_c0_exe1_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe2 = lvb_bb3_c0_exe2_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe3 = lvb_bb3_c0_exe3_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe4 = lvb_bb3_c0_exe4_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe5 = lvb_bb3_c0_exe5_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe6 = lvb_bb3_c0_exe6_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe7 = lvb_bb3_c0_exe7_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe8 = lvb_bb3_c0_exe8_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe9 = lvb_bb3_c0_exe9_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe10 = lvb_bb3_c0_exe10_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe11 = lvb_bb3_c0_exe11_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe12 = lvb_bb3_c0_exe12_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe13 = lvb_bb3_c0_exe13_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe14 = lvb_bb3_c0_exe14_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe15 = lvb_bb3_c0_exe15_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_forked16_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe1_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe2_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe3_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe4_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe5_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe6_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe7_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe8_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe9_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe10_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe11_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe12_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe13_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe14_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe15_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_forked16_reg_NO_SHIFT_REG <= rnode_10to11_forked16_0_NO_SHIFT_REG;
			lvb_bb3_c0_exe1_reg_NO_SHIFT_REG <= local_bb3_c0_exe1;
			lvb_bb3_c0_exe2_reg_NO_SHIFT_REG <= local_bb3_c0_exe2;
			lvb_bb3_c0_exe3_reg_NO_SHIFT_REG <= local_bb3_c0_exe3;
			lvb_bb3_c0_exe4_reg_NO_SHIFT_REG <= local_bb3_c0_exe4;
			lvb_bb3_c0_exe5_reg_NO_SHIFT_REG <= local_bb3_c0_exe5;
			lvb_bb3_c0_exe6_reg_NO_SHIFT_REG <= local_bb3_c0_exe6;
			lvb_bb3_c0_exe7_reg_NO_SHIFT_REG <= local_bb3_c0_exe7;
			lvb_bb3_c0_exe8_reg_NO_SHIFT_REG <= local_bb3_c0_exe8;
			lvb_bb3_c0_exe9_reg_NO_SHIFT_REG <= local_bb3_c0_exe9;
			lvb_bb3_c0_exe10_reg_NO_SHIFT_REG <= local_bb3_c0_exe10;
			lvb_bb3_c0_exe11_reg_NO_SHIFT_REG <= local_bb3_c0_exe11;
			lvb_bb3_c0_exe12_reg_NO_SHIFT_REG <= local_bb3_c0_exe12;
			lvb_bb3_c0_exe13_reg_NO_SHIFT_REG <= local_bb3_c0_exe13;
			lvb_bb3_c0_exe14_reg_NO_SHIFT_REG <= local_bb3_c0_exe14;
			lvb_bb3_c0_exe15_reg_NO_SHIFT_REG <= local_bb3_c0_exe15;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_4
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_in,
		input [31:0] 		input_r,
		input [31:0] 		input_e_d,
		input [31:0] 		input_wii_div,
		input [31:0] 		input_wii_div1,
		input 		input_wii_cmp19,
		input [31:0] 		input_wii_add7,
		input [31:0] 		input_wii_sub20,
		input [31:0] 		input_wii_sub22,
		input 		input_wii_var_,
		input 		input_wii_var__u17,
		input 		input_wii_var__u18,
		input 		input_wii_var__u19,
		input 		valid_in_0,
		output 		stall_out_0,
		input 		input_forked_0,
		input [31:0] 		input_pixel_y_020_pop821_0,
		input [31:0] 		input_mul3724_0,
		input 		input_notcmp1127_0,
		input 		input_notexitcond1430_0,
		input 		input_memdep_phi1_pop933_0,
		input [31:0] 		input_mul535_0,
		input [63:0] 		input_indvars_iv_pop1037_0,
		input [31:0] 		input_var__u20_0,
		input 		input_memdep_phi1_or39_0,
		input [31:0] 		input_var__u21_0,
		input 		input_notcmp41_0,
		input 		input_notexitcond943_0,
		input 		input_forked1644_0,
		input [31:0] 		input_mul2445_0,
		input 		input_var__u22_0,
		input 		input_notexitcond546_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input 		input_forked_1,
		input [31:0] 		input_pixel_y_020_pop821_1,
		input [31:0] 		input_mul3724_1,
		input 		input_notcmp1127_1,
		input 		input_notexitcond1430_1,
		input 		input_memdep_phi1_pop933_1,
		input [31:0] 		input_mul535_1,
		input [63:0] 		input_indvars_iv_pop1037_1,
		input [31:0] 		input_var__u20_1,
		input 		input_memdep_phi1_or39_1,
		input [31:0] 		input_var__u21_1,
		input 		input_notcmp41_1,
		input 		input_notexitcond943_1,
		input 		input_forked1644_1,
		input [31:0] 		input_mul2445_1,
		input 		input_var__u22_1,
		input 		input_notexitcond546_1,
		output 		valid_out_0,
		input 		stall_in_0,
		output [447:0] 		lvb_bb4_c0_exit87_c0_exi1386_0,
		output [31:0] 		lvb_bb4_c0_exe794_0,
		output 		lvb_bb4_c0_exe895_0,
		output 		lvb_bb4_c0_exe996_0,
		output [63:0] 		lvb_bb4_c0_exe1097_0,
		output 		lvb_bb4_c0_exe1198_0,
		output 		lvb_bb4_c0_exe1299_0,
		output [31:0] 		lvb_bb4_c1_exe1_0,
		output [31:0] 		lvb_bb4_c1_exe2_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [447:0] 		lvb_bb4_c0_exit87_c0_exi1386_1,
		output [31:0] 		lvb_bb4_c0_exe794_1,
		output 		lvb_bb4_c0_exe895_1,
		output 		lvb_bb4_c0_exe996_1,
		output [63:0] 		lvb_bb4_c0_exe1097_1,
		output 		lvb_bb4_c0_exe1198_1,
		output 		lvb_bb4_c0_exe1299_1,
		output [31:0] 		lvb_bb4_c1_exe1_1,
		output [31:0] 		lvb_bb4_c1_exe2_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		feedback_valid_in_30,
		output 		feedback_stall_out_30,
		input [31:0] 		feedback_data_in_30,
		input 		feedback_valid_in_40,
		output 		feedback_stall_out_40,
		input [31:0] 		feedback_data_in_40,
		output 		feedback_stall_out_0,
		input 		feedback_valid_in_1,
		output 		feedback_stall_out_1,
		input 		feedback_data_in_1,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		input 		feedback_valid_in_46,
		output 		feedback_stall_out_46,
		input [31:0] 		feedback_data_in_46,
		input 		feedback_valid_in_45,
		output 		feedback_stall_out_45,
		input 		feedback_data_in_45,
		input 		feedback_valid_in_41,
		output 		feedback_stall_out_41,
		input 		feedback_data_in_41,
		input 		feedback_valid_in_42,
		output 		feedback_stall_out_42,
		input [31:0] 		feedback_data_in_42,
		input 		feedback_valid_in_33,
		output 		feedback_stall_out_33,
		input [31:0] 		feedback_data_in_33,
		input 		feedback_valid_in_34,
		output 		feedback_stall_out_34,
		input [31:0] 		feedback_data_in_34,
		input 		feedback_valid_in_35,
		output 		feedback_stall_out_35,
		input 		feedback_data_in_35,
		input 		feedback_valid_in_36,
		output 		feedback_stall_out_36,
		input 		feedback_data_in_36,
		input 		feedback_valid_in_37,
		output 		feedback_stall_out_37,
		input 		feedback_data_in_37,
		input 		feedback_valid_in_38,
		output 		feedback_stall_out_38,
		input [31:0] 		feedback_data_in_38,
		input 		feedback_valid_in_39,
		output 		feedback_stall_out_39,
		input [63:0] 		feedback_data_in_39,
		input 		feedback_valid_in_43,
		output 		feedback_stall_out_43,
		input 		feedback_data_in_43,
		input 		feedback_valid_in_44,
		output 		feedback_stall_out_44,
		input 		feedback_data_in_44,
		input 		feedback_valid_in_47,
		output 		feedback_stall_out_47,
		input 		feedback_data_in_47,
		output 		feedback_valid_out_1,
		input 		feedback_stall_in_1,
		output 		feedback_data_out_1,
		output 		feedback_valid_out_30,
		input 		feedback_stall_in_30,
		output [31:0] 		feedback_data_out_30,
		output 		feedback_valid_out_45,
		input 		feedback_stall_in_45,
		output 		feedback_data_out_45,
		output 		feedback_valid_out_42,
		input 		feedback_stall_in_42,
		output [31:0] 		feedback_data_out_42,
		output 		feedback_valid_out_41,
		input 		feedback_stall_in_41,
		output 		feedback_data_out_41,
		output 		feedback_valid_out_40,
		input 		feedback_stall_in_40,
		output [31:0] 		feedback_data_out_40,
		output 		feedback_valid_out_33,
		input 		feedback_stall_in_33,
		output [31:0] 		feedback_data_out_33,
		output 		feedback_valid_out_34,
		input 		feedback_stall_in_34,
		output [31:0] 		feedback_data_out_34,
		output 		feedback_valid_out_35,
		input 		feedback_stall_in_35,
		output 		feedback_data_out_35,
		output 		feedback_valid_out_36,
		input 		feedback_stall_in_36,
		output 		feedback_data_out_36,
		output 		feedback_valid_out_37,
		input 		feedback_stall_in_37,
		output 		feedback_data_out_37,
		output 		feedback_valid_out_38,
		input 		feedback_stall_in_38,
		output [31:0] 		feedback_data_out_38,
		output 		feedback_valid_out_39,
		input 		feedback_stall_in_39,
		output [63:0] 		feedback_data_out_39,
		output 		feedback_valid_out_43,
		input 		feedback_stall_in_43,
		output 		feedback_data_out_43,
		output 		feedback_valid_out_44,
		input 		feedback_stall_in_44,
		output 		feedback_data_out_44,
		output 		feedback_valid_out_47,
		input 		feedback_stall_in_47,
		output 		feedback_data_out_47,
		output 		feedback_valid_out_46,
		input 		feedback_stall_in_46,
		output [31:0] 		feedback_data_out_46,
		input [511:0] 		avm_local_bb4_ld__readdata,
		input 		avm_local_bb4_ld__readdatavalid,
		input 		avm_local_bb4_ld__waitrequest,
		output [32:0] 		avm_local_bb4_ld__address,
		output 		avm_local_bb4_ld__read,
		output 		avm_local_bb4_ld__write,
		input 		avm_local_bb4_ld__writeack,
		output [511:0] 		avm_local_bb4_ld__writedata,
		output [63:0] 		avm_local_bb4_ld__byteenable,
		output [4:0] 		avm_local_bb4_ld__burstcount,
		output 		local_bb4_ld__active,
		input 		clock2x,
		input 		feedback_valid_in_48,
		output 		feedback_stall_out_48,
		input 		feedback_data_in_48,
		output 		feedback_valid_out_48,
		input 		feedback_stall_in_48,
		output 		feedback_data_out_48,
		input 		feedback_valid_in_31,
		output 		feedback_stall_out_31,
		input [31:0] 		feedback_data_in_31,
		input 		feedback_valid_in_32,
		output 		feedback_stall_out_32,
		input [31:0] 		feedback_data_in_32,
		output 		feedback_valid_out_32,
		input 		feedback_stall_in_32,
		output [31:0] 		feedback_data_out_32,
		output 		feedback_valid_out_31,
		input 		feedback_stall_in_31,
		output [31:0] 		feedback_data_out_31
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_node_stall_in_8;
 reg merge_node_valid_out_8_NO_SHIFT_REG;
wire merge_node_stall_in_9;
 reg merge_node_valid_out_9_NO_SHIFT_REG;
wire merge_node_stall_in_10;
 reg merge_node_valid_out_10_NO_SHIFT_REG;
wire merge_node_stall_in_11;
 reg merge_node_valid_out_11_NO_SHIFT_REG;
wire merge_node_stall_in_12;
 reg merge_node_valid_out_12_NO_SHIFT_REG;
wire merge_node_stall_in_13;
 reg merge_node_valid_out_13_NO_SHIFT_REG;
wire merge_node_stall_in_14;
 reg merge_node_valid_out_14_NO_SHIFT_REG;
wire merge_node_stall_in_15;
 reg merge_node_valid_out_15_NO_SHIFT_REG;
wire merge_node_stall_in_16;
 reg merge_node_valid_out_16_NO_SHIFT_REG;
wire merge_node_stall_in_17;
 reg merge_node_valid_out_17_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg input_forked_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pixel_y_020_pop821_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul3724_0_staging_reg_NO_SHIFT_REG;
 reg input_notcmp1127_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1430_0_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_pop933_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul535_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_pop1037_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u20_0_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_or39_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u21_0_staging_reg_NO_SHIFT_REG;
 reg input_notcmp41_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond943_0_staging_reg_NO_SHIFT_REG;
 reg input_forked1644_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul2445_0_staging_reg_NO_SHIFT_REG;
 reg input_var__u22_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond546_0_staging_reg_NO_SHIFT_REG;
 reg local_lvm_forked_NO_SHIFT_REG;
 reg [31:0] local_lvm_pixel_y_020_pop821_NO_SHIFT_REG;
 reg [31:0] local_lvm_mul3724_NO_SHIFT_REG;
 reg local_lvm_notcmp1127_NO_SHIFT_REG;
 reg local_lvm_notexitcond1430_NO_SHIFT_REG;
 reg local_lvm_memdep_phi1_pop933_NO_SHIFT_REG;
 reg [31:0] local_lvm_mul535_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv_pop1037_NO_SHIFT_REG;
 reg [31:0] local_lvm_var__u20_NO_SHIFT_REG;
 reg local_lvm_memdep_phi1_or39_NO_SHIFT_REG;
 reg [31:0] local_lvm_var__u21_NO_SHIFT_REG;
 reg local_lvm_notcmp41_NO_SHIFT_REG;
 reg local_lvm_notexitcond943_NO_SHIFT_REG;
 reg local_lvm_forked1644_NO_SHIFT_REG;
 reg [31:0] local_lvm_mul2445_NO_SHIFT_REG;
 reg local_lvm_var__u22_NO_SHIFT_REG;
 reg local_lvm_notexitcond546_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg input_forked_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pixel_y_020_pop821_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul3724_1_staging_reg_NO_SHIFT_REG;
 reg input_notcmp1127_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1430_1_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_pop933_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul535_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_pop1037_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u20_1_staging_reg_NO_SHIFT_REG;
 reg input_memdep_phi1_or39_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_var__u21_1_staging_reg_NO_SHIFT_REG;
 reg input_notcmp41_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond943_1_staging_reg_NO_SHIFT_REG;
 reg input_forked1644_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_mul2445_1_staging_reg_NO_SHIFT_REG;
 reg input_var__u22_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond546_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG) | (merge_node_stall_in_8 & merge_node_valid_out_8_NO_SHIFT_REG) | (merge_node_stall_in_9 & merge_node_valid_out_9_NO_SHIFT_REG) | (merge_node_stall_in_10 & merge_node_valid_out_10_NO_SHIFT_REG) | (merge_node_stall_in_11 & merge_node_valid_out_11_NO_SHIFT_REG) | (merge_node_stall_in_12 & merge_node_valid_out_12_NO_SHIFT_REG) | (merge_node_stall_in_13 & merge_node_valid_out_13_NO_SHIFT_REG) | (merge_node_stall_in_14 & merge_node_valid_out_14_NO_SHIFT_REG) | (merge_node_stall_in_15 & merge_node_valid_out_15_NO_SHIFT_REG) | (merge_node_stall_in_16 & merge_node_valid_out_16_NO_SHIFT_REG) | (merge_node_stall_in_17 & merge_node_valid_out_17_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_forked_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_pixel_y_020_pop821_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul3724_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp1127_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1430_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_pop933_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul535_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_pop1037_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u20_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_or39_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u21_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp41_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond943_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_forked1644_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul2445_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u22_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond546_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_forked_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_pixel_y_020_pop821_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul3724_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp1127_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1430_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_pop933_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul535_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_pop1037_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u20_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_memdep_phi1_or39_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u21_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notcmp41_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond943_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_forked1644_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_mul2445_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u22_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond546_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_forked_0_staging_reg_NO_SHIFT_REG <= input_forked_0;
				input_pixel_y_020_pop821_0_staging_reg_NO_SHIFT_REG <= input_pixel_y_020_pop821_0;
				input_mul3724_0_staging_reg_NO_SHIFT_REG <= input_mul3724_0;
				input_notcmp1127_0_staging_reg_NO_SHIFT_REG <= input_notcmp1127_0;
				input_notexitcond1430_0_staging_reg_NO_SHIFT_REG <= input_notexitcond1430_0;
				input_memdep_phi1_pop933_0_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_pop933_0;
				input_mul535_0_staging_reg_NO_SHIFT_REG <= input_mul535_0;
				input_indvars_iv_pop1037_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv_pop1037_0;
				input_var__u20_0_staging_reg_NO_SHIFT_REG <= input_var__u20_0;
				input_memdep_phi1_or39_0_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_or39_0;
				input_var__u21_0_staging_reg_NO_SHIFT_REG <= input_var__u21_0;
				input_notcmp41_0_staging_reg_NO_SHIFT_REG <= input_notcmp41_0;
				input_notexitcond943_0_staging_reg_NO_SHIFT_REG <= input_notexitcond943_0;
				input_forked1644_0_staging_reg_NO_SHIFT_REG <= input_forked1644_0;
				input_mul2445_0_staging_reg_NO_SHIFT_REG <= input_mul2445_0;
				input_var__u22_0_staging_reg_NO_SHIFT_REG <= input_var__u22_0;
				input_notexitcond546_0_staging_reg_NO_SHIFT_REG <= input_notexitcond546_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_forked_1_staging_reg_NO_SHIFT_REG <= input_forked_1;
				input_pixel_y_020_pop821_1_staging_reg_NO_SHIFT_REG <= input_pixel_y_020_pop821_1;
				input_mul3724_1_staging_reg_NO_SHIFT_REG <= input_mul3724_1;
				input_notcmp1127_1_staging_reg_NO_SHIFT_REG <= input_notcmp1127_1;
				input_notexitcond1430_1_staging_reg_NO_SHIFT_REG <= input_notexitcond1430_1;
				input_memdep_phi1_pop933_1_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_pop933_1;
				input_mul535_1_staging_reg_NO_SHIFT_REG <= input_mul535_1;
				input_indvars_iv_pop1037_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv_pop1037_1;
				input_var__u20_1_staging_reg_NO_SHIFT_REG <= input_var__u20_1;
				input_memdep_phi1_or39_1_staging_reg_NO_SHIFT_REG <= input_memdep_phi1_or39_1;
				input_var__u21_1_staging_reg_NO_SHIFT_REG <= input_var__u21_1;
				input_notcmp41_1_staging_reg_NO_SHIFT_REG <= input_notcmp41_1;
				input_notexitcond943_1_staging_reg_NO_SHIFT_REG <= input_notexitcond943_1;
				input_forked1644_1_staging_reg_NO_SHIFT_REG <= input_forked1644_1;
				input_mul2445_1_staging_reg_NO_SHIFT_REG <= input_mul2445_1;
				input_var__u22_1_staging_reg_NO_SHIFT_REG <= input_var__u22_1;
				input_notexitcond546_1_staging_reg_NO_SHIFT_REG <= input_notexitcond546_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_0_staging_reg_NO_SHIFT_REG;
					local_lvm_pixel_y_020_pop821_NO_SHIFT_REG <= input_pixel_y_020_pop821_0_staging_reg_NO_SHIFT_REG;
					local_lvm_mul3724_NO_SHIFT_REG <= input_mul3724_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp1127_NO_SHIFT_REG <= input_notcmp1127_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1430_NO_SHIFT_REG <= input_notexitcond1430_0_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_pop933_NO_SHIFT_REG <= input_memdep_phi1_pop933_0_staging_reg_NO_SHIFT_REG;
					local_lvm_mul535_NO_SHIFT_REG <= input_mul535_0_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_pop1037_NO_SHIFT_REG <= input_indvars_iv_pop1037_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_0_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_or39_NO_SHIFT_REG <= input_memdep_phi1_or39_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u21_NO_SHIFT_REG <= input_var__u21_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp41_NO_SHIFT_REG <= input_notcmp41_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond943_NO_SHIFT_REG <= input_notexitcond943_0_staging_reg_NO_SHIFT_REG;
					local_lvm_forked1644_NO_SHIFT_REG <= input_forked1644_0_staging_reg_NO_SHIFT_REG;
					local_lvm_mul2445_NO_SHIFT_REG <= input_mul2445_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u22_NO_SHIFT_REG <= input_var__u22_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond546_NO_SHIFT_REG <= input_notexitcond546_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_0;
					local_lvm_pixel_y_020_pop821_NO_SHIFT_REG <= input_pixel_y_020_pop821_0;
					local_lvm_mul3724_NO_SHIFT_REG <= input_mul3724_0;
					local_lvm_notcmp1127_NO_SHIFT_REG <= input_notcmp1127_0;
					local_lvm_notexitcond1430_NO_SHIFT_REG <= input_notexitcond1430_0;
					local_lvm_memdep_phi1_pop933_NO_SHIFT_REG <= input_memdep_phi1_pop933_0;
					local_lvm_mul535_NO_SHIFT_REG <= input_mul535_0;
					local_lvm_indvars_iv_pop1037_NO_SHIFT_REG <= input_indvars_iv_pop1037_0;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_0;
					local_lvm_memdep_phi1_or39_NO_SHIFT_REG <= input_memdep_phi1_or39_0;
					local_lvm_var__u21_NO_SHIFT_REG <= input_var__u21_0;
					local_lvm_notcmp41_NO_SHIFT_REG <= input_notcmp41_0;
					local_lvm_notexitcond943_NO_SHIFT_REG <= input_notexitcond943_0;
					local_lvm_forked1644_NO_SHIFT_REG <= input_forked1644_0;
					local_lvm_mul2445_NO_SHIFT_REG <= input_mul2445_0;
					local_lvm_var__u22_NO_SHIFT_REG <= input_var__u22_0;
					local_lvm_notexitcond546_NO_SHIFT_REG <= input_notexitcond546_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_1_staging_reg_NO_SHIFT_REG;
					local_lvm_pixel_y_020_pop821_NO_SHIFT_REG <= input_pixel_y_020_pop821_1_staging_reg_NO_SHIFT_REG;
					local_lvm_mul3724_NO_SHIFT_REG <= input_mul3724_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp1127_NO_SHIFT_REG <= input_notcmp1127_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1430_NO_SHIFT_REG <= input_notexitcond1430_1_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_pop933_NO_SHIFT_REG <= input_memdep_phi1_pop933_1_staging_reg_NO_SHIFT_REG;
					local_lvm_mul535_NO_SHIFT_REG <= input_mul535_1_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_pop1037_NO_SHIFT_REG <= input_indvars_iv_pop1037_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_1_staging_reg_NO_SHIFT_REG;
					local_lvm_memdep_phi1_or39_NO_SHIFT_REG <= input_memdep_phi1_or39_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u21_NO_SHIFT_REG <= input_var__u21_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notcmp41_NO_SHIFT_REG <= input_notcmp41_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond943_NO_SHIFT_REG <= input_notexitcond943_1_staging_reg_NO_SHIFT_REG;
					local_lvm_forked1644_NO_SHIFT_REG <= input_forked1644_1_staging_reg_NO_SHIFT_REG;
					local_lvm_mul2445_NO_SHIFT_REG <= input_mul2445_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u22_NO_SHIFT_REG <= input_var__u22_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond546_NO_SHIFT_REG <= input_notexitcond546_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_1;
					local_lvm_pixel_y_020_pop821_NO_SHIFT_REG <= input_pixel_y_020_pop821_1;
					local_lvm_mul3724_NO_SHIFT_REG <= input_mul3724_1;
					local_lvm_notcmp1127_NO_SHIFT_REG <= input_notcmp1127_1;
					local_lvm_notexitcond1430_NO_SHIFT_REG <= input_notexitcond1430_1;
					local_lvm_memdep_phi1_pop933_NO_SHIFT_REG <= input_memdep_phi1_pop933_1;
					local_lvm_mul535_NO_SHIFT_REG <= input_mul535_1;
					local_lvm_indvars_iv_pop1037_NO_SHIFT_REG <= input_indvars_iv_pop1037_1;
					local_lvm_var__u20_NO_SHIFT_REG <= input_var__u20_1;
					local_lvm_memdep_phi1_or39_NO_SHIFT_REG <= input_memdep_phi1_or39_1;
					local_lvm_var__u21_NO_SHIFT_REG <= input_var__u21_1;
					local_lvm_notcmp41_NO_SHIFT_REG <= input_notcmp41_1;
					local_lvm_notexitcond943_NO_SHIFT_REG <= input_notexitcond943_1;
					local_lvm_forked1644_NO_SHIFT_REG <= input_forked1644_1;
					local_lvm_mul2445_NO_SHIFT_REG <= input_mul2445_1;
					local_lvm_var__u22_NO_SHIFT_REG <= input_var__u22_1;
					local_lvm_notexitcond546_NO_SHIFT_REG <= input_notexitcond546_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_9_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_10_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_11_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_12_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_13_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_14_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_15_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_16_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_17_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_8_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_9_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_10_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_11_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_12_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_13_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_14_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_15_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_16_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_17_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_8))
			begin
				merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_9))
			begin
				merge_node_valid_out_9_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_10))
			begin
				merge_node_valid_out_10_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_11))
			begin
				merge_node_valid_out_11_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_12))
			begin
				merge_node_valid_out_12_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_13))
			begin
				merge_node_valid_out_13_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_14))
			begin
				merge_node_valid_out_14_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_15))
			begin
				merge_node_valid_out_15_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_16))
			begin
				merge_node_valid_out_16_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_17))
			begin
				merge_node_valid_out_17_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni147_stall_local;
wire [447:0] local_bb4_c0_eni147;

assign local_bb4_c0_eni147[7:0] = 8'bx;
assign local_bb4_c0_eni147[8] = local_lvm_forked1644_NO_SHIFT_REG;
assign local_bb4_c0_eni147[447:9] = 439'bx;

// Register node:
//  * latency = 14
//  * capacity = 14
 logic rnode_1to15_var__u17_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to15_var__u17_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to15_var__u17_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to15_var__u17_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_1to15_var__u17_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_1to15_var__u17_0_stall_out_reg_15_NO_SHIFT_REG;
wire [1:0] rci_rcnode_1to175_rc17_forked_0_reg_1;

acl_data_fifo rnode_1to15_var__u17_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to15_var__u17_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to15_var__u17_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_1to15_var__u17_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_1to15_var__u17_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to15_var__u17_0_reg_15_fifo.DEPTH = 15;
defparam rnode_1to15_var__u17_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_1to15_var__u17_0_reg_15_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to15_var__u17_0_reg_15_fifo.IMPL = "ram";

assign rnode_1to15_var__u17_0_reg_15_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_16_NO_SHIFT_REG;
assign merge_node_stall_in_16 = rnode_1to15_var__u17_0_stall_out_reg_15_NO_SHIFT_REG;
assign rnode_1to15_var__u17_0_stall_in_reg_15_NO_SHIFT_REG = rnode_1to15_var__u17_0_stall_in_NO_SHIFT_REG;
assign rnode_1to15_var__u17_0_valid_out_NO_SHIFT_REG = rnode_1to15_var__u17_0_valid_out_reg_15_NO_SHIFT_REG;
assign rci_rcnode_1to175_rc17_forked_0_reg_1[0] = local_lvm_forked_NO_SHIFT_REG;
assign rci_rcnode_1to175_rc17_forked_0_reg_1[1] = local_lvm_notexitcond546_NO_SHIFT_REG;

// Register node:
//  * latency = 174
//  * capacity = 174
 logic rcnode_1to175_rc17_forked_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to175_rc17_forked_0_stall_in_NO_SHIFT_REG;
 logic [1:0] rcnode_1to175_rc17_forked_0_NO_SHIFT_REG;
 logic rcnode_1to175_rc17_forked_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [1:0] rcnode_1to175_rc17_forked_0_reg_175_NO_SHIFT_REG;
 logic rcnode_1to175_rc17_forked_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rcnode_1to175_rc17_forked_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rcnode_1to175_rc17_forked_0_stall_out_reg_175_IP_NO_SHIFT_REG;
 logic rcnode_1to175_rc17_forked_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rcnode_1to175_rc17_forked_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to175_rc17_forked_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to175_rc17_forked_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rcnode_1to175_rc17_forked_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rcnode_1to175_rc17_forked_0_stall_out_reg_175_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to175_rc17_forked_0_reg_1),
	.data_out(rcnode_1to175_rc17_forked_0_reg_175_NO_SHIFT_REG)
);

defparam rcnode_1to175_rc17_forked_0_reg_175_fifo.DEPTH = 175;
defparam rcnode_1to175_rc17_forked_0_reg_175_fifo.DATA_WIDTH = 2;
defparam rcnode_1to175_rc17_forked_0_reg_175_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to175_rc17_forked_0_reg_175_fifo.IMPL = "ram";

assign rcnode_1to175_rc17_forked_0_reg_175_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_17_NO_SHIFT_REG;
assign rcnode_1to175_rc17_forked_0_stall_out_reg_175_NO_SHIFT_REG = (~(rcnode_1to175_rc17_forked_0_reg_175_inputs_ready_NO_SHIFT_REG) | rcnode_1to175_rc17_forked_0_stall_out_reg_175_IP_NO_SHIFT_REG);
assign merge_node_stall_in_17 = rcnode_1to175_rc17_forked_0_stall_out_reg_175_NO_SHIFT_REG;
assign rcnode_1to175_rc17_forked_0_NO_SHIFT_REG = rcnode_1to175_rc17_forked_0_reg_175_NO_SHIFT_REG;
assign rcnode_1to175_rc17_forked_0_stall_in_reg_175_NO_SHIFT_REG = rcnode_1to175_rc17_forked_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to175_rc17_forked_0_valid_out_NO_SHIFT_REG = rcnode_1to175_rc17_forked_0_valid_out_reg_175_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni248_stall_local;
wire [447:0] local_bb4_c0_eni248;

assign local_bb4_c0_eni248[15:0] = local_bb4_c0_eni147[15:0];
assign local_bb4_c0_eni248[16] = local_lvm_forked_NO_SHIFT_REG;
assign local_bb4_c0_eni248[447:17] = local_bb4_c0_eni147[447:17];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_var__u17_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_var__u17_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_var__u17_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_var__u17_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_var__u17_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_var__u17_0_stall_out_reg_16_NO_SHIFT_REG;
wire [1:0] rci_rcnode_175to176_rc0_forked_0_reg_175;

acl_data_fifo rnode_15to16_var__u17_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_var__u17_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_var__u17_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_var__u17_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_var__u17_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_var__u17_0_reg_16_fifo.DEPTH = 2;
defparam rnode_15to16_var__u17_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_var__u17_0_reg_16_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_15to16_var__u17_0_reg_16_fifo.IMPL = "ll_reg";

assign rnode_15to16_var__u17_0_reg_16_inputs_ready_NO_SHIFT_REG = rnode_1to15_var__u17_0_valid_out_NO_SHIFT_REG;
assign rnode_1to15_var__u17_0_stall_in_NO_SHIFT_REG = rnode_15to16_var__u17_0_stall_out_reg_16_NO_SHIFT_REG;
assign rnode_15to16_var__u17_0_stall_in_reg_16_NO_SHIFT_REG = rnode_15to16_var__u17_0_stall_in_NO_SHIFT_REG;
assign rnode_15to16_var__u17_0_valid_out_NO_SHIFT_REG = rnode_15to16_var__u17_0_valid_out_reg_16_NO_SHIFT_REG;
assign rci_rcnode_175to176_rc0_forked_0_reg_175[0] = rcnode_1to175_rc17_forked_0_NO_SHIFT_REG[0];
assign rci_rcnode_175to176_rc0_forked_0_reg_175[1] = rcnode_1to175_rc17_forked_0_NO_SHIFT_REG[1];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_175to176_rc0_forked_0_valid_out_0_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_stall_in_0_NO_SHIFT_REG;
 logic [1:0] rcnode_175to176_rc0_forked_0_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_valid_out_1_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_stall_in_1_NO_SHIFT_REG;
 logic [1:0] rcnode_175to176_rc0_forked_1_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_valid_out_2_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_stall_in_2_NO_SHIFT_REG;
 logic [1:0] rcnode_175to176_rc0_forked_2_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [1:0] rcnode_175to176_rc0_forked_0_reg_176_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_stall_out_reg_176_IP_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_forked_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rcnode_175to176_rc0_forked_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_175to176_rc0_forked_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_175to176_rc0_forked_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rcnode_175to176_rc0_forked_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rcnode_175to176_rc0_forked_0_stall_out_reg_176_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_175to176_rc0_forked_0_reg_175),
	.data_out(rcnode_175to176_rc0_forked_0_reg_176_NO_SHIFT_REG)
);

defparam rcnode_175to176_rc0_forked_0_reg_176_fifo.DEPTH = 1;
defparam rcnode_175to176_rc0_forked_0_reg_176_fifo.DATA_WIDTH = 2;
defparam rcnode_175to176_rc0_forked_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_175to176_rc0_forked_0_reg_176_fifo.IMPL = "ll_reg";

assign rcnode_175to176_rc0_forked_0_reg_176_inputs_ready_NO_SHIFT_REG = rcnode_1to175_rc17_forked_0_valid_out_NO_SHIFT_REG;
assign rcnode_175to176_rc0_forked_0_stall_out_reg_176_NO_SHIFT_REG = (~(rcnode_175to176_rc0_forked_0_reg_176_inputs_ready_NO_SHIFT_REG) | rcnode_175to176_rc0_forked_0_stall_out_reg_176_IP_NO_SHIFT_REG);
assign rcnode_1to175_rc17_forked_0_stall_in_NO_SHIFT_REG = rcnode_175to176_rc0_forked_0_stall_out_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_forked_0_stall_in_0_reg_176_NO_SHIFT_REG = (rcnode_175to176_rc0_forked_0_stall_in_0_NO_SHIFT_REG | rcnode_175to176_rc0_forked_0_stall_in_1_NO_SHIFT_REG | rcnode_175to176_rc0_forked_0_stall_in_2_NO_SHIFT_REG);
assign rcnode_175to176_rc0_forked_0_valid_out_0_NO_SHIFT_REG = rcnode_175to176_rc0_forked_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_forked_0_valid_out_1_NO_SHIFT_REG = rcnode_175to176_rc0_forked_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_forked_0_valid_out_2_NO_SHIFT_REG = rcnode_175to176_rc0_forked_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_forked_0_NO_SHIFT_REG = rcnode_175to176_rc0_forked_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_forked_1_NO_SHIFT_REG = rcnode_175to176_rc0_forked_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_forked_2_NO_SHIFT_REG = rcnode_175to176_rc0_forked_0_reg_176_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni349_stall_local;
wire [447:0] local_bb4_c0_eni349;

assign local_bb4_c0_eni349[31:0] = local_bb4_c0_eni248[31:0];
assign local_bb4_c0_eni349[63:32] = local_lvm_var__u20_NO_SHIFT_REG;
assign local_bb4_c0_eni349[447:64] = local_bb4_c0_eni248[447:64];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni1_stall_local;
wire [127:0] local_bb4_c1_eni1;

assign local_bb4_c1_eni1[7:0] = 8'bx;
assign local_bb4_c1_eni1[8] = rcnode_175to176_rc0_forked_0_NO_SHIFT_REG[0];
assign local_bb4_c1_eni1[127:9] = 119'bx;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni450_stall_local;
wire [447:0] local_bb4_c0_eni450;

assign local_bb4_c0_eni450[63:0] = local_bb4_c0_eni349[63:0];
assign local_bb4_c0_eni450[95:64] = local_lvm_mul2445_NO_SHIFT_REG;
assign local_bb4_c0_eni450[447:96] = local_bb4_c0_eni349[447:96];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni551_stall_local;
wire [447:0] local_bb4_c0_eni551;

assign local_bb4_c0_eni551[95:0] = local_bb4_c0_eni450[95:0];
assign local_bb4_c0_eni551[96] = local_lvm_memdep_phi1_or39_NO_SHIFT_REG;
assign local_bb4_c0_eni551[447:97] = local_bb4_c0_eni450[447:97];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni652_stall_local;
wire [447:0] local_bb4_c0_eni652;

assign local_bb4_c0_eni652[127:0] = local_bb4_c0_eni551[127:0];
assign local_bb4_c0_eni652[159:128] = local_lvm_var__u21_NO_SHIFT_REG;
assign local_bb4_c0_eni652[447:160] = local_bb4_c0_eni551[447:160];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni753_stall_local;
wire [447:0] local_bb4_c0_eni753;

assign local_bb4_c0_eni753[159:0] = local_bb4_c0_eni652[159:0];
assign local_bb4_c0_eni753[191:160] = local_lvm_pixel_y_020_pop821_NO_SHIFT_REG;
assign local_bb4_c0_eni753[447:192] = local_bb4_c0_eni652[447:192];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni854_stall_local;
wire [447:0] local_bb4_c0_eni854;

assign local_bb4_c0_eni854[191:0] = local_bb4_c0_eni753[191:0];
assign local_bb4_c0_eni854[223:192] = local_lvm_mul3724_NO_SHIFT_REG;
assign local_bb4_c0_eni854[447:224] = local_bb4_c0_eni753[447:224];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni955_stall_local;
wire [447:0] local_bb4_c0_eni955;

assign local_bb4_c0_eni955[223:0] = local_bb4_c0_eni854[223:0];
assign local_bb4_c0_eni955[224] = local_lvm_notcmp1127_NO_SHIFT_REG;
assign local_bb4_c0_eni955[447:225] = local_bb4_c0_eni854[447:225];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni1056_stall_local;
wire [447:0] local_bb4_c0_eni1056;

assign local_bb4_c0_eni1056[231:0] = local_bb4_c0_eni955[231:0];
assign local_bb4_c0_eni1056[232] = local_lvm_notexitcond1430_NO_SHIFT_REG;
assign local_bb4_c0_eni1056[447:233] = local_bb4_c0_eni955[447:233];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni1157_stall_local;
wire [447:0] local_bb4_c0_eni1157;

assign local_bb4_c0_eni1157[239:0] = local_bb4_c0_eni1056[239:0];
assign local_bb4_c0_eni1157[240] = local_lvm_memdep_phi1_pop933_NO_SHIFT_REG;
assign local_bb4_c0_eni1157[447:241] = local_bb4_c0_eni1056[447:241];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni1258_stall_local;
wire [447:0] local_bb4_c0_eni1258;

assign local_bb4_c0_eni1258[255:0] = local_bb4_c0_eni1157[255:0];
assign local_bb4_c0_eni1258[287:256] = local_lvm_mul535_NO_SHIFT_REG;
assign local_bb4_c0_eni1258[447:288] = local_bb4_c0_eni1157[447:288];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni1359_stall_local;
wire [447:0] local_bb4_c0_eni1359;

assign local_bb4_c0_eni1359[319:0] = local_bb4_c0_eni1258[319:0];
assign local_bb4_c0_eni1359[383:320] = local_lvm_indvars_iv_pop1037_NO_SHIFT_REG;
assign local_bb4_c0_eni1359[447:384] = local_bb4_c0_eni1258[447:384];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni14_stall_local;
wire [447:0] local_bb4_c0_eni14;

assign local_bb4_c0_eni14[383:0] = local_bb4_c0_eni1359[383:0];
assign local_bb4_c0_eni14[384] = local_lvm_notcmp41_NO_SHIFT_REG;
assign local_bb4_c0_eni14[447:385] = local_bb4_c0_eni1359[447:385];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni15_stall_local;
wire [447:0] local_bb4_c0_eni15;

assign local_bb4_c0_eni15[391:0] = local_bb4_c0_eni14[391:0];
assign local_bb4_c0_eni15[392] = local_lvm_notexitcond943_NO_SHIFT_REG;
assign local_bb4_c0_eni15[447:393] = local_bb4_c0_eni14[447:393];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni16_stall_local;
wire [447:0] local_bb4_c0_eni16;

assign local_bb4_c0_eni16[399:0] = local_bb4_c0_eni15[399:0];
assign local_bb4_c0_eni16[400] = local_lvm_var__u22_NO_SHIFT_REG;
assign local_bb4_c0_eni16[447:401] = local_bb4_c0_eni15[447:401];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene161_valid_out;
wire local_bb4_c0_ene161_stall_in;
wire local_bb4_c0_ene262_valid_out;
wire local_bb4_c0_ene262_stall_in;
wire local_bb4_c0_ene363_valid_out;
wire local_bb4_c0_ene363_stall_in;
wire local_bb4_c0_ene464_valid_out;
wire local_bb4_c0_ene464_stall_in;
wire local_bb4_c0_ene565_valid_out;
wire local_bb4_c0_ene565_stall_in;
wire local_bb4_c0_ene666_valid_out;
wire local_bb4_c0_ene666_stall_in;
wire local_bb4_c0_ene767_valid_out;
wire local_bb4_c0_ene767_stall_in;
wire local_bb4_c0_ene868_valid_out;
wire local_bb4_c0_ene868_stall_in;
wire local_bb4_c0_ene969_valid_out;
wire local_bb4_c0_ene969_stall_in;
wire local_bb4_c0_ene1070_valid_out;
wire local_bb4_c0_ene1070_stall_in;
wire local_bb4_c0_ene1171_valid_out;
wire local_bb4_c0_ene1171_stall_in;
wire local_bb4_c0_ene1272_valid_out;
wire local_bb4_c0_ene1272_stall_in;
wire local_bb4_c0_ene1373_valid_out;
wire local_bb4_c0_ene1373_stall_in;
wire local_bb4_c0_ene14_valid_out;
wire local_bb4_c0_ene14_stall_in;
wire local_bb4_c0_ene15_valid_out;
wire local_bb4_c0_ene15_stall_in;
wire local_bb4_c0_ene16_valid_out;
wire local_bb4_c0_ene16_stall_in;
wire SFC_2_VALID_1_1_0_valid_out;
wire SFC_2_VALID_1_1_0_stall_in;
wire local_bb4_c0_enter60_c0_eni16_inputs_ready;
wire local_bb4_c0_enter60_c0_eni16_stall_local;
wire local_bb4_c0_enter60_c0_eni16_input_accepted;
wire [447:0] local_bb4_c0_enter60_c0_eni16;
wire local_bb4_c0_exit87_c0_exi1386_entry_stall;
wire local_bb4_c0_enter60_c0_eni16_valid_bit;
wire local_bb4_c0_exit87_c0_exi1386_output_regs_ready;
wire local_bb4_c0_exit87_c0_exi1386_valid_in;
wire local_bb4_c0_exit87_c0_exi1386_phases;
wire local_bb4_c0_enter60_c0_eni16_inc_pipelined_thread;
wire local_bb4_c0_enter60_c0_eni16_dec_pipelined_thread;
wire local_bb4_c0_enter60_c0_eni16_fu_stall_out;

assign local_bb4_c0_enter60_c0_eni16_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_3_NO_SHIFT_REG & merge_node_valid_out_4_NO_SHIFT_REG & merge_node_valid_out_5_NO_SHIFT_REG & merge_node_valid_out_6_NO_SHIFT_REG & merge_node_valid_out_7_NO_SHIFT_REG & merge_node_valid_out_8_NO_SHIFT_REG & merge_node_valid_out_9_NO_SHIFT_REG & merge_node_valid_out_10_NO_SHIFT_REG & merge_node_valid_out_11_NO_SHIFT_REG & merge_node_valid_out_12_NO_SHIFT_REG & merge_node_valid_out_13_NO_SHIFT_REG & merge_node_valid_out_14_NO_SHIFT_REG & merge_node_valid_out_15_NO_SHIFT_REG);
assign local_bb4_c0_enter60_c0_eni16 = local_bb4_c0_eni16;
assign local_bb4_c0_enter60_c0_eni16_input_accepted = (local_bb4_c0_enter60_c0_eni16_inputs_ready && !(local_bb4_c0_exit87_c0_exi1386_entry_stall));
assign local_bb4_c0_enter60_c0_eni16_valid_bit = local_bb4_c0_enter60_c0_eni16_input_accepted;
assign local_bb4_c0_enter60_c0_eni16_inc_pipelined_thread = 1'b1;
assign local_bb4_c0_enter60_c0_eni16_dec_pipelined_thread = ~(1'b0);
assign local_bb4_c0_enter60_c0_eni16_fu_stall_out = (~(local_bb4_c0_enter60_c0_eni16_inputs_ready) | local_bb4_c0_exit87_c0_exi1386_entry_stall);
assign local_bb4_c0_enter60_c0_eni16_stall_local = (local_bb4_c0_ene161_stall_in | local_bb4_c0_ene262_stall_in | local_bb4_c0_ene363_stall_in | local_bb4_c0_ene464_stall_in | local_bb4_c0_ene565_stall_in | local_bb4_c0_ene666_stall_in | local_bb4_c0_ene767_stall_in | local_bb4_c0_ene868_stall_in | local_bb4_c0_ene969_stall_in | local_bb4_c0_ene1070_stall_in | local_bb4_c0_ene1171_stall_in | local_bb4_c0_ene1272_stall_in | local_bb4_c0_ene1373_stall_in | local_bb4_c0_ene14_stall_in | local_bb4_c0_ene15_stall_in | local_bb4_c0_ene16_stall_in | SFC_2_VALID_1_1_0_stall_in);
assign local_bb4_c0_ene161_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene262_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene363_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene464_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene565_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene666_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene767_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene868_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene969_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene1070_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene1171_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene1272_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene1373_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene14_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene15_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign local_bb4_c0_ene16_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign SFC_2_VALID_1_1_0_valid_out = local_bb4_c0_enter60_c0_eni16_inputs_ready;
assign merge_node_stall_in_0 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_1 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_2 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_3 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_4 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_5 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_6 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_7 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_8 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_9 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_10 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_11 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_12 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_13 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_14 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));
assign merge_node_stall_in_15 = (local_bb4_c0_enter60_c0_eni16_fu_stall_out | ~(local_bb4_c0_enter60_c0_eni16_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene161_stall_local;
wire local_bb4_c0_ene161;

assign local_bb4_c0_ene161 = local_bb4_c0_enter60_c0_eni16[8];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene262_stall_local;
wire local_bb4_c0_ene262;

assign local_bb4_c0_ene262 = local_bb4_c0_enter60_c0_eni16[16];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene363_stall_local;
wire [31:0] local_bb4_c0_ene363;

assign local_bb4_c0_ene363 = local_bb4_c0_enter60_c0_eni16[63:32];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene464_stall_local;
wire [31:0] local_bb4_c0_ene464;

assign local_bb4_c0_ene464 = local_bb4_c0_enter60_c0_eni16[95:64];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene565_stall_local;
wire local_bb4_c0_ene565;

assign local_bb4_c0_ene565 = local_bb4_c0_enter60_c0_eni16[96];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene666_stall_local;
wire [31:0] local_bb4_c0_ene666;

assign local_bb4_c0_ene666 = local_bb4_c0_enter60_c0_eni16[159:128];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene767_stall_local;
wire [31:0] local_bb4_c0_ene767;

assign local_bb4_c0_ene767 = local_bb4_c0_enter60_c0_eni16[191:160];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene868_stall_local;
wire [31:0] local_bb4_c0_ene868;

assign local_bb4_c0_ene868 = local_bb4_c0_enter60_c0_eni16[223:192];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene969_stall_local;
wire local_bb4_c0_ene969;

assign local_bb4_c0_ene969 = local_bb4_c0_enter60_c0_eni16[224];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene1070_stall_local;
wire local_bb4_c0_ene1070;

assign local_bb4_c0_ene1070 = local_bb4_c0_enter60_c0_eni16[232];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene1171_stall_local;
wire local_bb4_c0_ene1171;

assign local_bb4_c0_ene1171 = local_bb4_c0_enter60_c0_eni16[240];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene1272_stall_local;
wire [31:0] local_bb4_c0_ene1272;

assign local_bb4_c0_ene1272 = local_bb4_c0_enter60_c0_eni16[287:256];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene1373_stall_local;
wire [63:0] local_bb4_c0_ene1373;

assign local_bb4_c0_ene1373 = local_bb4_c0_enter60_c0_eni16[383:320];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene14_stall_local;
wire local_bb4_c0_ene14;

assign local_bb4_c0_ene14 = local_bb4_c0_enter60_c0_eni16[384];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene15_stall_local;
wire local_bb4_c0_ene15;

assign local_bb4_c0_ene15 = local_bb4_c0_enter60_c0_eni16[392];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene16_stall_local;
wire local_bb4_c0_ene16;

assign local_bb4_c0_ene16 = local_bb4_c0_enter60_c0_eni16[400];

// This section implements an unregistered operation.
// 
wire SFC_2_VALID_1_1_0_stall_local;
wire SFC_2_VALID_1_1_0;

assign SFC_2_VALID_1_1_0 = local_bb4_c0_enter60_c0_eni16_valid_bit;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene161_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene161_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene161_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene161_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene161_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene161_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene161_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene161_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene161_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene161_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene161_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene161_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene161_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene161),
	.data_out(rnode_1to2_bb4_c0_ene161_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene161_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene161_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene161_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene161_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene161_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene161_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene161_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene161_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene161_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene161_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene262_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene262_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene262_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene262_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene262_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene262_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene262_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene262_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene262_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene262_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene262_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene262_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene262_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene262),
	.data_out(rnode_1to2_bb4_c0_ene262_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene262_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene262_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene262_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene262_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene262_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene262_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene262_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene262_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene262_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene262_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene363_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene363_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene363_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene363_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene363_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene363_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene363_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene363_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene363_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene363_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene363_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene363_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene363_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene363),
	.data_out(rnode_1to2_bb4_c0_ene363_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene363_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene363_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene363_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene363_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene363_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene363_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene363_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene363_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene363_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene363_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene464_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene464_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene464_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene464_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene464_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene464_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene464_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene464_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene464_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene464_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene464_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene464_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene464_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene464),
	.data_out(rnode_1to2_bb4_c0_ene464_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene464_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene464_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene464_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene464_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene464_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene464_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene464_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene464_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene464_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene464_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene565_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene565_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene565_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene565_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene565_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene565_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene565_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene565_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene565_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene565_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene565_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene565_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene565_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene565),
	.data_out(rnode_1to2_bb4_c0_ene565_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene565_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene565_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene565_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene565_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene565_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene565_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene565_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene565_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene565_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene565_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene666_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene666_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene666_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene666_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene666_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene666_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene666_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene666_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene666_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene666_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene666_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene666_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene666_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene666),
	.data_out(rnode_1to2_bb4_c0_ene666_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene666_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene666_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene666_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene666_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene666_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene666_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene666_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene666_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene666_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene666_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene767_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene767_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene767_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene767_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene767_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene767_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene767_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene767_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene767_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene767_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene767_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene767_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene767_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene767),
	.data_out(rnode_1to2_bb4_c0_ene767_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene767_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene767_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene767_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene767_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene767_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene767_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene767_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene767_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene767_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene767_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene868_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene868_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene868_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene868_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene868_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene868_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene868_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene868_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene868_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene868_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene868_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene868_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene868_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene868),
	.data_out(rnode_1to2_bb4_c0_ene868_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene868_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene868_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene868_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene868_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene868_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene868_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene868_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene868_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene868_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene868_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene969_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene969_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene969_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene969_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene969_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene969_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene969_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene969_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene969_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene969_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene969_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene969_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene969_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene969),
	.data_out(rnode_1to2_bb4_c0_ene969_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene969_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene969_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene969_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene969_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene969_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene969_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene969_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene969_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene969_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene969_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene1070_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1070_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1070_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1070_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1070_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1070_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1070_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1070_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene1070_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene1070_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene1070_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene1070_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene1070_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene1070),
	.data_out(rnode_1to2_bb4_c0_ene1070_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene1070_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene1070_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene1070_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene1070_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene1070_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene1070_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene1070_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene1070_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene1070_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene1070_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene1171_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1171_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1171_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1171_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1171_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1171_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1171_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1171_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene1171_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene1171_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene1171_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene1171_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene1171_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene1171),
	.data_out(rnode_1to2_bb4_c0_ene1171_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene1171_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene1171_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene1171_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene1171_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene1171_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene1171_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene1171_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene1171_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene1171_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene1171_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene1272_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1272_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene1272_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1272_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene1272_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1272_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1272_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1272_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene1272_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene1272_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene1272_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene1272_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene1272_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene1272),
	.data_out(rnode_1to2_bb4_c0_ene1272_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene1272_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene1272_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene1272_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene1272_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene1272_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene1272_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene1272_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene1272_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene1272_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene1272_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene1373_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1373_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb4_c0_ene1373_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1373_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb4_c0_ene1373_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1373_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1373_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene1373_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene1373_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene1373_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene1373_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene1373_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene1373_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene1373),
	.data_out(rnode_1to2_bb4_c0_ene1373_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene1373_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene1373_0_reg_2_fifo.DATA_WIDTH = 64;
defparam rnode_1to2_bb4_c0_ene1373_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene1373_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene1373_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene1373_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene1373_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene1373_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene1373_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene1373_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene14_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene14_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene14_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene14_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene14_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene14_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene14_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene14_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene14_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene14_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene14_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene14_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene14_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene14),
	.data_out(rnode_1to2_bb4_c0_ene14_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene14_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene14_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene14_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene14_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene14_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene14_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene14_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene14_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene14_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene14_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene15_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene15_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene15_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene15_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene15_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene15_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene15_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene15_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene15_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene15_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene15_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene15_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene15_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene15),
	.data_out(rnode_1to2_bb4_c0_ene15_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene15_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene15_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene15_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene15_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene15_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene15_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene15_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene15_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene15_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene15_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene16_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene16_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene16_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene16_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene16_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene16_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene16_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene16_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene16_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene16_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene16_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene16_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene16_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene16),
	.data_out(rnode_1to2_bb4_c0_ene16_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene16_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene16_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene16_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene16_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene16_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene16_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene16_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene16_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene16_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene16_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_1_2_0_inputs_ready;
 reg SFC_2_VALID_1_2_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_1_2_0_stall_in;
wire SFC_2_VALID_1_2_0_output_regs_ready;
 reg SFC_2_VALID_1_2_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_1_2_0_causedstall;

assign SFC_2_VALID_1_2_0_inputs_ready = 1'b1;
assign SFC_2_VALID_1_2_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_1_1_0_stall_in = 1'b0;
assign SFC_2_VALID_1_2_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_1_2_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_1_2_0_output_regs_ready)
		begin
			SFC_2_VALID_1_2_0_NO_SHIFT_REG <= SFC_2_VALID_1_1_0;
		end
	end
end


// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_2to8_bb4_c0_ene161_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene161_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene161_0_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene161_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene161_0_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene161_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene161_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene161_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_2to8_bb4_c0_ene161_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to8_bb4_c0_ene161_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to8_bb4_c0_ene161_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_2to8_bb4_c0_ene161_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_2to8_bb4_c0_ene161_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene161_0_NO_SHIFT_REG),
	.data_out(rnode_2to8_bb4_c0_ene161_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_2to8_bb4_c0_ene161_0_reg_8_fifo.DEPTH = 6;
defparam rnode_2to8_bb4_c0_ene161_0_reg_8_fifo.DATA_WIDTH = 1;
defparam rnode_2to8_bb4_c0_ene161_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to8_bb4_c0_ene161_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_2to8_bb4_c0_ene161_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene161_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene161_0_NO_SHIFT_REG = rnode_2to8_bb4_c0_ene161_0_reg_8_NO_SHIFT_REG;
assign rnode_2to8_bb4_c0_ene161_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene161_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_2to6_bb4_c0_ene262_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene262_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene262_0_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene262_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene262_0_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene262_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene262_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene262_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_2to6_bb4_c0_ene262_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to6_bb4_c0_ene262_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to6_bb4_c0_ene262_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_2to6_bb4_c0_ene262_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_2to6_bb4_c0_ene262_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene262_0_NO_SHIFT_REG),
	.data_out(rnode_2to6_bb4_c0_ene262_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_2to6_bb4_c0_ene262_0_reg_6_fifo.DEPTH = 4;
defparam rnode_2to6_bb4_c0_ene262_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_2to6_bb4_c0_ene262_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to6_bb4_c0_ene262_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_2to6_bb4_c0_ene262_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene262_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to6_bb4_c0_ene262_0_NO_SHIFT_REG = rnode_2to6_bb4_c0_ene262_0_reg_6_NO_SHIFT_REG;
assign rnode_2to6_bb4_c0_ene262_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_2to6_bb4_c0_ene262_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_2to6_bb4_c0_ene363_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene363_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to6_bb4_c0_ene363_0_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene363_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to6_bb4_c0_ene363_0_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene363_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene363_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_2to6_bb4_c0_ene363_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_2to6_bb4_c0_ene363_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to6_bb4_c0_ene363_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to6_bb4_c0_ene363_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_2to6_bb4_c0_ene363_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_2to6_bb4_c0_ene363_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene363_0_NO_SHIFT_REG),
	.data_out(rnode_2to6_bb4_c0_ene363_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_2to6_bb4_c0_ene363_0_reg_6_fifo.DEPTH = 4;
defparam rnode_2to6_bb4_c0_ene363_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_2to6_bb4_c0_ene363_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to6_bb4_c0_ene363_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_2to6_bb4_c0_ene363_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene363_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to6_bb4_c0_ene363_0_NO_SHIFT_REG = rnode_2to6_bb4_c0_ene363_0_reg_6_NO_SHIFT_REG;
assign rnode_2to6_bb4_c0_ene363_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_2to6_bb4_c0_ene363_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_2to8_bb4_c0_ene464_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene464_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to8_bb4_c0_ene464_0_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene464_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to8_bb4_c0_ene464_0_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene464_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene464_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene464_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_2to8_bb4_c0_ene464_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to8_bb4_c0_ene464_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to8_bb4_c0_ene464_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_2to8_bb4_c0_ene464_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_2to8_bb4_c0_ene464_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene464_0_NO_SHIFT_REG),
	.data_out(rnode_2to8_bb4_c0_ene464_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_2to8_bb4_c0_ene464_0_reg_8_fifo.DEPTH = 6;
defparam rnode_2to8_bb4_c0_ene464_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_2to8_bb4_c0_ene464_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to8_bb4_c0_ene464_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_2to8_bb4_c0_ene464_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene464_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene464_0_NO_SHIFT_REG = rnode_2to8_bb4_c0_ene464_0_reg_8_NO_SHIFT_REG;
assign rnode_2to8_bb4_c0_ene464_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene464_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene565_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene565_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene565_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene565_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene565_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene565_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene565_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene565_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene565_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene565_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene565_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene565_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene565_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene565_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene565_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene565_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene565_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene565_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene565_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene565_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene565_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene565_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene565_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene565_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene565_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene666_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene666_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene666_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene666_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene666_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene666_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene666_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene666_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene666_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene666_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene666_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene666_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene666_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene666_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene666_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene666_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene666_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_2to9_bb4_c0_ene666_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene666_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene666_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene666_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene666_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene666_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene666_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene666_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene767_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene767_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene767_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene767_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene767_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene767_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene767_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene767_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene767_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene767_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene767_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene767_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene767_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene767_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene767_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene767_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene767_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_2to9_bb4_c0_ene767_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene767_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene767_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene767_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene767_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene767_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene767_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene767_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene868_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene868_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene868_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene868_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene868_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene868_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene868_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene868_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene868_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene868_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene868_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene868_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene868_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene868_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene868_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene868_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene868_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_2to9_bb4_c0_ene868_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene868_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene868_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene868_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene868_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene868_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene868_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene868_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene969_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene969_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene969_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene969_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene969_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene969_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene969_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene969_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene969_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene969_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene969_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene969_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene969_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene969_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene969_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene969_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene969_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene969_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene969_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene969_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene969_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene969_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene969_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene969_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene969_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene1070_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1070_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1070_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1070_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1070_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1070_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1070_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1070_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene1070_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene1070_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene1070_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene1070_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene1070_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene1070_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene1070_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene1070_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene1070_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene1070_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene1070_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene1070_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene1070_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1070_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene1070_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene1070_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1070_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene1171_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1171_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1171_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1171_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1171_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1171_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1171_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1171_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene1171_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene1171_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene1171_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene1171_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene1171_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene1171_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene1171_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene1171_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene1171_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene1171_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene1171_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene1171_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene1171_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1171_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene1171_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene1171_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1171_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene1272_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1272_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene1272_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1272_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to9_bb4_c0_ene1272_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1272_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1272_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1272_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene1272_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene1272_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene1272_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene1272_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene1272_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene1272_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene1272_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene1272_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene1272_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_2to9_bb4_c0_ene1272_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene1272_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene1272_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene1272_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1272_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene1272_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene1272_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1272_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene1373_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1373_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_2to9_bb4_c0_ene1373_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1373_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_2to9_bb4_c0_ene1373_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1373_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1373_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene1373_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene1373_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene1373_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene1373_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene1373_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene1373_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene1373_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene1373_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene1373_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene1373_0_reg_9_fifo.DATA_WIDTH = 64;
defparam rnode_2to9_bb4_c0_ene1373_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene1373_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene1373_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene1373_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1373_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene1373_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene1373_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene1373_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene14_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene14_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene14_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene14_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene14_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene14_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene14_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene14_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene14_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene14_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene14_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene14_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene14_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene14_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene14_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene14_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene14_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene14_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene14_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene14_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene14_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene14_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene14_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene14_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene14_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene15_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene15_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene15_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene15_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene15_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene15_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene15_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene15_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene15_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene15_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene15_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene15_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene15_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene15_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene15_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene15_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene15_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene15_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene15_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene15_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene15_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene15_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene15_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene15_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene15_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene16_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene16_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene16_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene16_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene16_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene16_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene16_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene16_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene16_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene16_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene16_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene16_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene16_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene16_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene16_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene16_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene16_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene16_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene16_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene16_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene16_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene16_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene16_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene16_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene16_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_2_3_0_inputs_ready;
 reg SFC_2_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_2_3_0_stall_in;
wire SFC_2_VALID_2_3_0_output_regs_ready;
 reg SFC_2_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_2_3_0_causedstall;

assign SFC_2_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_1_2_0_stall_in = 1'b0;
assign SFC_2_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_2_3_0_output_regs_ready)
		begin
			SFC_2_VALID_2_3_0_NO_SHIFT_REG <= SFC_2_VALID_1_2_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_c0_ene161_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_valid_out_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_stall_in_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene161_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_c0_ene161_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_c0_ene161_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_c0_ene161_0_stall_in_0_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_c0_ene161_0_valid_out_0_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_c0_ene161_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_2to8_bb4_c0_ene161_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_c0_ene161_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_c0_ene161_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_c0_ene161_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_c0_ene161_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_c0_ene161_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_c0_ene161_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to8_bb4_c0_ene161_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene161_0_stall_in_0_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene161_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_c0_ene161_0_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene161_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_c0_ene161_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_c0_ene161_1_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene161_0_reg_9_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_1_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_2_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_valid_out_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_stall_in_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene262_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_c0_ene262_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_c0_ene262_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_c0_ene262_0_stall_in_0_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_c0_ene262_0_valid_out_0_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_c0_ene262_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(rnode_2to6_bb4_c0_ene262_0_NO_SHIFT_REG),
	.data_out(rnode_6to7_bb4_c0_ene262_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_c0_ene262_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_c0_ene262_0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_6to7_bb4_c0_ene262_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_c0_ene262_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_c0_ene262_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to6_bb4_c0_ene262_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene262_0_stall_in_0_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene262_0_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene262_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene262_1_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene262_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_c0_ene262_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene262_2_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene262_0_reg_7_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_c0_ene363_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene363_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_c0_ene363_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene363_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_c0_ene363_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene363_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene363_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene363_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_c0_ene363_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_c0_ene363_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_c0_ene363_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_c0_ene363_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_c0_ene363_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(rnode_2to6_bb4_c0_ene363_0_NO_SHIFT_REG),
	.data_out(rnode_6to7_bb4_c0_ene363_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_c0_ene363_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_c0_ene363_0_reg_7_fifo.DATA_WIDTH = 32;
defparam rnode_6to7_bb4_c0_ene363_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_c0_ene363_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_c0_ene363_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to6_bb4_c0_ene363_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene363_0_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene363_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_c0_ene363_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene363_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_c0_ene464_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene464_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_c0_ene464_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene464_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_c0_ene464_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene464_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene464_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene464_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_c0_ene464_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_c0_ene464_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_c0_ene464_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_c0_ene464_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_c0_ene464_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_2to8_bb4_c0_ene464_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_c0_ene464_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_c0_ene464_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_c0_ene464_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4_c0_ene464_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_c0_ene464_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_c0_ene464_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to8_bb4_c0_ene464_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene464_0_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene464_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_c0_ene464_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene464_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene565_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene565_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene565_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene565_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene565_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene565_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene565_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene565_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene565_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene565_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene565_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene565_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene565_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene565_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene565_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene565_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene565_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene565_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene565_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene565_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene565_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene565_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene565_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene565_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene565_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene666_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene666_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene666_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene666_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene666_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene666_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene666_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene666_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene666_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene666_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene666_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene666_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene666_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene666_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene666_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene666_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene666_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_c0_ene666_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene666_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene666_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene666_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene666_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene666_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene666_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene666_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene767_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene767_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene767_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene767_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene767_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene767_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene767_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene767_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene767_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene767_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene767_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene767_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene767_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene767_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene767_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene767_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene767_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_c0_ene767_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene767_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene767_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene767_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene767_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene767_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene767_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene767_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene868_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene868_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene868_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene868_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene868_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene868_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene868_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene868_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene868_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene868_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene868_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene868_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene868_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene868_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene868_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene868_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene868_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_c0_ene868_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene868_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene868_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene868_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene868_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene868_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene868_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene868_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene969_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene969_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene969_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene969_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene969_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene969_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene969_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene969_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene969_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene969_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene969_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene969_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene969_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene969_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene969_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene969_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene969_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene969_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene969_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene969_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene969_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene969_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene969_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene969_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene969_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene1070_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1070_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1070_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1070_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1070_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1070_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1070_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1070_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene1070_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene1070_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene1070_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene1070_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene1070_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene1070_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene1070_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene1070_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene1070_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene1070_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene1070_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene1070_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene1070_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1070_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene1070_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene1070_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1070_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene1171_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1171_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1171_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1171_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1171_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1171_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1171_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1171_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene1171_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene1171_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene1171_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene1171_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene1171_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene1171_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene1171_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene1171_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene1171_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene1171_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene1171_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene1171_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene1171_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1171_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene1171_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene1171_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1171_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene1272_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1272_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene1272_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1272_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_c0_ene1272_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1272_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1272_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1272_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene1272_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene1272_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene1272_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene1272_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene1272_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene1272_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene1272_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene1272_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene1272_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_c0_ene1272_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene1272_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene1272_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene1272_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1272_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene1272_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene1272_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1272_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene1373_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1373_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_9to10_bb4_c0_ene1373_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1373_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_9to10_bb4_c0_ene1373_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1373_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1373_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene1373_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene1373_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene1373_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene1373_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene1373_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene1373_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene1373_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene1373_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene1373_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene1373_0_reg_10_fifo.DATA_WIDTH = 64;
defparam rnode_9to10_bb4_c0_ene1373_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene1373_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene1373_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene1373_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1373_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene1373_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene1373_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1373_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene14_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene14_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene14_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene14_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene14_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene14_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene14_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene14_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene14_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene14_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene14_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene14_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene14_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene14_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene14_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene14_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene14_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene14_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene14_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene14_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene14_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene14_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene14_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene14_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene14_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene15_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene15_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene15_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene15_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene15_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene15_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene15_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene15_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene15_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene15_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene15_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene15_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene15_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene15_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene15_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene15_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene15_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene15_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene15_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene15_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene15_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene15_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene15_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene15_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene15_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene16_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene16_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene16_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene16_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene16_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene16_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene16_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene16_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene16_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene16_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene16_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene16_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene16_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene16_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene16_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene16_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene16_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene16_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene16_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene16_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene16_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene16_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene16_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene16_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene16_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_3_4_0_inputs_ready;
 reg SFC_2_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_3_4_0_stall_in;
wire SFC_2_VALID_3_4_0_output_regs_ready;
 reg SFC_2_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_3_4_0_causedstall;

assign SFC_2_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_stall_in = 1'b0;
assign SFC_2_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_3_4_0_output_regs_ready)
		begin
			SFC_2_VALID_3_4_0_NO_SHIFT_REG <= SFC_2_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene161_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene161_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene161_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene161_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene161_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene161_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene161_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene161_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene161_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene161_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene161_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene161_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene161_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_8to9_bb4_c0_ene161_1_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene161_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene161_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene161_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene161_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene161_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene161_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_c0_ene161_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene161_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene161_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene161_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene161_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_7to9_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_1_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_valid_out_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_stall_in_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_c0_ene262_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_7to9_bb4_c0_ene262_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to9_bb4_c0_ene262_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to9_bb4_c0_ene262_0_stall_in_0_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_7to9_bb4_c0_ene262_0_valid_out_0_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_7to9_bb4_c0_ene262_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_c0_ene262_2_NO_SHIFT_REG),
	.data_out(rnode_7to9_bb4_c0_ene262_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_7to9_bb4_c0_ene262_0_reg_9_fifo.DEPTH = 2;
defparam rnode_7to9_bb4_c0_ene262_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_7to9_bb4_c0_ene262_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to9_bb4_c0_ene262_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_7to9_bb4_c0_ene262_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene262_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_7to9_bb4_c0_ene262_0_stall_in_0_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_7to9_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene262_0_NO_SHIFT_REG = rnode_7to9_bb4_c0_ene262_0_reg_9_NO_SHIFT_REG;
assign rnode_7to9_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene262_1_NO_SHIFT_REG = rnode_7to9_bb4_c0_ene262_0_reg_9_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_2_VALID_4_5_0_inputs_ready;
 reg SFC_2_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_4_5_0_stall_in;
wire SFC_2_VALID_4_5_0_output_regs_ready;
 reg SFC_2_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_4_5_0_causedstall;

assign SFC_2_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_stall_in = 1'b0;
assign SFC_2_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_4_5_0_output_regs_ready)
		begin
			SFC_2_VALID_4_5_0_NO_SHIFT_REG <= SFC_2_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_2_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_3_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_4_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_4_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_5_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_5_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_5_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_6_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_6_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_6_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_7_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_7_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_7_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_8_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_8_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_8_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_9_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_9_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_9_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_11_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_11_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_11_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_12_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_12_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_12_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_valid_out_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_in_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene262_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene262_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene262_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene262_0_stall_in_0_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene262_0_valid_out_0_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene262_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_7to9_bb4_c0_ene262_1_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene262_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene262_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene262_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene262_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene262_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_c0_ene262_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_0_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_1_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_2_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_3_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_4_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_5_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_5_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_6_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_6_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_7_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_7_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_8_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_8_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_9_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_9_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_10_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_10_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_11_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_11_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene262_0_valid_out_12_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene262_12_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene262_0_reg_10_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_2_VALID_5_6_0_inputs_ready;
 reg SFC_2_VALID_5_6_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_5_6_0_stall_in;
wire SFC_2_VALID_5_6_0_output_regs_ready;
 reg SFC_2_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_5_6_0_causedstall;

assign SFC_2_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_stall_in = 1'b0;
assign SFC_2_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_5_6_0_output_regs_ready)
		begin
			SFC_2_VALID_5_6_0_NO_SHIFT_REG <= SFC_2_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_6_7_0_inputs_ready;
 reg SFC_2_VALID_6_7_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_6_7_0_stall_in_0;
 reg SFC_2_VALID_6_7_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_6_7_0_stall_in_1;
 reg SFC_2_VALID_6_7_0_valid_out_2_NO_SHIFT_REG;
wire SFC_2_VALID_6_7_0_stall_in_2;
wire SFC_2_VALID_6_7_0_output_regs_ready;
 reg SFC_2_VALID_6_7_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_6_7_0_causedstall;

assign SFC_2_VALID_6_7_0_inputs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_stall_in = 1'b0;
assign SFC_2_VALID_6_7_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_6_7_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_6_7_0_output_regs_ready)
		begin
			SFC_2_VALID_6_7_0_NO_SHIFT_REG <= SFC_2_VALID_5_6_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_2_VALID_7_8_0_inputs_ready;
 reg SFC_2_VALID_7_8_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_7_8_0_stall_in;
wire SFC_2_VALID_7_8_0_output_regs_ready;
 reg SFC_2_VALID_7_8_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_7_8_0_causedstall;

assign SFC_2_VALID_7_8_0_inputs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_7_8_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_7_8_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_7_8_0_output_regs_ready)
		begin
			SFC_2_VALID_7_8_0_NO_SHIFT_REG <= SFC_2_VALID_6_7_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_j_35_pop30_add7_stall_local;
wire [31:0] local_bb4_j_35_pop30_add7;
wire local_bb4_j_35_pop30_add7_fu_valid_out;
wire local_bb4_j_35_pop30_add7_fu_stall_out;

acl_pop local_bb4_j_35_pop30_add7_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_6to7_bb4_c0_ene262_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(input_wii_add7),
	.stall_out(local_bb4_j_35_pop30_add7_fu_stall_out),
	.valid_in(SFC_2_VALID_6_7_0_NO_SHIFT_REG),
	.valid_out(local_bb4_j_35_pop30_add7_fu_valid_out),
	.stall_in(local_bb4_j_35_pop30_add7_stall_local),
	.data_out(local_bb4_j_35_pop30_add7),
	.feedback_in(feedback_data_in_30),
	.feedback_valid_in(feedback_valid_in_30),
	.feedback_stall_out(feedback_stall_out_30)
);

defparam local_bb4_j_35_pop30_add7_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_j_35_pop30_add7_feedback.DATA_WIDTH = 32;
defparam local_bb4_j_35_pop30_add7_feedback.STYLE = "REGULAR";

assign local_bb4_j_35_pop30_add7_stall_local = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__pop40_c0_ene363_stall_local;
wire [31:0] local_bb4__pop40_c0_ene363;
wire local_bb4__pop40_c0_ene363_fu_valid_out;
wire local_bb4__pop40_c0_ene363_fu_stall_out;

acl_pop local_bb4__pop40_c0_ene363_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_6to7_bb4_c0_ene262_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_6to7_bb4_c0_ene363_0_NO_SHIFT_REG),
	.stall_out(local_bb4__pop40_c0_ene363_fu_stall_out),
	.valid_in(SFC_2_VALID_6_7_0_NO_SHIFT_REG),
	.valid_out(local_bb4__pop40_c0_ene363_fu_valid_out),
	.stall_in(local_bb4__pop40_c0_ene363_stall_local),
	.data_out(local_bb4__pop40_c0_ene363),
	.feedback_in(feedback_data_in_40),
	.feedback_valid_in(feedback_valid_in_40),
	.feedback_stall_out(feedback_stall_out_40)
);

defparam local_bb4__pop40_c0_ene363_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4__pop40_c0_ene363_feedback.DATA_WIDTH = 32;
defparam local_bb4__pop40_c0_ene363_feedback.STYLE = "REGULAR";

assign local_bb4__pop40_c0_ene363_stall_local = 1'b0;

// This section implements a registered operation.
// 
wire SFC_2_VALID_8_9_0_inputs_ready;
 reg SFC_2_VALID_8_9_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_0;
 reg SFC_2_VALID_8_9_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_1;
 reg SFC_2_VALID_8_9_0_valid_out_2_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_2;
 reg SFC_2_VALID_8_9_0_valid_out_3_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_3;
 reg SFC_2_VALID_8_9_0_valid_out_4_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_4;
wire SFC_2_VALID_8_9_0_output_regs_ready;
 reg SFC_2_VALID_8_9_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_8_9_0_causedstall;

assign SFC_2_VALID_8_9_0_inputs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_stall_in = 1'b0;
assign SFC_2_VALID_8_9_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_8_9_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_8_9_0_output_regs_ready)
		begin
			SFC_2_VALID_8_9_0_NO_SHIFT_REG <= SFC_2_VALID_7_8_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_inc_stall_local;
wire [31:0] local_bb4_inc;

assign local_bb4_inc = (local_bb4_j_35_pop30_add7 + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_add16_valid_out;
wire local_bb4_add16_stall_in;
wire local_bb4_inc_valid_out;
wire local_bb4_inc_stall_in;
wire local_bb4__pop40_c0_ene363_valid_out_1;
wire local_bb4__pop40_c0_ene363_stall_in_1;
wire local_bb4_add16_inputs_ready;
wire local_bb4_add16_stall_local;
wire [31:0] local_bb4_add16;

assign local_bb4_add16_inputs_ready = (SFC_2_VALID_6_7_0_valid_out_1_NO_SHIFT_REG & rnode_6to7_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG & SFC_2_VALID_6_7_0_valid_out_2_NO_SHIFT_REG & rnode_6to7_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG & rnode_6to7_bb4_c0_ene363_0_valid_out_NO_SHIFT_REG);
assign local_bb4_add16 = (local_bb4_j_35_pop30_add7 + local_bb4__pop40_c0_ene363);
assign local_bb4_add16_valid_out = 1'b1;
assign local_bb4_inc_valid_out = 1'b1;
assign local_bb4__pop40_c0_ene363_valid_out_1 = 1'b1;
assign SFC_2_VALID_6_7_0_stall_in_1 = 1'b0;
assign rnode_6to7_bb4_c0_ene262_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign SFC_2_VALID_6_7_0_stall_in_2 = 1'b0;
assign rnode_6to7_bb4_c0_ene262_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene363_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_2_VALID_9_10_0_inputs_ready;
 reg SFC_2_VALID_9_10_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_0;
 reg SFC_2_VALID_9_10_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_1;
 reg SFC_2_VALID_9_10_0_valid_out_2_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_2;
 reg SFC_2_VALID_9_10_0_valid_out_3_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_3;
 reg SFC_2_VALID_9_10_0_valid_out_4_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_4;
 reg SFC_2_VALID_9_10_0_valid_out_5_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_5;
 reg SFC_2_VALID_9_10_0_valid_out_6_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_6;
 reg SFC_2_VALID_9_10_0_valid_out_7_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_7;
 reg SFC_2_VALID_9_10_0_valid_out_8_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_8;
 reg SFC_2_VALID_9_10_0_valid_out_9_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_9;
 reg SFC_2_VALID_9_10_0_valid_out_10_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_10;
 reg SFC_2_VALID_9_10_0_valid_out_11_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_11;
 reg SFC_2_VALID_9_10_0_valid_out_12_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_12;
 reg SFC_2_VALID_9_10_0_valid_out_13_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_13;
 reg SFC_2_VALID_9_10_0_valid_out_14_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_14;
 reg SFC_2_VALID_9_10_0_valid_out_15_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_15;
 reg SFC_2_VALID_9_10_0_valid_out_16_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_16;
 reg SFC_2_VALID_9_10_0_valid_out_17_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_17;
 reg SFC_2_VALID_9_10_0_valid_out_18_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_18;
 reg SFC_2_VALID_9_10_0_valid_out_19_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_19;
 reg SFC_2_VALID_9_10_0_valid_out_20_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_20;
 reg SFC_2_VALID_9_10_0_valid_out_21_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_21;
 reg SFC_2_VALID_9_10_0_valid_out_22_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_22;
 reg SFC_2_VALID_9_10_0_valid_out_23_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_23;
 reg SFC_2_VALID_9_10_0_valid_out_24_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_24;
 reg SFC_2_VALID_9_10_0_valid_out_25_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_25;
 reg SFC_2_VALID_9_10_0_valid_out_26_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_26;
 reg SFC_2_VALID_9_10_0_valid_out_27_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_27;
 reg SFC_2_VALID_9_10_0_valid_out_28_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_28;
wire SFC_2_VALID_9_10_0_output_regs_ready;
 reg SFC_2_VALID_9_10_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_9_10_0_causedstall;

assign SFC_2_VALID_9_10_0_inputs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_9_10_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_9_10_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_9_10_0_output_regs_ready)
		begin
			SFC_2_VALID_9_10_0_NO_SHIFT_REG <= SFC_2_VALID_8_9_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_keep_going_acl_pipeline_1_inputs_ready;
 reg local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb4_keep_going_acl_pipeline_1_stall_in;
wire local_bb4_keep_going_acl_pipeline_1_output_regs_ready;
wire local_bb4_keep_going_acl_pipeline_1_keep_going;
wire local_bb4_keep_going_acl_pipeline_1_fu_valid_out;
wire local_bb4_keep_going_acl_pipeline_1_fu_stall_out;
 reg local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb4_keep_going_acl_pipeline_1_feedback_pipelined;
wire local_bb4_keep_going_acl_pipeline_1_causedstall;

acl_pipeline local_bb4_keep_going_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb4_keep_going_acl_pipeline_1_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_keep_going_acl_pipeline_1_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_keep_going_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_0),
	.not_exitcond_in(feedback_data_in_1),
	.not_exitcond_valid_in(feedback_valid_in_1),
	.not_exitcond_stall_out(feedback_stall_out_1),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb4_keep_going_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb4_keep_going_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb4_keep_going_acl_pipeline_1_inputs_ready = 1'b1;
assign local_bb4_keep_going_acl_pipeline_1_output_regs_ready = 1'b1;
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign SFC_2_VALID_8_9_0_stall_in_1 = 1'b0;
assign rnode_8to9_bb4_c0_ene161_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb4_keep_going_acl_pipeline_1_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_keep_going_acl_pipeline_1_output_regs_ready)
		begin
			local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG <= local_bb4_keep_going_acl_pipeline_1_keep_going;
			local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_keep_going_acl_pipeline_1_stall_in))
			begin
				local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_mul2445_pop46_c0_ene464_stall_local;
wire [31:0] local_bb4_mul2445_pop46_c0_ene464;
wire local_bb4_mul2445_pop46_c0_ene464_fu_valid_out;
wire local_bb4_mul2445_pop46_c0_ene464_fu_stall_out;

acl_pop local_bb4_mul2445_pop46_c0_ene464_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_7to9_bb4_c0_ene262_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_8to9_bb4_c0_ene464_0_NO_SHIFT_REG),
	.stall_out(local_bb4_mul2445_pop46_c0_ene464_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_mul2445_pop46_c0_ene464_fu_valid_out),
	.stall_in(local_bb4_mul2445_pop46_c0_ene464_stall_local),
	.data_out(local_bb4_mul2445_pop46_c0_ene464),
	.feedback_in(feedback_data_in_46),
	.feedback_valid_in(feedback_valid_in_46),
	.feedback_stall_out(feedback_stall_out_46)
);

defparam local_bb4_mul2445_pop46_c0_ene464_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_mul2445_pop46_c0_ene464_feedback.DATA_WIDTH = 32;
defparam local_bb4_mul2445_pop46_c0_ene464_feedback.STYLE = "REGULAR";

assign local_bb4_mul2445_pop46_c0_ene464_stall_local = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_add16_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add16_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add16_1_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add16_2_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add16_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_valid_out_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_stall_in_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add16_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_add16_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_add16_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_add16_0_stall_in_0_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_add16_0_valid_out_0_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_add16_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_bb4_add16),
	.data_out(rnode_7to8_bb4_add16_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_add16_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_add16_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_7to8_bb4_add16_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_add16_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_add16_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add16_stall_in = 1'b0;
assign rnode_7to8_bb4_add16_0_stall_in_0_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_add16_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add16_0_NO_SHIFT_REG = rnode_7to8_bb4_add16_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_add16_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add16_1_NO_SHIFT_REG = rnode_7to8_bb4_add16_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_add16_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add16_2_NO_SHIFT_REG = rnode_7to8_bb4_add16_0_reg_8_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_inc_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_inc_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_inc_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_inc_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_7to8_bb4_inc_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_inc_1_NO_SHIFT_REG;
 logic rnode_7to8_bb4_inc_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_inc_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_inc_0_valid_out_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_inc_0_stall_in_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_inc_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_inc_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_inc_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_inc_0_stall_in_0_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_inc_0_valid_out_0_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_inc_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_bb4_inc),
	.data_out(rnode_7to8_bb4_inc_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_inc_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_inc_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_7to8_bb4_inc_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_inc_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_inc_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_inc_stall_in = 1'b0;
assign rnode_7to8_bb4_inc_0_stall_in_0_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_inc_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_inc_0_NO_SHIFT_REG = rnode_7to8_bb4_inc_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_inc_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_inc_1_NO_SHIFT_REG = rnode_7to8_bb4_inc_0_reg_8_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4__pop40_c0_ene363_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb4__pop40_c0_ene363_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4__pop40_c0_ene363_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4__pop40_c0_ene363_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4__pop40_c0_ene363_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4__pop40_c0_ene363_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4__pop40_c0_ene363_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4__pop40_c0_ene363_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4__pop40_c0_ene363_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_bb4__pop40_c0_ene363),
	.data_out(rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__pop40_c0_ene363_stall_in_1 = 1'b0;
assign rnode_7to8_bb4__pop40_c0_ene363_0_NO_SHIFT_REG = rnode_7to8_bb4__pop40_c0_ene363_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4__pop40_c0_ene363_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4__pop40_c0_ene363_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_10_11_0_inputs_ready;
 reg SFC_2_VALID_10_11_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_10_11_0_stall_in;
wire SFC_2_VALID_10_11_0_output_regs_ready;
 reg SFC_2_VALID_10_11_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_10_11_0_causedstall;

assign SFC_2_VALID_10_11_0_inputs_ready = 1'b1;
assign SFC_2_VALID_10_11_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_10_11_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_10_11_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_10_11_0_output_regs_ready)
		begin
			SFC_2_VALID_10_11_0_NO_SHIFT_REG <= SFC_2_VALID_9_10_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_forked1644_pop45_c0_ene161_valid_out_0;
wire local_bb4_forked1644_pop45_c0_ene161_stall_in_0;
wire local_bb4_forked1644_pop45_c0_ene161_valid_out_1;
wire local_bb4_forked1644_pop45_c0_ene161_stall_in_1;
wire local_bb4_forked1644_pop45_c0_ene161_inputs_ready;
wire local_bb4_forked1644_pop45_c0_ene161_stall_local;
wire local_bb4_forked1644_pop45_c0_ene161;
wire local_bb4_forked1644_pop45_c0_ene161_fu_valid_out;
wire local_bb4_forked1644_pop45_c0_ene161_fu_stall_out;

acl_pop local_bb4_forked1644_pop45_c0_ene161_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene161_0_NO_SHIFT_REG),
	.stall_out(local_bb4_forked1644_pop45_c0_ene161_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_forked1644_pop45_c0_ene161_fu_valid_out),
	.stall_in(local_bb4_forked1644_pop45_c0_ene161_stall_local),
	.data_out(local_bb4_forked1644_pop45_c0_ene161),
	.feedback_in(feedback_data_in_45),
	.feedback_valid_in(feedback_valid_in_45),
	.feedback_stall_out(feedback_stall_out_45)
);

defparam local_bb4_forked1644_pop45_c0_ene161_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_forked1644_pop45_c0_ene161_feedback.DATA_WIDTH = 1;
defparam local_bb4_forked1644_pop45_c0_ene161_feedback.STYLE = "REGULAR";

assign local_bb4_forked1644_pop45_c0_ene161_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_1_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene161_0_valid_out_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_forked1644_pop45_c0_ene161_stall_local = 1'b0;
assign local_bb4_forked1644_pop45_c0_ene161_valid_out_0 = 1'b1;
assign local_bb4_forked1644_pop45_c0_ene161_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_1 = 1'b0;
assign rnode_9to10_bb4_c0_ene161_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_valid_out_0;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_stall_in_0;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_valid_out_1;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_stall_in_1;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_inputs_ready;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_stall_local;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_fu_valid_out;
wire local_bb4_memdep_phi1_or39_pop41_c0_ene565_fu_stall_out;

acl_pop local_bb4_memdep_phi1_or39_pop41_c0_ene565_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene565_0_NO_SHIFT_REG),
	.stall_out(local_bb4_memdep_phi1_or39_pop41_c0_ene565_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_memdep_phi1_or39_pop41_c0_ene565_fu_valid_out),
	.stall_in(local_bb4_memdep_phi1_or39_pop41_c0_ene565_stall_local),
	.data_out(local_bb4_memdep_phi1_or39_pop41_c0_ene565),
	.feedback_in(feedback_data_in_41),
	.feedback_valid_in(feedback_valid_in_41),
	.feedback_stall_out(feedback_stall_out_41)
);

defparam local_bb4_memdep_phi1_or39_pop41_c0_ene565_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_memdep_phi1_or39_pop41_c0_ene565_feedback.DATA_WIDTH = 1;
defparam local_bb4_memdep_phi1_or39_pop41_c0_ene565_feedback.STYLE = "REGULAR";

assign local_bb4_memdep_phi1_or39_pop41_c0_ene565_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_2_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_1_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene565_0_valid_out_NO_SHIFT_REG);
assign local_bb4_memdep_phi1_or39_pop41_c0_ene565_stall_local = 1'b0;
assign local_bb4_memdep_phi1_or39_pop41_c0_ene565_valid_out_0 = 1'b1;
assign local_bb4_memdep_phi1_or39_pop41_c0_ene565_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_2 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene565_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__pop42_c0_ene666_valid_out_0;
wire local_bb4__pop42_c0_ene666_stall_in_0;
wire local_bb4__pop42_c0_ene666_valid_out_1;
wire local_bb4__pop42_c0_ene666_stall_in_1;
wire local_bb4__pop42_c0_ene666_inputs_ready;
wire local_bb4__pop42_c0_ene666_stall_local;
wire [31:0] local_bb4__pop42_c0_ene666;
wire local_bb4__pop42_c0_ene666_fu_valid_out;
wire local_bb4__pop42_c0_ene666_fu_stall_out;

acl_pop local_bb4__pop42_c0_ene666_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_2_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene666_0_NO_SHIFT_REG),
	.stall_out(local_bb4__pop42_c0_ene666_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__pop42_c0_ene666_fu_valid_out),
	.stall_in(local_bb4__pop42_c0_ene666_stall_local),
	.data_out(local_bb4__pop42_c0_ene666),
	.feedback_in(feedback_data_in_42),
	.feedback_valid_in(feedback_valid_in_42),
	.feedback_stall_out(feedback_stall_out_42)
);

defparam local_bb4__pop42_c0_ene666_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4__pop42_c0_ene666_feedback.DATA_WIDTH = 32;
defparam local_bb4__pop42_c0_ene666_feedback.STYLE = "REGULAR";

assign local_bb4__pop42_c0_ene666_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_3_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_2_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene666_0_valid_out_NO_SHIFT_REG);
assign local_bb4__pop42_c0_ene666_stall_local = 1'b0;
assign local_bb4__pop42_c0_ene666_valid_out_0 = 1'b1;
assign local_bb4__pop42_c0_ene666_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_3 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene666_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_pixel_y_020_pop821_pop33_c0_ene767_valid_out;
wire local_bb4_pixel_y_020_pop821_pop33_c0_ene767_stall_in;
wire local_bb4_pixel_y_020_pop821_pop33_c0_ene767_inputs_ready;
wire local_bb4_pixel_y_020_pop821_pop33_c0_ene767_stall_local;
wire [31:0] local_bb4_pixel_y_020_pop821_pop33_c0_ene767;
wire local_bb4_pixel_y_020_pop821_pop33_c0_ene767_fu_valid_out;
wire local_bb4_pixel_y_020_pop821_pop33_c0_ene767_fu_stall_out;

acl_pop local_bb4_pixel_y_020_pop821_pop33_c0_ene767_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_3_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene767_0_NO_SHIFT_REG),
	.stall_out(local_bb4_pixel_y_020_pop821_pop33_c0_ene767_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_pixel_y_020_pop821_pop33_c0_ene767_fu_valid_out),
	.stall_in(local_bb4_pixel_y_020_pop821_pop33_c0_ene767_stall_local),
	.data_out(local_bb4_pixel_y_020_pop821_pop33_c0_ene767),
	.feedback_in(feedback_data_in_33),
	.feedback_valid_in(feedback_valid_in_33),
	.feedback_stall_out(feedback_stall_out_33)
);

defparam local_bb4_pixel_y_020_pop821_pop33_c0_ene767_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_pixel_y_020_pop821_pop33_c0_ene767_feedback.DATA_WIDTH = 32;
defparam local_bb4_pixel_y_020_pop821_pop33_c0_ene767_feedback.STYLE = "REGULAR";

assign local_bb4_pixel_y_020_pop821_pop33_c0_ene767_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_4_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_3_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene767_0_valid_out_NO_SHIFT_REG);
assign local_bb4_pixel_y_020_pop821_pop33_c0_ene767_stall_local = 1'b0;
assign local_bb4_pixel_y_020_pop821_pop33_c0_ene767_valid_out = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_4 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene767_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_mul3724_pop34_c0_ene868_valid_out_0;
wire local_bb4_mul3724_pop34_c0_ene868_stall_in_0;
wire local_bb4_mul3724_pop34_c0_ene868_valid_out_1;
wire local_bb4_mul3724_pop34_c0_ene868_stall_in_1;
wire local_bb4_mul3724_pop34_c0_ene868_inputs_ready;
wire local_bb4_mul3724_pop34_c0_ene868_stall_local;
wire [31:0] local_bb4_mul3724_pop34_c0_ene868;
wire local_bb4_mul3724_pop34_c0_ene868_fu_valid_out;
wire local_bb4_mul3724_pop34_c0_ene868_fu_stall_out;

acl_pop local_bb4_mul3724_pop34_c0_ene868_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_4_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene868_0_NO_SHIFT_REG),
	.stall_out(local_bb4_mul3724_pop34_c0_ene868_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_mul3724_pop34_c0_ene868_fu_valid_out),
	.stall_in(local_bb4_mul3724_pop34_c0_ene868_stall_local),
	.data_out(local_bb4_mul3724_pop34_c0_ene868),
	.feedback_in(feedback_data_in_34),
	.feedback_valid_in(feedback_valid_in_34),
	.feedback_stall_out(feedback_stall_out_34)
);

defparam local_bb4_mul3724_pop34_c0_ene868_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_mul3724_pop34_c0_ene868_feedback.DATA_WIDTH = 32;
defparam local_bb4_mul3724_pop34_c0_ene868_feedback.STYLE = "REGULAR";

assign local_bb4_mul3724_pop34_c0_ene868_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_5_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_4_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene868_0_valid_out_NO_SHIFT_REG);
assign local_bb4_mul3724_pop34_c0_ene868_stall_local = 1'b0;
assign local_bb4_mul3724_pop34_c0_ene868_valid_out_0 = 1'b1;
assign local_bb4_mul3724_pop34_c0_ene868_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_5 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene868_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notcmp1127_pop35_c0_ene969_valid_out_0;
wire local_bb4_notcmp1127_pop35_c0_ene969_stall_in_0;
wire local_bb4_notcmp1127_pop35_c0_ene969_valid_out_1;
wire local_bb4_notcmp1127_pop35_c0_ene969_stall_in_1;
wire local_bb4_notcmp1127_pop35_c0_ene969_inputs_ready;
wire local_bb4_notcmp1127_pop35_c0_ene969_stall_local;
wire local_bb4_notcmp1127_pop35_c0_ene969;
wire local_bb4_notcmp1127_pop35_c0_ene969_fu_valid_out;
wire local_bb4_notcmp1127_pop35_c0_ene969_fu_stall_out;

acl_pop local_bb4_notcmp1127_pop35_c0_ene969_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_5_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene969_0_NO_SHIFT_REG),
	.stall_out(local_bb4_notcmp1127_pop35_c0_ene969_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notcmp1127_pop35_c0_ene969_fu_valid_out),
	.stall_in(local_bb4_notcmp1127_pop35_c0_ene969_stall_local),
	.data_out(local_bb4_notcmp1127_pop35_c0_ene969),
	.feedback_in(feedback_data_in_35),
	.feedback_valid_in(feedback_valid_in_35),
	.feedback_stall_out(feedback_stall_out_35)
);

defparam local_bb4_notcmp1127_pop35_c0_ene969_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_notcmp1127_pop35_c0_ene969_feedback.DATA_WIDTH = 1;
defparam local_bb4_notcmp1127_pop35_c0_ene969_feedback.STYLE = "REGULAR";

assign local_bb4_notcmp1127_pop35_c0_ene969_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_6_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_5_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene969_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notcmp1127_pop35_c0_ene969_stall_local = 1'b0;
assign local_bb4_notcmp1127_pop35_c0_ene969_valid_out_0 = 1'b1;
assign local_bb4_notcmp1127_pop35_c0_ene969_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_6 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_5_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene969_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notexitcond1430_pop36_c0_ene1070_valid_out_0;
wire local_bb4_notexitcond1430_pop36_c0_ene1070_stall_in_0;
wire local_bb4_notexitcond1430_pop36_c0_ene1070_valid_out_1;
wire local_bb4_notexitcond1430_pop36_c0_ene1070_stall_in_1;
wire local_bb4_notexitcond1430_pop36_c0_ene1070_inputs_ready;
wire local_bb4_notexitcond1430_pop36_c0_ene1070_stall_local;
wire local_bb4_notexitcond1430_pop36_c0_ene1070;
wire local_bb4_notexitcond1430_pop36_c0_ene1070_fu_valid_out;
wire local_bb4_notexitcond1430_pop36_c0_ene1070_fu_stall_out;

acl_pop local_bb4_notexitcond1430_pop36_c0_ene1070_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene1070_0_NO_SHIFT_REG),
	.stall_out(local_bb4_notexitcond1430_pop36_c0_ene1070_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond1430_pop36_c0_ene1070_fu_valid_out),
	.stall_in(local_bb4_notexitcond1430_pop36_c0_ene1070_stall_local),
	.data_out(local_bb4_notexitcond1430_pop36_c0_ene1070),
	.feedback_in(feedback_data_in_36),
	.feedback_valid_in(feedback_valid_in_36),
	.feedback_stall_out(feedback_stall_out_36)
);

defparam local_bb4_notexitcond1430_pop36_c0_ene1070_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_notexitcond1430_pop36_c0_ene1070_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond1430_pop36_c0_ene1070_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond1430_pop36_c0_ene1070_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_7_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_6_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene1070_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notexitcond1430_pop36_c0_ene1070_stall_local = 1'b0;
assign local_bb4_notexitcond1430_pop36_c0_ene1070_valid_out_0 = 1'b1;
assign local_bb4_notexitcond1430_pop36_c0_ene1070_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_7 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_6_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1070_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_valid_out;
wire local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_stall_in;
wire local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_inputs_ready;
wire local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_stall_local;
wire local_bb4_memdep_phi1_pop933_pop37_c0_ene1171;
wire local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_fu_valid_out;
wire local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_fu_stall_out;

acl_pop local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_7_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene1171_0_NO_SHIFT_REG),
	.stall_out(local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_fu_valid_out),
	.stall_in(local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_stall_local),
	.data_out(local_bb4_memdep_phi1_pop933_pop37_c0_ene1171),
	.feedback_in(feedback_data_in_37),
	.feedback_valid_in(feedback_valid_in_37),
	.feedback_stall_out(feedback_stall_out_37)
);

defparam local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_feedback.DATA_WIDTH = 1;
defparam local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_feedback.STYLE = "REGULAR";

assign local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_8_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_7_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene1171_0_valid_out_NO_SHIFT_REG);
assign local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_stall_local = 1'b0;
assign local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_valid_out = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_8 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_7_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1171_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_mul535_pop38_c0_ene1272_valid_out;
wire local_bb4_mul535_pop38_c0_ene1272_stall_in;
wire local_bb4_mul535_pop38_c0_ene1272_inputs_ready;
wire local_bb4_mul535_pop38_c0_ene1272_stall_local;
wire [31:0] local_bb4_mul535_pop38_c0_ene1272;
wire local_bb4_mul535_pop38_c0_ene1272_fu_valid_out;
wire local_bb4_mul535_pop38_c0_ene1272_fu_stall_out;

acl_pop local_bb4_mul535_pop38_c0_ene1272_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_8_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene1272_0_NO_SHIFT_REG),
	.stall_out(local_bb4_mul535_pop38_c0_ene1272_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_mul535_pop38_c0_ene1272_fu_valid_out),
	.stall_in(local_bb4_mul535_pop38_c0_ene1272_stall_local),
	.data_out(local_bb4_mul535_pop38_c0_ene1272),
	.feedback_in(feedback_data_in_38),
	.feedback_valid_in(feedback_valid_in_38),
	.feedback_stall_out(feedback_stall_out_38)
);

defparam local_bb4_mul535_pop38_c0_ene1272_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_mul535_pop38_c0_ene1272_feedback.DATA_WIDTH = 32;
defparam local_bb4_mul535_pop38_c0_ene1272_feedback.STYLE = "REGULAR";

assign local_bb4_mul535_pop38_c0_ene1272_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_9_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_8_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene1272_0_valid_out_NO_SHIFT_REG);
assign local_bb4_mul535_pop38_c0_ene1272_stall_local = 1'b0;
assign local_bb4_mul535_pop38_c0_ene1272_valid_out = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_9 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_8_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1272_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_valid_out_0;
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_stall_in_0;
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_valid_out_1;
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_stall_in_1;
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_inputs_ready;
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_stall_local;
wire [63:0] local_bb4_indvars_iv_pop1037_pop39_c0_ene1373;
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_fu_valid_out;
wire local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_fu_stall_out;

acl_pop local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_9_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene1373_0_NO_SHIFT_REG),
	.stall_out(local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_fu_valid_out),
	.stall_in(local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_stall_local),
	.data_out(local_bb4_indvars_iv_pop1037_pop39_c0_ene1373),
	.feedback_in(feedback_data_in_39),
	.feedback_valid_in(feedback_valid_in_39),
	.feedback_stall_out(feedback_stall_out_39)
);

defparam local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_feedback.DATA_WIDTH = 64;
defparam local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_feedback.STYLE = "REGULAR";

assign local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_10_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_9_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene1373_0_valid_out_NO_SHIFT_REG);
assign local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_stall_local = 1'b0;
assign local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_valid_out_0 = 1'b1;
assign local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_10 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_9_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene1373_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notcmp41_pop43_c0_ene14_valid_out_0;
wire local_bb4_notcmp41_pop43_c0_ene14_stall_in_0;
wire local_bb4_notcmp41_pop43_c0_ene14_valid_out_1;
wire local_bb4_notcmp41_pop43_c0_ene14_stall_in_1;
wire local_bb4_notcmp41_pop43_c0_ene14_inputs_ready;
wire local_bb4_notcmp41_pop43_c0_ene14_stall_local;
wire local_bb4_notcmp41_pop43_c0_ene14;
wire local_bb4_notcmp41_pop43_c0_ene14_fu_valid_out;
wire local_bb4_notcmp41_pop43_c0_ene14_fu_stall_out;

acl_pop local_bb4_notcmp41_pop43_c0_ene14_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_10_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene14_0_NO_SHIFT_REG),
	.stall_out(local_bb4_notcmp41_pop43_c0_ene14_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notcmp41_pop43_c0_ene14_fu_valid_out),
	.stall_in(local_bb4_notcmp41_pop43_c0_ene14_stall_local),
	.data_out(local_bb4_notcmp41_pop43_c0_ene14),
	.feedback_in(feedback_data_in_43),
	.feedback_valid_in(feedback_valid_in_43),
	.feedback_stall_out(feedback_stall_out_43)
);

defparam local_bb4_notcmp41_pop43_c0_ene14_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_notcmp41_pop43_c0_ene14_feedback.DATA_WIDTH = 1;
defparam local_bb4_notcmp41_pop43_c0_ene14_feedback.STYLE = "REGULAR";

assign local_bb4_notcmp41_pop43_c0_ene14_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_11_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_10_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene14_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notcmp41_pop43_c0_ene14_stall_local = 1'b0;
assign local_bb4_notcmp41_pop43_c0_ene14_valid_out_0 = 1'b1;
assign local_bb4_notcmp41_pop43_c0_ene14_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_11 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene14_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notexitcond943_pop44_c0_ene15_valid_out_0;
wire local_bb4_notexitcond943_pop44_c0_ene15_stall_in_0;
wire local_bb4_notexitcond943_pop44_c0_ene15_valid_out_1;
wire local_bb4_notexitcond943_pop44_c0_ene15_stall_in_1;
wire local_bb4_notexitcond943_pop44_c0_ene15_inputs_ready;
wire local_bb4_notexitcond943_pop44_c0_ene15_stall_local;
wire local_bb4_notexitcond943_pop44_c0_ene15;
wire local_bb4_notexitcond943_pop44_c0_ene15_fu_valid_out;
wire local_bb4_notexitcond943_pop44_c0_ene15_fu_stall_out;

acl_pop local_bb4_notexitcond943_pop44_c0_ene15_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_11_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene15_0_NO_SHIFT_REG),
	.stall_out(local_bb4_notexitcond943_pop44_c0_ene15_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond943_pop44_c0_ene15_fu_valid_out),
	.stall_in(local_bb4_notexitcond943_pop44_c0_ene15_stall_local),
	.data_out(local_bb4_notexitcond943_pop44_c0_ene15),
	.feedback_in(feedback_data_in_44),
	.feedback_valid_in(feedback_valid_in_44),
	.feedback_stall_out(feedback_stall_out_44)
);

defparam local_bb4_notexitcond943_pop44_c0_ene15_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_notexitcond943_pop44_c0_ene15_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond943_pop44_c0_ene15_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond943_pop44_c0_ene15_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_12_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_11_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene15_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notexitcond943_pop44_c0_ene15_stall_local = 1'b0;
assign local_bb4_notexitcond943_pop44_c0_ene15_valid_out_0 = 1'b1;
assign local_bb4_notexitcond943_pop44_c0_ene15_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_12 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_11_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene15_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__pop47_c0_ene16_valid_out_0;
wire local_bb4__pop47_c0_ene16_stall_in_0;
wire local_bb4__pop47_c0_ene16_valid_out_1;
wire local_bb4__pop47_c0_ene16_stall_in_1;
wire local_bb4__pop47_c0_ene16_inputs_ready;
wire local_bb4__pop47_c0_ene16_stall_local;
wire local_bb4__pop47_c0_ene16;
wire local_bb4__pop47_c0_ene16_fu_valid_out;
wire local_bb4__pop47_c0_ene16_fu_stall_out;

acl_pop local_bb4__pop47_c0_ene16_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene262_12_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene16_0_NO_SHIFT_REG),
	.stall_out(local_bb4__pop47_c0_ene16_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__pop47_c0_ene16_fu_valid_out),
	.stall_in(local_bb4__pop47_c0_ene16_stall_local),
	.data_out(local_bb4__pop47_c0_ene16),
	.feedback_in(feedback_data_in_47),
	.feedback_valid_in(feedback_valid_in_47),
	.feedback_stall_out(feedback_stall_out_47)
);

defparam local_bb4__pop47_c0_ene16_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4__pop47_c0_ene16_feedback.DATA_WIDTH = 1;
defparam local_bb4__pop47_c0_ene16_feedback.STYLE = "REGULAR";

assign local_bb4__pop47_c0_ene16_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_13_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene262_0_valid_out_12_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene16_0_valid_out_NO_SHIFT_REG);
assign local_bb4__pop47_c0_ene16_stall_local = 1'b0;
assign local_bb4__pop47_c0_ene16_valid_out_0 = 1'b1;
assign local_bb4__pop47_c0_ene16_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_13 = 1'b0;
assign rnode_9to10_bb4_c0_ene262_0_stall_in_12_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene16_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_keep_going_acl_pipeline_1_stall_in = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_NO_SHIFT_REG = rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i_i_valid_out;
wire local_bb4_cmp_i_i_stall_in;
wire local_bb4_cmp_i_i_inputs_ready;
wire local_bb4_cmp_i_i_stall_local;
wire local_bb4_cmp_i_i;

assign local_bb4_cmp_i_i_inputs_ready = rnode_7to8_bb4_add16_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_cmp_i_i = ($signed(rnode_7to8_bb4_add16_0_NO_SHIFT_REG) < $signed(32'h0));
assign local_bb4_cmp_i_i_valid_out = 1'b1;
assign rnode_7to8_bb4_add16_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp1_i_i_valid_out;
wire local_bb4_cmp1_i_i_stall_in;
wire local_bb4_cmp1_i_i_inputs_ready;
wire local_bb4_cmp1_i_i_stall_local;
wire local_bb4_cmp1_i_i;

assign local_bb4_cmp1_i_i_inputs_ready = rnode_7to8_bb4_add16_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp1_i_i = ($signed(rnode_7to8_bb4_add16_1_NO_SHIFT_REG) > $signed(input_wii_sub20));
assign local_bb4_cmp1_i_i_valid_out = 1'b1;
assign rnode_7to8_bb4_add16_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_add16_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add16_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_add16_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add16_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_add16_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add16_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add16_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add16_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_add16_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_add16_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_add16_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_add16_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_add16_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_7to8_bb4_add16_2_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_add16_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_add16_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_add16_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4_add16_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_add16_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_add16_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add16_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_add16_0_NO_SHIFT_REG = rnode_8to9_bb4_add16_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_add16_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_add16_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp14_valid_out;
wire local_bb4_cmp14_stall_in;
wire local_bb4_cmp14_inputs_ready;
wire local_bb4_cmp14_stall_local;
wire local_bb4_cmp14;

assign local_bb4_cmp14_inputs_ready = rnode_7to8_bb4_inc_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_cmp14 = ($signed(rnode_7to8_bb4_inc_0_NO_SHIFT_REG) > $signed(input_r));
assign local_bb4_cmp14_valid_out = 1'b1;
assign rnode_7to8_bb4_inc_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_inc_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_inc_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_inc_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_inc_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_inc_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_inc_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_inc_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_inc_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_inc_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_inc_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_inc_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_inc_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_inc_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_7to8_bb4_inc_1_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_inc_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_inc_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_inc_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4_inc_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_inc_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_inc_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_inc_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_inc_0_NO_SHIFT_REG = rnode_8to9_bb4_inc_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_inc_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_inc_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4__pop40_c0_ene363_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4__pop40_c0_ene363_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4__pop40_c0_ene363_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4__pop40_c0_ene363_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4__pop40_c0_ene363_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4__pop40_c0_ene363_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4__pop40_c0_ene363_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4__pop40_c0_ene363_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4__pop40_c0_ene363_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_7to8_bb4__pop40_c0_ene363_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4__pop40_c0_ene363_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4__pop40_c0_ene363_0_NO_SHIFT_REG = rnode_8to9_bb4__pop40_c0_ene363_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4__pop40_c0_ene363_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4__pop40_c0_ene363_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_forked1644_pop45_c0_ene161),
	.data_out(rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_forked1644_pop45_c0_ene161_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_NO_SHIFT_REG = rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_memdep_phi1_or39_pop41_c0_ene565),
	.data_out(rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_memdep_phi1_or39_pop41_c0_ene565_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_NO_SHIFT_REG = rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4__pop42_c0_ene666_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop42_c0_ene666_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4__pop42_c0_ene666_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop42_c0_ene666_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop42_c0_ene666_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop42_c0_ene666_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4__pop42_c0_ene666_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4__pop42_c0_ene666_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4__pop42_c0_ene666_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4__pop42_c0_ene666),
	.data_out(rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_fifo.DATA_WIDTH = 32;
defparam rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__pop42_c0_ene666_stall_in_1 = 1'b0;
assign rnode_10to11_bb4__pop42_c0_ene666_0_NO_SHIFT_REG = rnode_10to11_bb4__pop42_c0_ene666_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4__pop42_c0_ene666_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__pop42_c0_ene666_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_mul3724_pop34_c0_ene868),
	.data_out(rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_fifo.DATA_WIDTH = 32;
defparam rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_mul3724_pop34_c0_ene868_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_NO_SHIFT_REG = rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notcmp1127_pop35_c0_ene969),
	.data_out(rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notcmp1127_pop35_c0_ene969_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_NO_SHIFT_REG = rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond1430_pop36_c0_ene1070),
	.data_out(rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond1430_pop36_c0_ene1070_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_NO_SHIFT_REG = rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_indvars_iv_pop1037_pop39_c0_ene1373),
	.data_out(rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_NO_SHIFT_REG = rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notcmp41_pop43_c0_ene14),
	.data_out(rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notcmp41_pop43_c0_ene14_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_NO_SHIFT_REG = rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond943_pop44_c0_ene15),
	.data_out(rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond943_pop44_c0_ene15_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_NO_SHIFT_REG = rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4__pop47_c0_ene16_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop47_c0_ene16_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop47_c0_ene16_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop47_c0_ene16_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop47_c0_ene16_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop47_c0_ene16_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4__pop47_c0_ene16_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4__pop47_c0_ene16_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4__pop47_c0_ene16_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4__pop47_c0_ene16),
	.data_out(rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__pop47_c0_ene16_stall_in_1 = 1'b0;
assign rnode_10to11_bb4__pop47_c0_ene16_0_NO_SHIFT_REG = rnode_10to11_bb4__pop47_c0_ene16_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4__pop47_c0_ene16_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__pop47_c0_ene16_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_cmp_i_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp_i_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp_i_i_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp_i_i_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp_i_i_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp_i_i_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp_i_i_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp_i_i_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_cmp_i_i_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_cmp_i_i_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_cmp_i_i_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_cmp_i_i_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_cmp_i_i_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(local_bb4_cmp_i_i),
	.data_out(rnode_8to9_bb4_cmp_i_i_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_cmp_i_i_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_cmp_i_i_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_cmp_i_i_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_cmp_i_i_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_cmp_i_i_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp_i_i_stall_in = 1'b0;
assign rnode_8to9_bb4_cmp_i_i_0_NO_SHIFT_REG = rnode_8to9_bb4_cmp_i_i_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_cmp_i_i_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_cmp_i_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_cmp1_i_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp1_i_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp1_i_i_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp1_i_i_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp1_i_i_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp1_i_i_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp1_i_i_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp1_i_i_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_cmp1_i_i_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_cmp1_i_i_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_cmp1_i_i_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_cmp1_i_i_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_cmp1_i_i_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(local_bb4_cmp1_i_i),
	.data_out(rnode_8to9_bb4_cmp1_i_i_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_cmp1_i_i_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_cmp1_i_i_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_cmp1_i_i_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_cmp1_i_i_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_cmp1_i_i_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp1_i_i_stall_in = 1'b0;
assign rnode_8to9_bb4_cmp1_i_i_0_NO_SHIFT_REG = rnode_8to9_bb4_cmp1_i_i_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_cmp1_i_i_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_cmp1_i_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_cmp14_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_cmp14_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_cmp14_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_cmp14_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_cmp14_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_cmp14_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_cmp14_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(local_bb4_cmp14),
	.data_out(rnode_8to9_bb4_cmp14_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_cmp14_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_cmp14_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp14_stall_in = 1'b0;
assign rnode_8to9_bb4_cmp14_0_NO_SHIFT_REG = rnode_8to9_bb4_cmp14_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_cmp14_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_cmp14_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4__pop40_c0_ene363_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4__pop40_c0_ene363_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4__pop40_c0_ene363_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4__pop40_c0_ene363_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4__pop40_c0_ene363_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4__pop40_c0_ene363_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4__pop40_c0_ene363_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4__pop40_c0_ene363_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4__pop40_c0_ene363_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_8to9_bb4__pop40_c0_ene363_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4__pop40_c0_ene363_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4__pop40_c0_ene363_0_NO_SHIFT_REG = rnode_9to10_bb4__pop40_c0_ene363_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4__pop40_c0_ene363_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4__pop40_c0_ene363_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi174_stall_local;
wire [447:0] local_bb4_c0_exi174;

assign local_bb4_c0_exi174[7:0] = 8'bx;
assign local_bb4_c0_exi174[8] = rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_NO_SHIFT_REG;
assign local_bb4_c0_exi174[447:9] = 439'bx;

// This section implements an unregistered operation.
// 
wire local_bb4___stall_local;
wire [31:0] local_bb4__;

assign local_bb4__ = (rnode_8to9_bb4_cmp1_i_i_0_NO_SHIFT_REG ? input_wii_sub20 : rnode_8to9_bb4_add16_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__stall_local;
wire local_bb4_var_;

assign local_bb4_var_ = (input_wii_var__u17 | rnode_8to9_bb4_cmp14_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4___u23_stall_local;
wire [31:0] local_bb4___u23;

assign local_bb4___u23 = (rnode_8to9_bb4_cmp_i_i_0_NO_SHIFT_REG ? 32'h0 : local_bb4__);

// This section implements an unregistered operation.
// 
wire local_bb4_var__valid_out_1;
wire local_bb4_var__stall_in_1;
wire local_bb4_notexit_valid_out_0;
wire local_bb4_notexit_stall_in_0;
wire local_bb4_notexit_valid_out_1;
wire local_bb4_notexit_stall_in_1;
wire local_bb4_notexit_inputs_ready;
wire local_bb4_notexit_stall_local;
wire local_bb4_notexit;

assign local_bb4_notexit_inputs_ready = rnode_8to9_bb4_cmp14_0_valid_out_NO_SHIFT_REG;
assign local_bb4_notexit = (local_bb4_var_ ^ 1'b1);
assign local_bb4_var__valid_out_1 = 1'b1;
assign local_bb4_notexit_valid_out_0 = 1'b1;
assign local_bb4_notexit_valid_out_1 = 1'b1;
assign rnode_8to9_bb4_cmp14_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_mul2445_pop46_c0_ene464_valid_out_1;
wire local_bb4_mul2445_pop46_c0_ene464_stall_in_1;
wire local_bb4_add25_valid_out;
wire local_bb4_add25_stall_in;
wire local_bb4_add25_inputs_ready;
wire local_bb4_add25_stall_local;
wire [31:0] local_bb4_add25;

assign local_bb4_add25_inputs_ready = (SFC_2_VALID_8_9_0_valid_out_2_NO_SHIFT_REG & rnode_7to9_bb4_c0_ene262_0_valid_out_0_NO_SHIFT_REG & rnode_8to9_bb4_c0_ene464_0_valid_out_NO_SHIFT_REG & rnode_8to9_bb4_cmp1_i_i_0_valid_out_NO_SHIFT_REG & rnode_8to9_bb4_add16_0_valid_out_NO_SHIFT_REG & rnode_8to9_bb4_cmp_i_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_add25 = (local_bb4_mul2445_pop46_c0_ene464 + local_bb4___u23);
assign local_bb4_mul2445_pop46_c0_ene464_valid_out_1 = 1'b1;
assign local_bb4_add25_valid_out = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in_2 = 1'b0;
assign rnode_7to9_bb4_c0_ene262_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene464_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_cmp1_i_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_add16_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_cmp_i_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_9to11_bb4_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__0_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__0_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_var__0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_9to11_bb4_var__0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to11_bb4_var__0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to11_bb4_var__0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_9to11_bb4_var__0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_9to11_bb4_var__0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_var_),
	.data_out(rnode_9to11_bb4_var__0_reg_11_NO_SHIFT_REG)
);

defparam rnode_9to11_bb4_var__0_reg_11_fifo.DEPTH = 2;
defparam rnode_9to11_bb4_var__0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_9to11_bb4_var__0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to11_bb4_var__0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_9to11_bb4_var__0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__stall_in_1 = 1'b0;
assign rnode_9to11_bb4_var__0_NO_SHIFT_REG = rnode_9to11_bb4_var__0_reg_11_NO_SHIFT_REG;
assign rnode_9to11_bb4_var__0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_var__0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_notexitcond_notexit_inputs_ready;
 reg local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_0;
 reg local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_1;
 reg local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_2;
 reg local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_3;
 reg local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_4;
 reg local_bb4_notexitcond_notexit_valid_out_5_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_5;
 reg local_bb4_notexitcond_notexit_valid_out_6_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_6;
 reg local_bb4_notexitcond_notexit_valid_out_7_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_7;
 reg local_bb4_notexitcond_notexit_valid_out_8_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_8;
 reg local_bb4_notexitcond_notexit_valid_out_9_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_9;
 reg local_bb4_notexitcond_notexit_valid_out_10_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_10;
 reg local_bb4_notexitcond_notexit_valid_out_11_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_11;
 reg local_bb4_notexitcond_notexit_valid_out_12_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_12;
 reg local_bb4_notexitcond_notexit_valid_out_13_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_13;
 reg local_bb4_notexitcond_notexit_valid_out_14_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_14;
 reg local_bb4_notexitcond_notexit_valid_out_15_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_15;
wire local_bb4_notexitcond_notexit_output_regs_ready;
wire local_bb4_notexitcond_notexit_result;
wire local_bb4_notexitcond_notexit_fu_valid_out;
wire local_bb4_notexitcond_notexit_fu_stall_out;
 reg local_bb4_notexitcond_notexit_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_causedstall;

acl_push local_bb4_notexitcond_notexit_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(local_bb4_notexit),
	.stall_out(local_bb4_notexitcond_notexit_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond_notexit_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond_notexit_result),
	.feedback_out(feedback_data_out_1),
	.feedback_valid_out(feedback_valid_out_1),
	.feedback_stall_in(feedback_stall_in_1)
);

defparam local_bb4_notexitcond_notexit_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond_notexit_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond_notexit_feedback.FIFO_DEPTH = 8;
defparam local_bb4_notexitcond_notexit_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_notexitcond_notexit_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond_notexit_inputs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_output_regs_ready = 1'b1;
assign local_bb4_notexit_stall_in_0 = 1'b0;
assign SFC_2_VALID_8_9_0_stall_in_3 = 1'b0;
assign local_bb4_notexitcond_notexit_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond_notexit_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_7_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_8_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_9_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_10_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_11_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_12_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_13_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_14_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_15_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond_notexit_output_regs_ready)
		begin
			local_bb4_notexitcond_notexit_NO_SHIFT_REG <= local_bb4_notexitcond_notexit_result;
			local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_6_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_7_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_8_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_9_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_10_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_11_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_12_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_13_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_14_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_15_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond_notexit_stall_in_0))
			begin
				local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_1))
			begin
				local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_2))
			begin
				local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_3))
			begin
				local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_4))
			begin
				local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_5))
			begin
				local_bb4_notexitcond_notexit_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_6))
			begin
				local_bb4_notexitcond_notexit_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_7))
			begin
				local_bb4_notexitcond_notexit_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_8))
			begin
				local_bb4_notexitcond_notexit_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_9))
			begin
				local_bb4_notexitcond_notexit_valid_out_9_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_10))
			begin
				local_bb4_notexitcond_notexit_valid_out_10_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_11))
			begin
				local_bb4_notexitcond_notexit_valid_out_11_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_12))
			begin
				local_bb4_notexitcond_notexit_valid_out_12_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_13))
			begin
				local_bb4_notexitcond_notexit_valid_out_13_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_14))
			begin
				local_bb4_notexitcond_notexit_valid_out_14_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_15))
			begin
				local_bb4_notexitcond_notexit_valid_out_15_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_j_35_push30_inc_inputs_ready;
 reg local_bb4_j_35_push30_inc_valid_out_NO_SHIFT_REG;
wire local_bb4_j_35_push30_inc_stall_in;
wire local_bb4_j_35_push30_inc_output_regs_ready;
wire [31:0] local_bb4_j_35_push30_inc_result;
wire local_bb4_j_35_push30_inc_fu_valid_out;
wire local_bb4_j_35_push30_inc_fu_stall_out;
 reg [31:0] local_bb4_j_35_push30_inc_NO_SHIFT_REG;
wire local_bb4_j_35_push30_inc_causedstall;

acl_push local_bb4_j_35_push30_inc_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexit),
	.predicate(1'b0),
	.data_in(rnode_8to9_bb4_inc_0_NO_SHIFT_REG),
	.stall_out(local_bb4_j_35_push30_inc_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_j_35_push30_inc_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_j_35_push30_inc_result),
	.feedback_out(feedback_data_out_30),
	.feedback_valid_out(feedback_valid_out_30),
	.feedback_stall_in(feedback_stall_in_30)
);

defparam local_bb4_j_35_push30_inc_feedback.STALLFREE = 1;
defparam local_bb4_j_35_push30_inc_feedback.DATA_WIDTH = 32;
defparam local_bb4_j_35_push30_inc_feedback.FIFO_DEPTH = 9;
defparam local_bb4_j_35_push30_inc_feedback.MIN_FIFO_LATENCY = 7;
defparam local_bb4_j_35_push30_inc_feedback.STYLE = "REGULAR";

assign local_bb4_j_35_push30_inc_inputs_ready = 1'b1;
assign local_bb4_j_35_push30_inc_output_regs_ready = 1'b1;
assign local_bb4_notexit_stall_in_1 = 1'b0;
assign SFC_2_VALID_8_9_0_stall_in_4 = 1'b0;
assign rnode_8to9_bb4_inc_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_j_35_push30_inc_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_j_35_push30_inc_NO_SHIFT_REG <= 'x;
		local_bb4_j_35_push30_inc_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_j_35_push30_inc_output_regs_ready)
		begin
			local_bb4_j_35_push30_inc_NO_SHIFT_REG <= local_bb4_j_35_push30_inc_result;
			local_bb4_j_35_push30_inc_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_j_35_push30_inc_stall_in))
			begin
				local_bb4_j_35_push30_inc_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(local_bb4_mul2445_pop46_c0_ene464),
	.data_out(rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_mul2445_pop46_c0_ene464_stall_in_1 = 1'b0;
assign rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_NO_SHIFT_REG = rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_add25_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_add25_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add25_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_add25_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add25_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add25_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add25_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_add25_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_add25_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_add25_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_add25_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_add25_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(local_bb4_add25),
	.data_out(rnode_9to10_bb4_add25_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_add25_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_add25_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_add25_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_add25_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_add25_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add25_stall_in = 1'b0;
assign rnode_9to10_bb4_add25_0_NO_SHIFT_REG = rnode_9to10_bb4_add25_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_add25_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_add25_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_forked1644_push45_forked1644_pop45_inputs_ready;
 reg local_bb4_forked1644_push45_forked1644_pop45_valid_out_NO_SHIFT_REG;
wire local_bb4_forked1644_push45_forked1644_pop45_stall_in;
wire local_bb4_forked1644_push45_forked1644_pop45_output_regs_ready;
wire local_bb4_forked1644_push45_forked1644_pop45_result;
wire local_bb4_forked1644_push45_forked1644_pop45_fu_valid_out;
wire local_bb4_forked1644_push45_forked1644_pop45_fu_stall_out;
 reg local_bb4_forked1644_push45_forked1644_pop45_NO_SHIFT_REG;
wire local_bb4_forked1644_push45_forked1644_pop45_causedstall;

acl_push local_bb4_forked1644_push45_forked1644_pop45_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_forked1644_pop45_c0_ene161),
	.stall_out(local_bb4_forked1644_push45_forked1644_pop45_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_forked1644_push45_forked1644_pop45_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_forked1644_push45_forked1644_pop45_result),
	.feedback_out(feedback_data_out_45),
	.feedback_valid_out(feedback_valid_out_45),
	.feedback_stall_in(feedback_stall_in_45)
);

defparam local_bb4_forked1644_push45_forked1644_pop45_feedback.STALLFREE = 1;
defparam local_bb4_forked1644_push45_forked1644_pop45_feedback.DATA_WIDTH = 1;
defparam local_bb4_forked1644_push45_forked1644_pop45_feedback.FIFO_DEPTH = 9;
defparam local_bb4_forked1644_push45_forked1644_pop45_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_forked1644_push45_forked1644_pop45_feedback.STYLE = "REGULAR";

assign local_bb4_forked1644_push45_forked1644_pop45_inputs_ready = 1'b1;
assign local_bb4_forked1644_push45_forked1644_pop45_output_regs_ready = 1'b1;
assign local_bb4_forked1644_pop45_c0_ene161_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_1 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_15 = 1'b0;
assign local_bb4_forked1644_push45_forked1644_pop45_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_forked1644_push45_forked1644_pop45_NO_SHIFT_REG <= 'x;
		local_bb4_forked1644_push45_forked1644_pop45_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_forked1644_push45_forked1644_pop45_output_regs_ready)
		begin
			local_bb4_forked1644_push45_forked1644_pop45_NO_SHIFT_REG <= local_bb4_forked1644_push45_forked1644_pop45_result;
			local_bb4_forked1644_push45_forked1644_pop45_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_forked1644_push45_forked1644_pop45_stall_in))
			begin
				local_bb4_forked1644_push45_forked1644_pop45_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4__push42__pop42_inputs_ready;
 reg local_bb4__push42__pop42_valid_out_NO_SHIFT_REG;
wire local_bb4__push42__pop42_stall_in;
wire local_bb4__push42__pop42_output_regs_ready;
wire [31:0] local_bb4__push42__pop42_result;
wire local_bb4__push42__pop42_fu_valid_out;
wire local_bb4__push42__pop42_fu_stall_out;
 reg [31:0] local_bb4__push42__pop42_NO_SHIFT_REG;
wire local_bb4__push42__pop42_causedstall;

acl_push local_bb4__push42__pop42_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4__pop42_c0_ene666),
	.stall_out(local_bb4__push42__pop42_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__push42__pop42_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4__push42__pop42_result),
	.feedback_out(feedback_data_out_42),
	.feedback_valid_out(feedback_valid_out_42),
	.feedback_stall_in(feedback_stall_in_42)
);

defparam local_bb4__push42__pop42_feedback.STALLFREE = 1;
defparam local_bb4__push42__pop42_feedback.DATA_WIDTH = 32;
defparam local_bb4__push42__pop42_feedback.FIFO_DEPTH = 9;
defparam local_bb4__push42__pop42_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4__push42__pop42_feedback.STYLE = "REGULAR";

assign local_bb4__push42__pop42_inputs_ready = 1'b1;
assign local_bb4__push42__pop42_output_regs_ready = 1'b1;
assign local_bb4__pop42_c0_ene666_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_2 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_16 = 1'b0;
assign local_bb4__push42__pop42_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4__push42__pop42_NO_SHIFT_REG <= 'x;
		local_bb4__push42__pop42_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4__push42__pop42_output_regs_ready)
		begin
			local_bb4__push42__pop42_NO_SHIFT_REG <= local_bb4__push42__pop42_result;
			local_bb4__push42__pop42_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4__push42__pop42_stall_in))
			begin
				local_bb4__push42__pop42_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_inputs_ready;
 reg local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_valid_out_NO_SHIFT_REG;
wire local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_stall_in;
wire local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_output_regs_ready;
wire local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_result;
wire local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_fu_valid_out;
wire local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_fu_stall_out;
 reg local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_NO_SHIFT_REG;
wire local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_causedstall;

acl_push local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_memdep_phi1_or39_pop41_c0_ene565),
	.stall_out(local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_result),
	.feedback_out(feedback_data_out_41),
	.feedback_valid_out(feedback_valid_out_41),
	.feedback_stall_in(feedback_stall_in_41)
);

defparam local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_feedback.STALLFREE = 1;
defparam local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_feedback.DATA_WIDTH = 1;
defparam local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_feedback.FIFO_DEPTH = 9;
defparam local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_feedback.STYLE = "REGULAR";

assign local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_inputs_ready = 1'b1;
assign local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_output_regs_ready = 1'b1;
assign local_bb4_memdep_phi1_or39_pop41_c0_ene565_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_3 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_17 = 1'b0;
assign local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_NO_SHIFT_REG <= 'x;
		local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_output_regs_ready)
		begin
			local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_NO_SHIFT_REG <= local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_result;
			local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_stall_in))
			begin
				local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4__push40__pop40_inputs_ready;
 reg local_bb4__push40__pop40_valid_out_NO_SHIFT_REG;
wire local_bb4__push40__pop40_stall_in;
wire local_bb4__push40__pop40_output_regs_ready;
wire [31:0] local_bb4__push40__pop40_result;
wire local_bb4__push40__pop40_fu_valid_out;
wire local_bb4__push40__pop40_fu_stall_out;
 reg [31:0] local_bb4__push40__pop40_NO_SHIFT_REG;
wire local_bb4__push40__pop40_causedstall;

acl_push local_bb4__push40__pop40_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4__pop40_c0_ene363_0_NO_SHIFT_REG),
	.stall_out(local_bb4__push40__pop40_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__push40__pop40_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4__push40__pop40_result),
	.feedback_out(feedback_data_out_40),
	.feedback_valid_out(feedback_valid_out_40),
	.feedback_stall_in(feedback_stall_in_40)
);

defparam local_bb4__push40__pop40_feedback.STALLFREE = 1;
defparam local_bb4__push40__pop40_feedback.DATA_WIDTH = 32;
defparam local_bb4__push40__pop40_feedback.FIFO_DEPTH = 9;
defparam local_bb4__push40__pop40_feedback.MIN_FIFO_LATENCY = 6;
defparam local_bb4__push40__pop40_feedback.STYLE = "REGULAR";

assign local_bb4__push40__pop40_inputs_ready = 1'b1;
assign local_bb4__push40__pop40_output_regs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_4 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_18 = 1'b0;
assign rnode_9to10_bb4__pop40_c0_ene363_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4__push40__pop40_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4__push40__pop40_NO_SHIFT_REG <= 'x;
		local_bb4__push40__pop40_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4__push40__pop40_output_regs_ready)
		begin
			local_bb4__push40__pop40_NO_SHIFT_REG <= local_bb4__push40__pop40_result;
			local_bb4__push40__pop40_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4__push40__pop40_stall_in))
			begin
				local_bb4__push40__pop40_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_inputs_ready;
 reg local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_valid_out_NO_SHIFT_REG;
wire local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_stall_in;
wire local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_output_regs_ready;
wire [31:0] local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_result;
wire local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_fu_valid_out;
wire local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_fu_stall_out;
 reg [31:0] local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_NO_SHIFT_REG;
wire local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_causedstall;

acl_push local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_pixel_y_020_pop821_pop33_c0_ene767),
	.stall_out(local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_result),
	.feedback_out(feedback_data_out_33),
	.feedback_valid_out(feedback_valid_out_33),
	.feedback_stall_in(feedback_stall_in_33)
);

defparam local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_feedback.STALLFREE = 1;
defparam local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_feedback.DATA_WIDTH = 32;
defparam local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_feedback.FIFO_DEPTH = 9;
defparam local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_feedback.STYLE = "REGULAR";

assign local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_inputs_ready = 1'b1;
assign local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_output_regs_ready = 1'b1;
assign local_bb4_pixel_y_020_pop821_pop33_c0_ene767_stall_in = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_5 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_19 = 1'b0;
assign local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_NO_SHIFT_REG <= 'x;
		local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_output_regs_ready)
		begin
			local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_NO_SHIFT_REG <= local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_result;
			local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_stall_in))
			begin
				local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_mul3724_push34_mul3724_pop34_inputs_ready;
 reg local_bb4_mul3724_push34_mul3724_pop34_valid_out_NO_SHIFT_REG;
wire local_bb4_mul3724_push34_mul3724_pop34_stall_in;
wire local_bb4_mul3724_push34_mul3724_pop34_output_regs_ready;
wire [31:0] local_bb4_mul3724_push34_mul3724_pop34_result;
wire local_bb4_mul3724_push34_mul3724_pop34_fu_valid_out;
wire local_bb4_mul3724_push34_mul3724_pop34_fu_stall_out;
 reg [31:0] local_bb4_mul3724_push34_mul3724_pop34_NO_SHIFT_REG;
wire local_bb4_mul3724_push34_mul3724_pop34_causedstall;

acl_push local_bb4_mul3724_push34_mul3724_pop34_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_mul3724_pop34_c0_ene868),
	.stall_out(local_bb4_mul3724_push34_mul3724_pop34_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_mul3724_push34_mul3724_pop34_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_mul3724_push34_mul3724_pop34_result),
	.feedback_out(feedback_data_out_34),
	.feedback_valid_out(feedback_valid_out_34),
	.feedback_stall_in(feedback_stall_in_34)
);

defparam local_bb4_mul3724_push34_mul3724_pop34_feedback.STALLFREE = 1;
defparam local_bb4_mul3724_push34_mul3724_pop34_feedback.DATA_WIDTH = 32;
defparam local_bb4_mul3724_push34_mul3724_pop34_feedback.FIFO_DEPTH = 9;
defparam local_bb4_mul3724_push34_mul3724_pop34_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_mul3724_push34_mul3724_pop34_feedback.STYLE = "REGULAR";

assign local_bb4_mul3724_push34_mul3724_pop34_inputs_ready = 1'b1;
assign local_bb4_mul3724_push34_mul3724_pop34_output_regs_ready = 1'b1;
assign local_bb4_mul3724_pop34_c0_ene868_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_6 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_20 = 1'b0;
assign local_bb4_mul3724_push34_mul3724_pop34_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul3724_push34_mul3724_pop34_NO_SHIFT_REG <= 'x;
		local_bb4_mul3724_push34_mul3724_pop34_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul3724_push34_mul3724_pop34_output_regs_ready)
		begin
			local_bb4_mul3724_push34_mul3724_pop34_NO_SHIFT_REG <= local_bb4_mul3724_push34_mul3724_pop34_result;
			local_bb4_mul3724_push34_mul3724_pop34_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul3724_push34_mul3724_pop34_stall_in))
			begin
				local_bb4_mul3724_push34_mul3724_pop34_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_notcmp1127_push35_notcmp1127_pop35_inputs_ready;
 reg local_bb4_notcmp1127_push35_notcmp1127_pop35_valid_out_NO_SHIFT_REG;
wire local_bb4_notcmp1127_push35_notcmp1127_pop35_stall_in;
wire local_bb4_notcmp1127_push35_notcmp1127_pop35_output_regs_ready;
wire local_bb4_notcmp1127_push35_notcmp1127_pop35_result;
wire local_bb4_notcmp1127_push35_notcmp1127_pop35_fu_valid_out;
wire local_bb4_notcmp1127_push35_notcmp1127_pop35_fu_stall_out;
 reg local_bb4_notcmp1127_push35_notcmp1127_pop35_NO_SHIFT_REG;
wire local_bb4_notcmp1127_push35_notcmp1127_pop35_causedstall;

acl_push local_bb4_notcmp1127_push35_notcmp1127_pop35_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_notcmp1127_pop35_c0_ene969),
	.stall_out(local_bb4_notcmp1127_push35_notcmp1127_pop35_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notcmp1127_push35_notcmp1127_pop35_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notcmp1127_push35_notcmp1127_pop35_result),
	.feedback_out(feedback_data_out_35),
	.feedback_valid_out(feedback_valid_out_35),
	.feedback_stall_in(feedback_stall_in_35)
);

defparam local_bb4_notcmp1127_push35_notcmp1127_pop35_feedback.STALLFREE = 1;
defparam local_bb4_notcmp1127_push35_notcmp1127_pop35_feedback.DATA_WIDTH = 1;
defparam local_bb4_notcmp1127_push35_notcmp1127_pop35_feedback.FIFO_DEPTH = 9;
defparam local_bb4_notcmp1127_push35_notcmp1127_pop35_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_notcmp1127_push35_notcmp1127_pop35_feedback.STYLE = "REGULAR";

assign local_bb4_notcmp1127_push35_notcmp1127_pop35_inputs_ready = 1'b1;
assign local_bb4_notcmp1127_push35_notcmp1127_pop35_output_regs_ready = 1'b1;
assign local_bb4_notcmp1127_pop35_c0_ene969_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_7 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_21 = 1'b0;
assign local_bb4_notcmp1127_push35_notcmp1127_pop35_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notcmp1127_push35_notcmp1127_pop35_NO_SHIFT_REG <= 'x;
		local_bb4_notcmp1127_push35_notcmp1127_pop35_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notcmp1127_push35_notcmp1127_pop35_output_regs_ready)
		begin
			local_bb4_notcmp1127_push35_notcmp1127_pop35_NO_SHIFT_REG <= local_bb4_notcmp1127_push35_notcmp1127_pop35_result;
			local_bb4_notcmp1127_push35_notcmp1127_pop35_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notcmp1127_push35_notcmp1127_pop35_stall_in))
			begin
				local_bb4_notcmp1127_push35_notcmp1127_pop35_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_notexitcond1430_push36_notexitcond1430_pop36_inputs_ready;
 reg local_bb4_notexitcond1430_push36_notexitcond1430_pop36_valid_out_NO_SHIFT_REG;
wire local_bb4_notexitcond1430_push36_notexitcond1430_pop36_stall_in;
wire local_bb4_notexitcond1430_push36_notexitcond1430_pop36_output_regs_ready;
wire local_bb4_notexitcond1430_push36_notexitcond1430_pop36_result;
wire local_bb4_notexitcond1430_push36_notexitcond1430_pop36_fu_valid_out;
wire local_bb4_notexitcond1430_push36_notexitcond1430_pop36_fu_stall_out;
 reg local_bb4_notexitcond1430_push36_notexitcond1430_pop36_NO_SHIFT_REG;
wire local_bb4_notexitcond1430_push36_notexitcond1430_pop36_causedstall;

acl_push local_bb4_notexitcond1430_push36_notexitcond1430_pop36_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_notexitcond1430_pop36_c0_ene1070),
	.stall_out(local_bb4_notexitcond1430_push36_notexitcond1430_pop36_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond1430_push36_notexitcond1430_pop36_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond1430_push36_notexitcond1430_pop36_result),
	.feedback_out(feedback_data_out_36),
	.feedback_valid_out(feedback_valid_out_36),
	.feedback_stall_in(feedback_stall_in_36)
);

defparam local_bb4_notexitcond1430_push36_notexitcond1430_pop36_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond1430_push36_notexitcond1430_pop36_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond1430_push36_notexitcond1430_pop36_feedback.FIFO_DEPTH = 9;
defparam local_bb4_notexitcond1430_push36_notexitcond1430_pop36_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_notexitcond1430_push36_notexitcond1430_pop36_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond1430_push36_notexitcond1430_pop36_inputs_ready = 1'b1;
assign local_bb4_notexitcond1430_push36_notexitcond1430_pop36_output_regs_ready = 1'b1;
assign local_bb4_notexitcond1430_pop36_c0_ene1070_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_8 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_22 = 1'b0;
assign local_bb4_notexitcond1430_push36_notexitcond1430_pop36_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond1430_push36_notexitcond1430_pop36_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond1430_push36_notexitcond1430_pop36_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond1430_push36_notexitcond1430_pop36_output_regs_ready)
		begin
			local_bb4_notexitcond1430_push36_notexitcond1430_pop36_NO_SHIFT_REG <= local_bb4_notexitcond1430_push36_notexitcond1430_pop36_result;
			local_bb4_notexitcond1430_push36_notexitcond1430_pop36_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond1430_push36_notexitcond1430_pop36_stall_in))
			begin
				local_bb4_notexitcond1430_push36_notexitcond1430_pop36_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_inputs_ready;
 reg local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_valid_out_NO_SHIFT_REG;
wire local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_stall_in;
wire local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_output_regs_ready;
wire local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_result;
wire local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_fu_valid_out;
wire local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_fu_stall_out;
 reg local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_NO_SHIFT_REG;
wire local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_causedstall;

acl_push local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_memdep_phi1_pop933_pop37_c0_ene1171),
	.stall_out(local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_result),
	.feedback_out(feedback_data_out_37),
	.feedback_valid_out(feedback_valid_out_37),
	.feedback_stall_in(feedback_stall_in_37)
);

defparam local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_feedback.STALLFREE = 1;
defparam local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_feedback.DATA_WIDTH = 1;
defparam local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_feedback.FIFO_DEPTH = 9;
defparam local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_feedback.STYLE = "REGULAR";

assign local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_inputs_ready = 1'b1;
assign local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_output_regs_ready = 1'b1;
assign local_bb4_memdep_phi1_pop933_pop37_c0_ene1171_stall_in = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_9 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_23 = 1'b0;
assign local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_NO_SHIFT_REG <= 'x;
		local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_output_regs_ready)
		begin
			local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_NO_SHIFT_REG <= local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_result;
			local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_stall_in))
			begin
				local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_mul535_push38_mul535_pop38_inputs_ready;
 reg local_bb4_mul535_push38_mul535_pop38_valid_out_NO_SHIFT_REG;
wire local_bb4_mul535_push38_mul535_pop38_stall_in;
wire local_bb4_mul535_push38_mul535_pop38_output_regs_ready;
wire [31:0] local_bb4_mul535_push38_mul535_pop38_result;
wire local_bb4_mul535_push38_mul535_pop38_fu_valid_out;
wire local_bb4_mul535_push38_mul535_pop38_fu_stall_out;
 reg [31:0] local_bb4_mul535_push38_mul535_pop38_NO_SHIFT_REG;
wire local_bb4_mul535_push38_mul535_pop38_causedstall;

acl_push local_bb4_mul535_push38_mul535_pop38_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_mul535_pop38_c0_ene1272),
	.stall_out(local_bb4_mul535_push38_mul535_pop38_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_mul535_push38_mul535_pop38_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_mul535_push38_mul535_pop38_result),
	.feedback_out(feedback_data_out_38),
	.feedback_valid_out(feedback_valid_out_38),
	.feedback_stall_in(feedback_stall_in_38)
);

defparam local_bb4_mul535_push38_mul535_pop38_feedback.STALLFREE = 1;
defparam local_bb4_mul535_push38_mul535_pop38_feedback.DATA_WIDTH = 32;
defparam local_bb4_mul535_push38_mul535_pop38_feedback.FIFO_DEPTH = 9;
defparam local_bb4_mul535_push38_mul535_pop38_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_mul535_push38_mul535_pop38_feedback.STYLE = "REGULAR";

assign local_bb4_mul535_push38_mul535_pop38_inputs_ready = 1'b1;
assign local_bb4_mul535_push38_mul535_pop38_output_regs_ready = 1'b1;
assign local_bb4_mul535_pop38_c0_ene1272_stall_in = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_10 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_24 = 1'b0;
assign local_bb4_mul535_push38_mul535_pop38_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul535_push38_mul535_pop38_NO_SHIFT_REG <= 'x;
		local_bb4_mul535_push38_mul535_pop38_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul535_push38_mul535_pop38_output_regs_ready)
		begin
			local_bb4_mul535_push38_mul535_pop38_NO_SHIFT_REG <= local_bb4_mul535_push38_mul535_pop38_result;
			local_bb4_mul535_push38_mul535_pop38_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul535_push38_mul535_pop38_stall_in))
			begin
				local_bb4_mul535_push38_mul535_pop38_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_inputs_ready;
 reg local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_valid_out_NO_SHIFT_REG;
wire local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_stall_in;
wire local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_output_regs_ready;
wire [63:0] local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_result;
wire local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_fu_valid_out;
wire local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_fu_stall_out;
 reg [63:0] local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_NO_SHIFT_REG;
wire local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_causedstall;

acl_push local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_indvars_iv_pop1037_pop39_c0_ene1373),
	.stall_out(local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_result),
	.feedback_out(feedback_data_out_39),
	.feedback_valid_out(feedback_valid_out_39),
	.feedback_stall_in(feedback_stall_in_39)
);

defparam local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_feedback.STALLFREE = 1;
defparam local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_feedback.DATA_WIDTH = 64;
defparam local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_feedback.FIFO_DEPTH = 9;
defparam local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_feedback.STYLE = "REGULAR";

assign local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_inputs_ready = 1'b1;
assign local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_output_regs_ready = 1'b1;
assign local_bb4_indvars_iv_pop1037_pop39_c0_ene1373_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_11 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_25 = 1'b0;
assign local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_NO_SHIFT_REG <= 'x;
		local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_output_regs_ready)
		begin
			local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_NO_SHIFT_REG <= local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_result;
			local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_stall_in))
			begin
				local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_notcmp41_push43_notcmp41_pop43_inputs_ready;
 reg local_bb4_notcmp41_push43_notcmp41_pop43_valid_out_NO_SHIFT_REG;
wire local_bb4_notcmp41_push43_notcmp41_pop43_stall_in;
wire local_bb4_notcmp41_push43_notcmp41_pop43_output_regs_ready;
wire local_bb4_notcmp41_push43_notcmp41_pop43_result;
wire local_bb4_notcmp41_push43_notcmp41_pop43_fu_valid_out;
wire local_bb4_notcmp41_push43_notcmp41_pop43_fu_stall_out;
 reg local_bb4_notcmp41_push43_notcmp41_pop43_NO_SHIFT_REG;
wire local_bb4_notcmp41_push43_notcmp41_pop43_causedstall;

acl_push local_bb4_notcmp41_push43_notcmp41_pop43_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_notcmp41_pop43_c0_ene14),
	.stall_out(local_bb4_notcmp41_push43_notcmp41_pop43_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notcmp41_push43_notcmp41_pop43_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notcmp41_push43_notcmp41_pop43_result),
	.feedback_out(feedback_data_out_43),
	.feedback_valid_out(feedback_valid_out_43),
	.feedback_stall_in(feedback_stall_in_43)
);

defparam local_bb4_notcmp41_push43_notcmp41_pop43_feedback.STALLFREE = 1;
defparam local_bb4_notcmp41_push43_notcmp41_pop43_feedback.DATA_WIDTH = 1;
defparam local_bb4_notcmp41_push43_notcmp41_pop43_feedback.FIFO_DEPTH = 9;
defparam local_bb4_notcmp41_push43_notcmp41_pop43_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_notcmp41_push43_notcmp41_pop43_feedback.STYLE = "REGULAR";

assign local_bb4_notcmp41_push43_notcmp41_pop43_inputs_ready = 1'b1;
assign local_bb4_notcmp41_push43_notcmp41_pop43_output_regs_ready = 1'b1;
assign local_bb4_notcmp41_pop43_c0_ene14_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_12 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_26 = 1'b0;
assign local_bb4_notcmp41_push43_notcmp41_pop43_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notcmp41_push43_notcmp41_pop43_NO_SHIFT_REG <= 'x;
		local_bb4_notcmp41_push43_notcmp41_pop43_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notcmp41_push43_notcmp41_pop43_output_regs_ready)
		begin
			local_bb4_notcmp41_push43_notcmp41_pop43_NO_SHIFT_REG <= local_bb4_notcmp41_push43_notcmp41_pop43_result;
			local_bb4_notcmp41_push43_notcmp41_pop43_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notcmp41_push43_notcmp41_pop43_stall_in))
			begin
				local_bb4_notcmp41_push43_notcmp41_pop43_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_notexitcond943_push44_notexitcond943_pop44_inputs_ready;
 reg local_bb4_notexitcond943_push44_notexitcond943_pop44_valid_out_NO_SHIFT_REG;
wire local_bb4_notexitcond943_push44_notexitcond943_pop44_stall_in;
wire local_bb4_notexitcond943_push44_notexitcond943_pop44_output_regs_ready;
wire local_bb4_notexitcond943_push44_notexitcond943_pop44_result;
wire local_bb4_notexitcond943_push44_notexitcond943_pop44_fu_valid_out;
wire local_bb4_notexitcond943_push44_notexitcond943_pop44_fu_stall_out;
 reg local_bb4_notexitcond943_push44_notexitcond943_pop44_NO_SHIFT_REG;
wire local_bb4_notexitcond943_push44_notexitcond943_pop44_causedstall;

acl_push local_bb4_notexitcond943_push44_notexitcond943_pop44_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_notexitcond943_pop44_c0_ene15),
	.stall_out(local_bb4_notexitcond943_push44_notexitcond943_pop44_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond943_push44_notexitcond943_pop44_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond943_push44_notexitcond943_pop44_result),
	.feedback_out(feedback_data_out_44),
	.feedback_valid_out(feedback_valid_out_44),
	.feedback_stall_in(feedback_stall_in_44)
);

defparam local_bb4_notexitcond943_push44_notexitcond943_pop44_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond943_push44_notexitcond943_pop44_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond943_push44_notexitcond943_pop44_feedback.FIFO_DEPTH = 9;
defparam local_bb4_notexitcond943_push44_notexitcond943_pop44_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_notexitcond943_push44_notexitcond943_pop44_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond943_push44_notexitcond943_pop44_inputs_ready = 1'b1;
assign local_bb4_notexitcond943_push44_notexitcond943_pop44_output_regs_ready = 1'b1;
assign local_bb4_notexitcond943_pop44_c0_ene15_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_13 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_27 = 1'b0;
assign local_bb4_notexitcond943_push44_notexitcond943_pop44_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond943_push44_notexitcond943_pop44_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond943_push44_notexitcond943_pop44_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond943_push44_notexitcond943_pop44_output_regs_ready)
		begin
			local_bb4_notexitcond943_push44_notexitcond943_pop44_NO_SHIFT_REG <= local_bb4_notexitcond943_push44_notexitcond943_pop44_result;
			local_bb4_notexitcond943_push44_notexitcond943_pop44_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond943_push44_notexitcond943_pop44_stall_in))
			begin
				local_bb4_notexitcond943_push44_notexitcond943_pop44_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4__push47__pop47_inputs_ready;
 reg local_bb4__push47__pop47_valid_out_NO_SHIFT_REG;
wire local_bb4__push47__pop47_stall_in;
wire local_bb4__push47__pop47_output_regs_ready;
wire local_bb4__push47__pop47_result;
wire local_bb4__push47__pop47_fu_valid_out;
wire local_bb4__push47__pop47_fu_stall_out;
 reg local_bb4__push47__pop47_NO_SHIFT_REG;
wire local_bb4__push47__pop47_causedstall;

acl_push local_bb4__push47__pop47_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4__pop47_c0_ene16),
	.stall_out(local_bb4__push47__pop47_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__push47__pop47_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4__push47__pop47_result),
	.feedback_out(feedback_data_out_47),
	.feedback_valid_out(feedback_valid_out_47),
	.feedback_stall_in(feedback_stall_in_47)
);

defparam local_bb4__push47__pop47_feedback.STALLFREE = 1;
defparam local_bb4__push47__pop47_feedback.DATA_WIDTH = 1;
defparam local_bb4__push47__pop47_feedback.FIFO_DEPTH = 9;
defparam local_bb4__push47__pop47_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4__push47__pop47_feedback.STYLE = "REGULAR";

assign local_bb4__push47__pop47_inputs_ready = 1'b1;
assign local_bb4__push47__pop47_output_regs_ready = 1'b1;
assign local_bb4__pop47_c0_ene16_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_14 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_28 = 1'b0;
assign local_bb4__push47__pop47_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4__push47__pop47_NO_SHIFT_REG <= 'x;
		local_bb4__push47__pop47_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4__push47__pop47_output_regs_ready)
		begin
			local_bb4__push47__pop47_NO_SHIFT_REG <= local_bb4__push47__pop47_result;
			local_bb4__push47__pop47_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4__push47__pop47_stall_in))
			begin
				local_bb4__push47__pop47_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notexitcond_notexit_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notexitcond_notexit_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_15 = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG = rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_j_35_push30_inc_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_j_35_push30_inc_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_j_35_push30_inc_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_j_35_push30_inc_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_j_35_push30_inc_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_j_35_push30_inc_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_j_35_push30_inc_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_j_35_push30_inc_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_j_35_push30_inc_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_j_35_push30_inc_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_j_35_push30_inc_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_j_35_push30_inc_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_j_35_push30_inc_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_j_35_push30_inc_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_j_35_push30_inc_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_j_35_push30_inc_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_j_35_push30_inc_0_reg_11_fifo.DATA_WIDTH = 32;
defparam rnode_10to11_bb4_j_35_push30_inc_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_j_35_push30_inc_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_j_35_push30_inc_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_j_35_push30_inc_stall_in = 1'b0;
assign rnode_10to11_bb4_j_35_push30_inc_0_NO_SHIFT_REG = rnode_10to11_bb4_j_35_push30_inc_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_j_35_push30_inc_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_j_35_push30_inc_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_mul2445_push46_mul2445_pop46_inputs_ready;
 reg local_bb4_mul2445_push46_mul2445_pop46_valid_out_NO_SHIFT_REG;
wire local_bb4_mul2445_push46_mul2445_pop46_stall_in;
wire local_bb4_mul2445_push46_mul2445_pop46_output_regs_ready;
wire [31:0] local_bb4_mul2445_push46_mul2445_pop46_result;
wire local_bb4_mul2445_push46_mul2445_pop46_fu_valid_out;
wire local_bb4_mul2445_push46_mul2445_pop46_fu_stall_out;
 reg [31:0] local_bb4_mul2445_push46_mul2445_pop46_NO_SHIFT_REG;
wire local_bb4_mul2445_push46_mul2445_pop46_causedstall;

acl_push local_bb4_mul2445_push46_mul2445_pop46_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_NO_SHIFT_REG),
	.stall_out(local_bb4_mul2445_push46_mul2445_pop46_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_mul2445_push46_mul2445_pop46_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_mul2445_push46_mul2445_pop46_result),
	.feedback_out(feedback_data_out_46),
	.feedback_valid_out(feedback_valid_out_46),
	.feedback_stall_in(feedback_stall_in_46)
);

defparam local_bb4_mul2445_push46_mul2445_pop46_feedback.STALLFREE = 1;
defparam local_bb4_mul2445_push46_mul2445_pop46_feedback.DATA_WIDTH = 32;
defparam local_bb4_mul2445_push46_mul2445_pop46_feedback.FIFO_DEPTH = 9;
defparam local_bb4_mul2445_push46_mul2445_pop46_feedback.MIN_FIFO_LATENCY = 8;
defparam local_bb4_mul2445_push46_mul2445_pop46_feedback.STYLE = "REGULAR";

assign local_bb4_mul2445_push46_mul2445_pop46_inputs_ready = 1'b1;
assign local_bb4_mul2445_push46_mul2445_pop46_output_regs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_0 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_14 = 1'b0;
assign rnode_9to10_bb4_mul2445_pop46_c0_ene464_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_mul2445_push46_mul2445_pop46_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul2445_push46_mul2445_pop46_NO_SHIFT_REG <= 'x;
		local_bb4_mul2445_push46_mul2445_pop46_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul2445_push46_mul2445_pop46_output_regs_ready)
		begin
			local_bb4_mul2445_push46_mul2445_pop46_NO_SHIFT_REG <= local_bb4_mul2445_push46_mul2445_pop46_result;
			local_bb4_mul2445_push46_mul2445_pop46_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul2445_push46_mul2445_pop46_stall_in))
			begin
				local_bb4_mul2445_push46_mul2445_pop46_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_idxprom26_stall_local;
wire [63:0] local_bb4_idxprom26;

assign local_bb4_idxprom26[63:32] = 32'h0;
assign local_bb4_idxprom26[31:0] = rnode_9to10_bb4_add25_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_arrayidx27_valid_out;
wire local_bb4_arrayidx27_stall_in;
wire local_bb4_arrayidx27_inputs_ready;
wire local_bb4_arrayidx27_stall_local;
wire [63:0] local_bb4_arrayidx27;

assign local_bb4_arrayidx27_inputs_ready = rnode_9to10_bb4_add25_0_valid_out_NO_SHIFT_REG;
assign local_bb4_arrayidx27 = ((input_in & 64'hFFFFFFFFFFFFFC00) + ((local_bb4_idxprom26 & 64'hFFFFFFFF) << 6'h2));
assign local_bb4_arrayidx27_valid_out = 1'b1;
assign rnode_9to10_bb4_add25_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_arrayidx27_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx27_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx27_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx27_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx27_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx27_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx27_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx27_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_arrayidx27_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_arrayidx27_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_arrayidx27_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_arrayidx27_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_arrayidx27_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in((local_bb4_arrayidx27 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_10to11_bb4_arrayidx27_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_arrayidx27_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_arrayidx27_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_arrayidx27_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_arrayidx27_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_arrayidx27_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_arrayidx27_stall_in = 1'b0;
assign rnode_10to11_bb4_arrayidx27_0_NO_SHIFT_REG = rnode_10to11_bb4_arrayidx27_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_arrayidx27_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx27_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi275_stall_local;
wire [447:0] local_bb4_c0_exi275;

assign local_bb4_c0_exi275[63:0] = local_bb4_c0_exi174[63:0];
assign local_bb4_c0_exi275[127:64] = (rnode_10to11_bb4_arrayidx27_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign local_bb4_c0_exi275[447:128] = local_bb4_c0_exi174[447:128];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi376_stall_local;
wire [447:0] local_bb4_c0_exi376;

assign local_bb4_c0_exi376[127:0] = local_bb4_c0_exi275[127:0];
assign local_bb4_c0_exi376[128] = rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_NO_SHIFT_REG;
assign local_bb4_c0_exi376[447:129] = local_bb4_c0_exi275[447:129];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi477_stall_local;
wire [447:0] local_bb4_c0_exi477;

assign local_bb4_c0_exi477[159:0] = local_bb4_c0_exi376[159:0];
assign local_bb4_c0_exi477[191:160] = rnode_10to11_bb4__pop42_c0_ene666_0_NO_SHIFT_REG;
assign local_bb4_c0_exi477[447:192] = local_bb4_c0_exi376[447:192];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi578_stall_local;
wire [447:0] local_bb4_c0_exi578;

assign local_bb4_c0_exi578[191:0] = local_bb4_c0_exi477[191:0];
assign local_bb4_c0_exi578[192] = rnode_9to11_bb4_var__0_NO_SHIFT_REG;
assign local_bb4_c0_exi578[447:193] = local_bb4_c0_exi477[447:193];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi679_stall_local;
wire [447:0] local_bb4_c0_exi679;

assign local_bb4_c0_exi679[199:0] = local_bb4_c0_exi578[199:0];
assign local_bb4_c0_exi679[200] = rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG;
assign local_bb4_c0_exi679[447:201] = local_bb4_c0_exi578[447:201];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi780_stall_local;
wire [447:0] local_bb4_c0_exi780;

assign local_bb4_c0_exi780[223:0] = local_bb4_c0_exi679[223:0];
assign local_bb4_c0_exi780[255:224] = rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_NO_SHIFT_REG;
assign local_bb4_c0_exi780[447:256] = local_bb4_c0_exi679[447:256];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi881_stall_local;
wire [447:0] local_bb4_c0_exi881;

assign local_bb4_c0_exi881[255:0] = local_bb4_c0_exi780[255:0];
assign local_bb4_c0_exi881[256] = rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_NO_SHIFT_REG;
assign local_bb4_c0_exi881[447:257] = local_bb4_c0_exi780[447:257];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi982_stall_local;
wire [447:0] local_bb4_c0_exi982;

assign local_bb4_c0_exi982[263:0] = local_bb4_c0_exi881[263:0];
assign local_bb4_c0_exi982[264] = rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_NO_SHIFT_REG;
assign local_bb4_c0_exi982[447:265] = local_bb4_c0_exi881[447:265];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi1083_stall_local;
wire [447:0] local_bb4_c0_exi1083;

assign local_bb4_c0_exi1083[319:0] = local_bb4_c0_exi982[319:0];
assign local_bb4_c0_exi1083[383:320] = rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_NO_SHIFT_REG;
assign local_bb4_c0_exi1083[447:384] = local_bb4_c0_exi982[447:384];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi1184_stall_local;
wire [447:0] local_bb4_c0_exi1184;

assign local_bb4_c0_exi1184[383:0] = local_bb4_c0_exi1083[383:0];
assign local_bb4_c0_exi1184[384] = rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_NO_SHIFT_REG;
assign local_bb4_c0_exi1184[447:385] = local_bb4_c0_exi1083[447:385];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi1285_stall_local;
wire [447:0] local_bb4_c0_exi1285;

assign local_bb4_c0_exi1285[391:0] = local_bb4_c0_exi1184[391:0];
assign local_bb4_c0_exi1285[392] = rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_NO_SHIFT_REG;
assign local_bb4_c0_exi1285[447:393] = local_bb4_c0_exi1184[447:393];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi1386_valid_out;
wire local_bb4_c0_exi1386_stall_in;
wire local_bb4_c0_exi1386_inputs_ready;
wire local_bb4_c0_exi1386_stall_local;
wire [447:0] local_bb4_c0_exi1386;

assign local_bb4_c0_exi1386_inputs_ready = (rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4__pop42_c0_ene666_0_valid_out_NO_SHIFT_REG & rnode_9to11_bb4_var__0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_arrayidx27_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4__pop47_c0_ene16_0_valid_out_NO_SHIFT_REG);
assign local_bb4_c0_exi1386[399:0] = local_bb4_c0_exi1285[399:0];
assign local_bb4_c0_exi1386[400] = rnode_10to11_bb4__pop47_c0_ene16_0_NO_SHIFT_REG;
assign local_bb4_c0_exi1386[447:401] = local_bb4_c0_exi1285[447:401];
assign local_bb4_c0_exi1386_valid_out = 1'b1;
assign rnode_10to11_bb4_memdep_phi1_or39_pop41_c0_ene565_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__pop42_c0_ene666_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_var__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_forked1644_pop45_c0_ene161_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx27_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_mul3724_pop34_c0_ene868_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notcmp1127_pop35_c0_ene969_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond1430_pop36_c0_ene1070_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_indvars_iv_pop1037_pop39_c0_ene1373_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notcmp41_pop43_c0_ene14_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond943_pop44_c0_ene15_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__pop47_c0_ene16_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_c0_exit87_c0_exi1386_inputs_ready;
 reg local_bb4_c0_exit87_c0_exi1386_valid_out_0_NO_SHIFT_REG;
wire local_bb4_c0_exit87_c0_exi1386_stall_in_0;
 reg local_bb4_c0_exit87_c0_exi1386_valid_out_1_NO_SHIFT_REG;
wire local_bb4_c0_exit87_c0_exi1386_stall_in_1;
 reg local_bb4_c0_exit87_c0_exi1386_valid_out_2_NO_SHIFT_REG;
wire local_bb4_c0_exit87_c0_exi1386_stall_in_2;
 reg [447:0] local_bb4_c0_exit87_c0_exi1386_NO_SHIFT_REG;
wire [447:0] local_bb4_c0_exit87_c0_exi1386_in;
wire local_bb4_c0_exit87_c0_exi1386_valid;
wire local_bb4_c0_exit87_c0_exi1386_causedstall;

acl_stall_free_sink local_bb4_c0_exit87_c0_exi1386_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb4_c0_exi1386),
	.data_out(local_bb4_c0_exit87_c0_exi1386_in),
	.input_accepted(local_bb4_c0_enter60_c0_eni16_input_accepted),
	.valid_out(local_bb4_c0_exit87_c0_exi1386_valid),
	.stall_in(~(local_bb4_c0_exit87_c0_exi1386_output_regs_ready)),
	.stall_entry(local_bb4_c0_exit87_c0_exi1386_entry_stall),
	.valid_in(local_bb4_c0_exit87_c0_exi1386_valid_in),
	.IIphases(local_bb4_c0_exit87_c0_exi1386_phases),
	.inc_pipelined_thread(local_bb4_c0_enter60_c0_eni16_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb4_c0_enter60_c0_eni16_dec_pipelined_thread)
);

defparam local_bb4_c0_exit87_c0_exi1386_instance.DATA_WIDTH = 448;
defparam local_bb4_c0_exit87_c0_exi1386_instance.PIPELINE_DEPTH = 15;
defparam local_bb4_c0_exit87_c0_exi1386_instance.SHARINGII = 1;
defparam local_bb4_c0_exit87_c0_exi1386_instance.SCHEDULEII = 1;
defparam local_bb4_c0_exit87_c0_exi1386_instance.ALWAYS_THROTTLE = 0;

assign local_bb4_c0_exit87_c0_exi1386_inputs_ready = 1'b1;
assign local_bb4_c0_exit87_c0_exi1386_output_regs_ready = ((~(local_bb4_c0_exit87_c0_exi1386_valid_out_0_NO_SHIFT_REG) | ~(local_bb4_c0_exit87_c0_exi1386_stall_in_0)) & (~(local_bb4_c0_exit87_c0_exi1386_valid_out_1_NO_SHIFT_REG) | ~(local_bb4_c0_exit87_c0_exi1386_stall_in_1)) & (~(local_bb4_c0_exit87_c0_exi1386_valid_out_2_NO_SHIFT_REG) | ~(local_bb4_c0_exit87_c0_exi1386_stall_in_2)));
assign local_bb4_c0_exit87_c0_exi1386_valid_in = SFC_2_VALID_10_11_0_NO_SHIFT_REG;
assign local_bb4_c0_exi1386_stall_in = 1'b0;
assign local_bb4_mul2445_push46_mul2445_pop46_stall_in = 1'b0;
assign local_bb4_forked1644_push45_forked1644_pop45_stall_in = 1'b0;
assign local_bb4__push42__pop42_stall_in = 1'b0;
assign local_bb4_memdep_phi1_or39_push41_memdep_phi1_or39_pop41_stall_in = 1'b0;
assign local_bb4__push40__pop40_stall_in = 1'b0;
assign local_bb4_pixel_y_020_pop821_push33_pixel_y_020_pop821_pop33_stall_in = 1'b0;
assign local_bb4_mul3724_push34_mul3724_pop34_stall_in = 1'b0;
assign local_bb4_notcmp1127_push35_notcmp1127_pop35_stall_in = 1'b0;
assign local_bb4_notexitcond1430_push36_notexitcond1430_pop36_stall_in = 1'b0;
assign local_bb4_memdep_phi1_pop933_push37_memdep_phi1_pop933_pop37_stall_in = 1'b0;
assign local_bb4_mul535_push38_mul535_pop38_stall_in = 1'b0;
assign local_bb4_indvars_iv_pop1037_push39_indvars_iv_pop1037_pop39_stall_in = 1'b0;
assign local_bb4_notcmp41_push43_notcmp41_pop43_stall_in = 1'b0;
assign local_bb4_notexitcond943_push44_notexitcond943_pop44_stall_in = 1'b0;
assign local_bb4__push47__pop47_stall_in = 1'b0;
assign SFC_2_VALID_10_11_0_stall_in = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_j_35_push30_inc_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_c0_exit87_c0_exi1386_causedstall = (1'b1 && (1'b0 && !(~(local_bb4_c0_exit87_c0_exi1386_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c0_exit87_c0_exi1386_NO_SHIFT_REG <= 'x;
		local_bb4_c0_exit87_c0_exi1386_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_c0_exit87_c0_exi1386_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_c0_exit87_c0_exi1386_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c0_exit87_c0_exi1386_output_regs_ready)
		begin
			local_bb4_c0_exit87_c0_exi1386_NO_SHIFT_REG <= local_bb4_c0_exit87_c0_exi1386_in;
			local_bb4_c0_exit87_c0_exi1386_valid_out_0_NO_SHIFT_REG <= local_bb4_c0_exit87_c0_exi1386_valid;
			local_bb4_c0_exit87_c0_exi1386_valid_out_1_NO_SHIFT_REG <= local_bb4_c0_exit87_c0_exi1386_valid;
			local_bb4_c0_exit87_c0_exi1386_valid_out_2_NO_SHIFT_REG <= local_bb4_c0_exit87_c0_exi1386_valid;
		end
		else
		begin
			if (~(local_bb4_c0_exit87_c0_exi1386_stall_in_0))
			begin
				local_bb4_c0_exit87_c0_exi1386_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c0_exit87_c0_exi1386_stall_in_1))
			begin
				local_bb4_c0_exit87_c0_exi1386_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c0_exit87_c0_exi1386_stall_in_2))
			begin
				local_bb4_c0_exit87_c0_exi1386_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe289_valid_out;
wire local_bb4_c0_exe289_stall_in;
wire local_bb4_c0_exe289_inputs_ready;
wire local_bb4_c0_exe289_stall_local;
wire [63:0] local_bb4_c0_exe289;

assign local_bb4_c0_exe289_inputs_ready = local_bb4_c0_exit87_c0_exi1386_valid_out_0_NO_SHIFT_REG;
assign local_bb4_c0_exe289 = local_bb4_c0_exit87_c0_exi1386_NO_SHIFT_REG[127:64];
assign local_bb4_c0_exe289_valid_out = local_bb4_c0_exe289_inputs_ready;
assign local_bb4_c0_exe289_stall_local = local_bb4_c0_exe289_stall_in;
assign local_bb4_c0_exit87_c0_exi1386_stall_in_0 = (|local_bb4_c0_exe289_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe390_valid_out;
wire local_bb4_c0_exe390_stall_in;
wire local_bb4_c0_exe390_inputs_ready;
wire local_bb4_c0_exe390_stall_local;
wire local_bb4_c0_exe390;

assign local_bb4_c0_exe390_inputs_ready = local_bb4_c0_exit87_c0_exi1386_valid_out_1_NO_SHIFT_REG;
assign local_bb4_c0_exe390 = local_bb4_c0_exit87_c0_exi1386_NO_SHIFT_REG[128];
assign local_bb4_c0_exe390_valid_out = local_bb4_c0_exe390_inputs_ready;
assign local_bb4_c0_exe390_stall_local = local_bb4_c0_exe390_stall_in;
assign local_bb4_c0_exit87_c0_exi1386_stall_in_1 = (|local_bb4_c0_exe390_stall_local);

// Register node:
//  * latency = 159
//  * capacity = 159
 logic rnode_16to175_bb4_c0_exit87_c0_exi1386_0_valid_out_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_in_NO_SHIFT_REG;
 logic [447:0] rnode_16to175_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [447:0] rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit87_c0_exi1386_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_16to175_bb4_c0_exit87_c0_exi1386_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb4_c0_exit87_c0_exi1386_NO_SHIFT_REG),
	.data_out(rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_fifo.DEPTH = 160;
defparam rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_fifo.DATA_WIDTH = 448;
defparam rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_fifo.IMPL = "ram";

assign rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_inputs_ready_NO_SHIFT_REG = local_bb4_c0_exit87_c0_exi1386_valid_out_2_NO_SHIFT_REG;
assign local_bb4_c0_exit87_c0_exi1386_stall_in_2 = rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_175_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit87_c0_exi1386_0_reg_175_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_in_reg_175_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_in_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit87_c0_exi1386_0_valid_out_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit87_c0_exi1386_0_valid_out_reg_175_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_ld__inputs_ready;
 reg local_bb4_ld__valid_out_NO_SHIFT_REG;
wire local_bb4_ld__stall_in;
wire local_bb4_ld__output_regs_ready;
wire local_bb4_ld__fu_stall_out;
wire local_bb4_ld__fu_valid_out;
wire [31:0] local_bb4_ld__lsu_dataout;
 reg [31:0] local_bb4_ld__NO_SHIFT_REG;
wire local_bb4_ld__causedstall;

lsu_top lsu_local_bb4_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb4_ld__fu_stall_out),
	.i_valid(local_bb4_ld__inputs_ready),
	.i_address((local_bb4_c0_exe289 & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(input_wii_var__u17),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb4_ld__output_regs_ready)),
	.o_valid(local_bb4_ld__fu_valid_out),
	.o_readdata(local_bb4_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb4_ld__active),
	.avm_address(avm_local_bb4_ld__address),
	.avm_read(avm_local_bb4_ld__read),
	.avm_readdata(avm_local_bb4_ld__readdata),
	.avm_write(avm_local_bb4_ld__write),
	.avm_writeack(avm_local_bb4_ld__writeack),
	.avm_burstcount(avm_local_bb4_ld__burstcount),
	.avm_writedata(avm_local_bb4_ld__writedata),
	.avm_byteenable(avm_local_bb4_ld__byteenable),
	.avm_waitrequest(avm_local_bb4_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb4_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb4_ld_.AWIDTH = 33;
defparam lsu_local_bb4_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb4_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb4_ld_.READ = 1;
defparam lsu_local_bb4_ld_.ATOMIC = 0;
defparam lsu_local_bb4_ld_.WIDTH = 32;
defparam lsu_local_bb4_ld_.MWIDTH = 512;
defparam lsu_local_bb4_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb4_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb4_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb4_ld_.MEMORY_SIDE_MEM_LATENCY = 99;
defparam lsu_local_bb4_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb4_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb4_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb4_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb4_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb4_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb4_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb4_ld_.USECACHING = 0;
defparam lsu_local_bb4_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb4_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb4_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb4_ld_.ADDRSPACE = 1;
defparam lsu_local_bb4_ld_.STYLE = "BURST-COALESCED";

assign local_bb4_ld__inputs_ready = (local_bb4_c0_exe289_valid_out & local_bb4_c0_exe390_valid_out & rnode_15to16_var__u17_0_valid_out_NO_SHIFT_REG);
assign local_bb4_ld__output_regs_ready = (&(~(local_bb4_ld__valid_out_NO_SHIFT_REG) | ~(local_bb4_ld__stall_in)));
assign local_bb4_c0_exe289_stall_in = (local_bb4_ld__fu_stall_out | ~(local_bb4_ld__inputs_ready));
assign local_bb4_c0_exe390_stall_in = (local_bb4_ld__fu_stall_out | ~(local_bb4_ld__inputs_ready));
assign rnode_15to16_var__u17_0_stall_in_NO_SHIFT_REG = (local_bb4_ld__fu_stall_out | ~(local_bb4_ld__inputs_ready));
assign local_bb4_ld__causedstall = (local_bb4_ld__inputs_ready && (local_bb4_ld__fu_stall_out && !(~(local_bb4_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_ld__NO_SHIFT_REG <= 'x;
		local_bb4_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_ld__output_regs_ready)
		begin
			local_bb4_ld__NO_SHIFT_REG <= local_bb4_ld__lsu_dataout;
			local_bb4_ld__valid_out_NO_SHIFT_REG <= local_bb4_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb4_ld__stall_in))
			begin
				local_bb4_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_NO_SHIFT_REG;
 logic [447:0] rnode_175to176_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_1_NO_SHIFT_REG;
 logic [447:0] rnode_175to176_bb4_c0_exit87_c0_exi1386_1_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_2_NO_SHIFT_REG;
 logic [447:0] rnode_175to176_bb4_c0_exit87_c0_exi1386_2_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_3_NO_SHIFT_REG;
 logic [447:0] rnode_175to176_bb4_c0_exit87_c0_exi1386_3_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [447:0] rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_176_NO_SHIFT_REG;
 reg rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_0_NO_SHIFT_REG;
 reg rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_3_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_16to175_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_fifo.DATA_WIDTH = 448;
defparam rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_fifo.IMPL = "ll_reg";

assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_inputs_ready_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit87_c0_exi1386_0_valid_out_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit87_c0_exi1386_0_stall_in_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_176_NO_SHIFT_REG = ((rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_0_NO_SHIFT_REG)) | 1'b0 | 1'b0 | (rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_3_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_3_NO_SHIFT_REG)));
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_NO_SHIFT_REG = (rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_0_NO_SHIFT_REG));
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_1_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_2_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_3_NO_SHIFT_REG = (rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_3_NO_SHIFT_REG));
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_1_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_2_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_3_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_reg_176_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_0_NO_SHIFT_REG <= (rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG & (rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_0_NO_SHIFT_REG | ~(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_NO_SHIFT_REG)) & rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_176_NO_SHIFT_REG);
		rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_3_NO_SHIFT_REG <= (rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_176_NO_SHIFT_REG & (rnode_175to176_bb4_c0_exit87_c0_exi1386_0_consumed_3_NO_SHIFT_REG | ~(rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_3_NO_SHIFT_REG)) & rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_176_NO_SHIFT_REG);
	end
end


// This section implements a staging register.
// 
wire rstag_176to176_bb4_ld__valid_out;
wire rstag_176to176_bb4_ld__stall_in;
wire rstag_176to176_bb4_ld__inputs_ready;
wire rstag_176to176_bb4_ld__stall_local;
 reg rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG;
wire rstag_176to176_bb4_ld__combined_valid;
 reg [31:0] rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_176to176_bb4_ld_;

assign rstag_176to176_bb4_ld__inputs_ready = local_bb4_ld__valid_out_NO_SHIFT_REG;
assign rstag_176to176_bb4_ld_ = (rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG ? rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG : local_bb4_ld__NO_SHIFT_REG);
assign rstag_176to176_bb4_ld__combined_valid = (rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG | rstag_176to176_bb4_ld__inputs_ready);
assign rstag_176to176_bb4_ld__valid_out = rstag_176to176_bb4_ld__combined_valid;
assign rstag_176to176_bb4_ld__stall_local = rstag_176to176_bb4_ld__stall_in;
assign local_bb4_ld__stall_in = (|rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_176to176_bb4_ld__stall_local)
		begin
			if (~(rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= rstag_176to176_bb4_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG <= local_bb4_ld__NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe188_stall_local;
wire local_bb4_c0_exe188;

assign local_bb4_c0_exe188 = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG[8];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe491_stall_local;
wire [31:0] local_bb4_c0_exe491;

assign local_bb4_c0_exe491 = rnode_175to176_bb4_c0_exit87_c0_exi1386_1_NO_SHIFT_REG[191:160];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe693_stall_local;
wire local_bb4_c0_exe693;

assign local_bb4_c0_exe693 = rnode_175to176_bb4_c0_exit87_c0_exi1386_2_NO_SHIFT_REG[200];

// Register node:
//  * latency = 16
//  * capacity = 16
 logic rnode_176to192_bb4_c0_exit87_c0_exi1386_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_in_NO_SHIFT_REG;
 logic [447:0] rnode_176to192_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG;
 logic rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_inputs_ready_NO_SHIFT_REG;
 logic [447:0] rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_NO_SHIFT_REG;
 logic rnode_176to192_bb4_c0_exit87_c0_exi1386_0_valid_out_reg_192_NO_SHIFT_REG;
 logic rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_in_reg_192_NO_SHIFT_REG;
 logic rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_192_NO_SHIFT_REG;

acl_data_fifo rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_in_reg_192_NO_SHIFT_REG),
	.valid_out(rnode_176to192_bb4_c0_exit87_c0_exi1386_0_valid_out_reg_192_NO_SHIFT_REG),
	.stall_out(rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_192_NO_SHIFT_REG),
	.data_in(rnode_175to176_bb4_c0_exit87_c0_exi1386_3_NO_SHIFT_REG),
	.data_out(rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_NO_SHIFT_REG)
);

defparam rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_fifo.DEPTH = 17;
defparam rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_fifo.DATA_WIDTH = 448;
defparam rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_fifo.IMPL = "ram";

assign rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_inputs_ready_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_3_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_3_NO_SHIFT_REG = rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_192_NO_SHIFT_REG;
assign rnode_176to192_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG = rnode_176to192_bb4_c0_exit87_c0_exi1386_0_reg_192_NO_SHIFT_REG;
assign rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_in_reg_192_NO_SHIFT_REG = rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_in_NO_SHIFT_REG;
assign rnode_176to192_bb4_c0_exit87_c0_exi1386_0_valid_out_NO_SHIFT_REG = rnode_176to192_bb4_c0_exit87_c0_exi1386_0_valid_out_reg_192_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni2_stall_local;
wire [127:0] local_bb4_c1_eni2;

assign local_bb4_c1_eni2[15:0] = local_bb4_c1_eni1[15:0];
assign local_bb4_c1_eni2[16] = local_bb4_c0_exe188;
assign local_bb4_c1_eni2[127:17] = local_bb4_c1_eni1[127:17];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_0_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_1_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_1_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_2_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_2_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_3_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_3_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_4_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_4_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_5_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_5_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_5_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_6_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_6_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_6_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_7_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_7_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_7_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_inputs_ready_NO_SHIFT_REG;
 logic [447:0] rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_193_NO_SHIFT_REG;
 logic rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_193_NO_SHIFT_REG;

acl_data_fifo rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_193_NO_SHIFT_REG),
	.valid_out(rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG),
	.stall_out(rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_193_NO_SHIFT_REG),
	.data_in(rnode_176to192_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG),
	.data_out(rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG)
);

defparam rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_fifo.DEPTH = 1;
defparam rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_fifo.DATA_WIDTH = 448;
defparam rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_fifo.IMPL = "ll_reg";

assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_inputs_ready_NO_SHIFT_REG = rnode_176to192_bb4_c0_exit87_c0_exi1386_0_valid_out_NO_SHIFT_REG;
assign rnode_176to192_bb4_c0_exit87_c0_exi1386_0_stall_in_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_out_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_0_reg_193_NO_SHIFT_REG = (rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_0_NO_SHIFT_REG | rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_1_NO_SHIFT_REG | rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_2_NO_SHIFT_REG | rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_3_NO_SHIFT_REG | rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_4_NO_SHIFT_REG | rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_5_NO_SHIFT_REG | rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_6_NO_SHIFT_REG | rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_7_NO_SHIFT_REG);
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_1_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_2_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_3_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_4_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_5_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_6_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_7_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_1_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_2_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_3_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_4_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_5_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_6_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_7_NO_SHIFT_REG = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_reg_193_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni3_stall_local;
wire [127:0] local_bb4_c1_eni3;

assign local_bb4_c1_eni3[31:0] = local_bb4_c1_eni2[31:0];
assign local_bb4_c1_eni3[63:32] = rstag_176to176_bb4_ld_;
assign local_bb4_c1_eni3[127:64] = local_bb4_c1_eni2[127:64];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe592_stall_local;
wire local_bb4_c0_exe592;

assign local_bb4_c0_exe592 = rnode_192to193_bb4_c0_exit87_c0_exi1386_0_NO_SHIFT_REG[192];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe794_stall_local;
wire [31:0] local_bb4_c0_exe794;

assign local_bb4_c0_exe794 = rnode_192to193_bb4_c0_exit87_c0_exi1386_1_NO_SHIFT_REG[255:224];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe895_stall_local;
wire local_bb4_c0_exe895;

assign local_bb4_c0_exe895 = rnode_192to193_bb4_c0_exit87_c0_exi1386_2_NO_SHIFT_REG[256];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe996_stall_local;
wire local_bb4_c0_exe996;

assign local_bb4_c0_exe996 = rnode_192to193_bb4_c0_exit87_c0_exi1386_3_NO_SHIFT_REG[264];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe1097_stall_local;
wire [63:0] local_bb4_c0_exe1097;

assign local_bb4_c0_exe1097 = rnode_192to193_bb4_c0_exit87_c0_exi1386_4_NO_SHIFT_REG[383:320];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe1198_stall_local;
wire local_bb4_c0_exe1198;

assign local_bb4_c0_exe1198 = rnode_192to193_bb4_c0_exit87_c0_exi1386_5_NO_SHIFT_REG[384];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe1299_valid_out;
wire local_bb4_c0_exe1299_stall_in;
wire local_bb4_c0_exe1198_valid_out;
wire local_bb4_c0_exe1198_stall_in;
wire local_bb4_c0_exe1097_valid_out;
wire local_bb4_c0_exe1097_stall_in;
wire local_bb4_c0_exe996_valid_out;
wire local_bb4_c0_exe996_stall_in;
wire local_bb4_c0_exe895_valid_out;
wire local_bb4_c0_exe895_stall_in;
wire local_bb4_c0_exe794_valid_out;
wire local_bb4_c0_exe794_stall_in;
wire local_bb4_c0_exe592_valid_out;
wire local_bb4_c0_exe592_stall_in;
wire local_bb4_c0_exe1299_inputs_ready;
wire local_bb4_c0_exe1299_stall_local;
wire local_bb4_c0_exe1299;

assign local_bb4_c0_exe1299_inputs_ready = (rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_6_NO_SHIFT_REG & rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_5_NO_SHIFT_REG & rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_4_NO_SHIFT_REG & rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_3_NO_SHIFT_REG & rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_2_NO_SHIFT_REG & rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_1_NO_SHIFT_REG & rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_c0_exe1299 = rnode_192to193_bb4_c0_exit87_c0_exi1386_6_NO_SHIFT_REG[392];
assign local_bb4_c0_exe1299_stall_local = (local_bb4_c0_exe1299_stall_in | local_bb4_c0_exe1198_stall_in | local_bb4_c0_exe1097_stall_in | local_bb4_c0_exe996_stall_in | local_bb4_c0_exe895_stall_in | local_bb4_c0_exe794_stall_in | local_bb4_c0_exe592_stall_in);
assign local_bb4_c0_exe1299_valid_out = local_bb4_c0_exe1299_inputs_ready;
assign local_bb4_c0_exe1198_valid_out = local_bb4_c0_exe1299_inputs_ready;
assign local_bb4_c0_exe1097_valid_out = local_bb4_c0_exe1299_inputs_ready;
assign local_bb4_c0_exe996_valid_out = local_bb4_c0_exe1299_inputs_ready;
assign local_bb4_c0_exe895_valid_out = local_bb4_c0_exe1299_inputs_ready;
assign local_bb4_c0_exe794_valid_out = local_bb4_c0_exe1299_inputs_ready;
assign local_bb4_c0_exe592_valid_out = local_bb4_c0_exe1299_inputs_ready;
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_6_NO_SHIFT_REG = (local_bb4_c0_exe1299_stall_local | ~(local_bb4_c0_exe1299_inputs_ready));
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_5_NO_SHIFT_REG = (local_bb4_c0_exe1299_stall_local | ~(local_bb4_c0_exe1299_inputs_ready));
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_4_NO_SHIFT_REG = (local_bb4_c0_exe1299_stall_local | ~(local_bb4_c0_exe1299_inputs_ready));
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_3_NO_SHIFT_REG = (local_bb4_c0_exe1299_stall_local | ~(local_bb4_c0_exe1299_inputs_ready));
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_2_NO_SHIFT_REG = (local_bb4_c0_exe1299_stall_local | ~(local_bb4_c0_exe1299_inputs_ready));
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_1_NO_SHIFT_REG = (local_bb4_c0_exe1299_stall_local | ~(local_bb4_c0_exe1299_inputs_ready));
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c0_exe1299_stall_local | ~(local_bb4_c0_exe1299_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni4_stall_local;
wire [127:0] local_bb4_c1_eni4;

assign local_bb4_c1_eni4[63:0] = local_bb4_c1_eni3[63:0];
assign local_bb4_c1_eni4[95:64] = local_bb4_c0_exe491;
assign local_bb4_c1_eni4[127:96] = local_bb4_c1_eni3[127:96];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni5_stall_local;
wire [127:0] local_bb4_c1_eni5;

assign local_bb4_c1_eni5[95:0] = local_bb4_c1_eni4[95:0];
assign local_bb4_c1_eni5[96] = rcnode_175to176_rc0_forked_0_NO_SHIFT_REG[1];
assign local_bb4_c1_eni5[127:97] = local_bb4_c1_eni4[127:97];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni6_valid_out;
wire local_bb4_c1_eni6_stall_in;
wire local_bb4_c0_exe693_valid_out_1;
wire local_bb4_c0_exe693_stall_in_1;
wire local_bb4_c1_eni6_inputs_ready;
wire local_bb4_c1_eni6_stall_local;
wire [127:0] local_bb4_c1_eni6;

assign local_bb4_c1_eni6_inputs_ready = (rcnode_175to176_rc0_forked_0_valid_out_0_NO_SHIFT_REG & rstag_176to176_bb4_ld__valid_out & rcnode_175to176_rc0_forked_0_valid_out_2_NO_SHIFT_REG & rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb4_c0_exit87_c0_exi1386_0_valid_out_2_NO_SHIFT_REG);
assign local_bb4_c1_eni6[103:0] = local_bb4_c1_eni5[103:0];
assign local_bb4_c1_eni6[104] = local_bb4_c0_exe693;
assign local_bb4_c1_eni6[127:105] = local_bb4_c1_eni5[127:105];
assign local_bb4_c1_eni6_stall_local = (local_bb4_c1_eni6_stall_in | local_bb4_c0_exe693_stall_in_1);
assign local_bb4_c1_eni6_valid_out = local_bb4_c1_eni6_inputs_ready;
assign local_bb4_c0_exe693_valid_out_1 = local_bb4_c1_eni6_inputs_ready;
assign rcnode_175to176_rc0_forked_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rstag_176to176_bb4_ld__stall_in = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rcnode_175to176_rc0_forked_0_stall_in_2_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_1_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rnode_175to176_bb4_c0_exit87_c0_exi1386_0_stall_in_2_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb4_c1_enter_c1_eni6_inputs_ready;
 reg local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_0;
 reg local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_1;
 reg local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_2;
 reg local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_3;
 reg local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_4;
 reg local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_5;
 reg local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_6;
wire local_bb4_c1_enter_c1_eni6_output_regs_ready;
 reg [127:0] local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_input_accepted;
 reg local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG;
wire local_bb4_c1_exit_c1_exi2_entry_stall;
wire local_bb4_c1_exit_c1_exi2_output_regs_ready;
wire [12:0] local_bb4_c1_exit_c1_exi2_valid_bits;
wire local_bb4_c1_exit_c1_exi2_valid_in;
wire local_bb4_c1_exit_c1_exi2_phases;
wire local_bb4_c1_enter_c1_eni6_inc_pipelined_thread;
wire local_bb4_c1_enter_c1_eni6_dec_pipelined_thread;
wire local_bb4_c1_enter_c1_eni6_causedstall;

assign local_bb4_c1_enter_c1_eni6_inputs_ready = (local_bb4_c1_eni6_valid_out & local_bb4_c0_exe693_valid_out_1 & rcnode_175to176_rc0_forked_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_c1_enter_c1_eni6_output_regs_ready = 1'b1;
assign local_bb4_c1_enter_c1_eni6_input_accepted = (local_bb4_c1_enter_c1_eni6_inputs_ready && !(local_bb4_c1_exit_c1_exi2_entry_stall));
assign local_bb4_c1_enter_c1_eni6_inc_pipelined_thread = rcnode_175to176_rc0_forked_0_NO_SHIFT_REG[0];
assign local_bb4_c1_enter_c1_eni6_dec_pipelined_thread = ~(local_bb4_c0_exe693);
assign local_bb4_c1_eni6_stall_in = ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign local_bb4_c0_exe693_stall_in_1 = ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign rcnode_175to176_rc0_forked_0_stall_in_1_NO_SHIFT_REG = ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign local_bb4_c1_enter_c1_eni6_causedstall = (1'b1 && ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG <= local_bb4_c1_enter_c1_eni6_input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG <= 'x;
		local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c1_enter_c1_eni6_output_regs_ready)
		begin
			local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG <= local_bb4_c1_eni6;
			local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_0))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_1))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_2))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_3))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_4))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_5))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_6))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene1_stall_local;
wire local_bb4_c1_ene1;

assign local_bb4_c1_ene1 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[8];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene2_stall_local;
wire local_bb4_c1_ene2;

assign local_bb4_c1_ene2 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[16];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene3_stall_local;
wire [31:0] local_bb4_c1_ene3;

assign local_bb4_c1_ene3 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene4_stall_local;
wire [31:0] local_bb4_c1_ene4;

assign local_bb4_c1_ene4 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[95:64];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene5_stall_local;
wire local_bb4_c1_ene5;

assign local_bb4_c1_ene5 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[96];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene6_stall_local;
wire local_bb4_c1_ene6;

assign local_bb4_c1_ene6 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[104];

// This section implements an unregistered operation.
// 
wire SFC_3_VALID_177_177_0_stall_local;
wire SFC_3_VALID_177_177_0;

assign SFC_3_VALID_177_177_0 = local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_forked_and_stall_local;
wire local_bb4_forked_and;

assign local_bb4_forked_and = (local_bb4_c1_ene1 & local_bb4_c1_ene2);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u24_stall_local;
wire [31:0] local_bb4_var__u24;

assign local_bb4_var__u24 = local_bb4_c1_ene3;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u25_stall_local;
wire [31:0] local_bb4_var__u25;

assign local_bb4_var__u25 = local_bb4_c1_ene4;

// This section implements an unregistered operation.
// 
wire local_bb4_notexitcond546_pop48_c1_ene5_stall_local;
wire local_bb4_notexitcond546_pop48_c1_ene5;
wire local_bb4_notexitcond546_pop48_c1_ene5_fu_valid_out;
wire local_bb4_notexitcond546_pop48_c1_ene5_fu_stall_out;

acl_pop local_bb4_notexitcond546_pop48_c1_ene5_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_c1_ene1),
	.predicate(1'b0),
	.data_in(local_bb4_c1_ene5),
	.stall_out(local_bb4_notexitcond546_pop48_c1_ene5_fu_stall_out),
	.valid_in(SFC_3_VALID_177_177_0),
	.valid_out(local_bb4_notexitcond546_pop48_c1_ene5_fu_valid_out),
	.stall_in(local_bb4_notexitcond546_pop48_c1_ene5_stall_local),
	.data_out(local_bb4_notexitcond546_pop48_c1_ene5),
	.feedback_in(feedback_data_in_48),
	.feedback_valid_in(feedback_valid_in_48),
	.feedback_stall_out(feedback_stall_out_48)
);

defparam local_bb4_notexitcond546_pop48_c1_ene5_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_notexitcond546_pop48_c1_ene5_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond546_pop48_c1_ene5_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond546_pop48_c1_ene5_stall_local = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and2_i_stall_local;
wire [31:0] local_bb4_and2_i;

assign local_bb4_and2_i = (local_bb4_var__u24 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i_stall_local;
wire [31:0] local_bb4_and12_i;

assign local_bb4_and12_i = (local_bb4_var__u24 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i_stall_local;
wire [31:0] local_bb4_xor_i;

assign local_bb4_xor_i = (local_bb4_var__u25 ^ 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_forked_and_valid_out;
wire local_bb4_forked_and_stall_in;
wire local_bb4_notexitcond546_pop48_c1_ene5_valid_out_0;
wire local_bb4_notexitcond546_pop48_c1_ene5_stall_in_0;
wire SFC_3_VALID_177_177_0_valid_out_0;
wire SFC_3_VALID_177_177_0_stall_in_0;
wire SFC_3_VALID_177_177_0_valid_out_2;
wire SFC_3_VALID_177_177_0_stall_in_2;
wire local_bb4_c1_ene6_valid_out_0;
wire local_bb4_c1_ene6_stall_in_0;
wire local_bb4_notexitcond_or_valid_out;
wire local_bb4_notexitcond_or_stall_in;
wire local_bb4_notexitcond_or_inputs_ready;
wire local_bb4_notexitcond_or_stall_local;
wire local_bb4_notexitcond_or;

assign local_bb4_notexitcond_or_inputs_ready = (local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG);
assign local_bb4_notexitcond_or = (local_bb4_c1_ene6 | local_bb4_notexitcond546_pop48_c1_ene5);
assign local_bb4_forked_and_valid_out = 1'b1;
assign local_bb4_notexitcond546_pop48_c1_ene5_valid_out_0 = 1'b1;
assign SFC_3_VALID_177_177_0_valid_out_0 = 1'b1;
assign SFC_3_VALID_177_177_0_valid_out_2 = 1'b1;
assign local_bb4_c1_ene6_valid_out_0 = 1'b1;
assign local_bb4_notexitcond_or_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_0 = 1'b0;
assign local_bb4_c1_enter_c1_eni6_stall_in_1 = 1'b0;
assign local_bb4_c1_enter_c1_eni6_stall_in_4 = 1'b0;
assign local_bb4_c1_enter_c1_eni6_stall_in_6 = 1'b0;
assign local_bb4_c1_enter_c1_eni6_stall_in_5 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_stall_local;
wire [31:0] local_bb4_shr3_i;

assign local_bb4_shr3_i = ((local_bb4_and2_i & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_stall_local;
wire [31:0] local_bb4_and_i;

assign local_bb4_and_i = (local_bb4_xor_i >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i_stall_local;
wire [31:0] local_bb4_and10_i;

assign local_bb4_and10_i = (local_bb4_xor_i & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_forked_and_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_forked_and_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_forked_and_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_forked_and_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_forked_and_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_forked_and_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_forked_and_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_forked_and),
	.data_out(rnode_177to178_bb4_forked_and_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_forked_and_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_forked_and_0_reg_178_fifo.DATA_WIDTH = 1;
defparam rnode_177to178_bb4_forked_and_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_forked_and_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_forked_and_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_forked_and_stall_in = 1'b0;
assign rnode_177to178_bb4_forked_and_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_forked_and_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_forked_and_0_NO_SHIFT_REG = rnode_177to178_bb4_forked_and_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_forked_and_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_forked_and_1_NO_SHIFT_REG = rnode_177to178_bb4_forked_and_0_reg_178_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_177_178_0_inputs_ready;
 reg SFC_3_VALID_177_178_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_177_178_0_stall_in_0;
 reg SFC_3_VALID_177_178_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_177_178_0_stall_in_1;
wire SFC_3_VALID_177_178_0_output_regs_ready;
 reg SFC_3_VALID_177_178_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_177_178_0_causedstall;

assign SFC_3_VALID_177_178_0_inputs_ready = 1'b1;
assign SFC_3_VALID_177_178_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_177_177_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_177_178_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_177_178_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_177_178_0_output_regs_ready)
		begin
			SFC_3_VALID_177_178_0_NO_SHIFT_REG <= SFC_3_VALID_177_177_0;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_notexitcond546_push48_notexitcond546_pop48_inputs_ready;
 reg local_bb4_notexitcond546_push48_notexitcond546_pop48_valid_out_NO_SHIFT_REG;
wire local_bb4_notexitcond546_push48_notexitcond546_pop48_stall_in;
wire local_bb4_notexitcond546_push48_notexitcond546_pop48_output_regs_ready;
wire local_bb4_notexitcond546_push48_notexitcond546_pop48_result;
wire local_bb4_notexitcond546_push48_notexitcond546_pop48_fu_valid_out;
wire local_bb4_notexitcond546_push48_notexitcond546_pop48_fu_stall_out;
 reg local_bb4_notexitcond546_push48_notexitcond546_pop48_NO_SHIFT_REG;
wire local_bb4_notexitcond546_push48_notexitcond546_pop48_causedstall;

acl_push local_bb4_notexitcond546_push48_notexitcond546_pop48_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_c1_ene6),
	.predicate(1'b0),
	.data_in(local_bb4_notexitcond546_pop48_c1_ene5),
	.stall_out(local_bb4_notexitcond546_push48_notexitcond546_pop48_fu_stall_out),
	.valid_in(SFC_3_VALID_177_177_0),
	.valid_out(local_bb4_notexitcond546_push48_notexitcond546_pop48_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond546_push48_notexitcond546_pop48_result),
	.feedback_out(feedback_data_out_48),
	.feedback_valid_out(feedback_valid_out_48),
	.feedback_stall_in(feedback_stall_in_48)
);

defparam local_bb4_notexitcond546_push48_notexitcond546_pop48_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond546_push48_notexitcond546_pop48_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond546_push48_notexitcond546_pop48_feedback.FIFO_DEPTH = 9;
defparam local_bb4_notexitcond546_push48_notexitcond546_pop48_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_notexitcond546_push48_notexitcond546_pop48_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond546_push48_notexitcond546_pop48_inputs_ready = 1'b1;
assign local_bb4_notexitcond546_push48_notexitcond546_pop48_output_regs_ready = 1'b1;
assign local_bb4_notexitcond546_pop48_c1_ene5_stall_in_0 = 1'b0;
assign local_bb4_c1_ene6_stall_in_0 = 1'b0;
assign SFC_3_VALID_177_177_0_stall_in_2 = 1'b0;
assign local_bb4_notexitcond546_push48_notexitcond546_pop48_causedstall = (SFC_3_VALID_177_177_0 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond546_push48_notexitcond546_pop48_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond546_push48_notexitcond546_pop48_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond546_push48_notexitcond546_pop48_output_regs_ready)
		begin
			local_bb4_notexitcond546_push48_notexitcond546_pop48_NO_SHIFT_REG <= local_bb4_notexitcond546_push48_notexitcond546_pop48_result;
			local_bb4_notexitcond546_push48_notexitcond546_pop48_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond546_push48_notexitcond546_pop48_stall_in))
			begin
				local_bb4_notexitcond546_push48_notexitcond546_pop48_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_notexitcond_or_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb4_notexitcond_or_0_stall_in_NO_SHIFT_REG;
 logic rnode_177to178_bb4_notexitcond_or_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_notexitcond_or_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic rnode_177to178_bb4_notexitcond_or_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_notexitcond_or_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_notexitcond_or_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_notexitcond_or_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_notexitcond_or_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_notexitcond_or_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_notexitcond_or_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_notexitcond_or_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_notexitcond_or_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond_or),
	.data_out(rnode_177to178_bb4_notexitcond_or_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_notexitcond_or_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_notexitcond_or_0_reg_178_fifo.DATA_WIDTH = 1;
defparam rnode_177to178_bb4_notexitcond_or_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_notexitcond_or_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_notexitcond_or_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond_or_stall_in = 1'b0;
assign rnode_177to178_bb4_notexitcond_or_0_NO_SHIFT_REG = rnode_177to178_bb4_notexitcond_or_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_notexitcond_or_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_notexitcond_or_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_stall_local;
wire [31:0] local_bb4_shr_i;

assign local_bb4_shr_i = ((local_bb4_and_i & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i_stall_local;
wire local_bb4_cmp13_i;

assign local_bb4_cmp13_i = ((local_bb4_and10_i & 32'hFFFF) > (local_bb4_and12_i & 32'hFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_forked_and_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to179_bb4_forked_and_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to179_bb4_forked_and_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_forked_and_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to179_bb4_forked_and_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_forked_and_0_valid_out_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_forked_and_0_stall_in_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_forked_and_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_forked_and_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_forked_and_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_forked_and_0_stall_in_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_forked_and_0_valid_out_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_forked_and_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_forked_and_1_NO_SHIFT_REG),
	.data_out(rnode_178to179_bb4_forked_and_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_forked_and_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4_forked_and_0_reg_179_fifo.DATA_WIDTH = 1;
defparam rnode_178to179_bb4_forked_and_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4_forked_and_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4_forked_and_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_forked_and_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_forked_and_0_NO_SHIFT_REG = rnode_178to179_bb4_forked_and_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_forked_and_0_stall_in_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_forked_and_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_178_179_0_inputs_ready;
 reg SFC_3_VALID_178_179_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_178_179_0_stall_in_0;
 reg SFC_3_VALID_178_179_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_178_179_0_stall_in_1;
wire SFC_3_VALID_178_179_0_output_regs_ready;
 reg SFC_3_VALID_178_179_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_178_179_0_causedstall;

assign SFC_3_VALID_178_179_0_inputs_ready = 1'b1;
assign SFC_3_VALID_178_179_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_177_178_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_178_179_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_178_179_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_178_179_0_output_regs_ready)
		begin
			SFC_3_VALID_178_179_0_NO_SHIFT_REG <= SFC_3_VALID_177_178_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_t_34_pop31__valid_out;
wire local_bb4_t_34_pop31__stall_in;
wire local_bb4_t_34_pop31__inputs_ready;
wire local_bb4_t_34_pop31__stall_local;
wire [31:0] local_bb4_t_34_pop31_;
wire local_bb4_t_34_pop31__fu_valid_out;
wire local_bb4_t_34_pop31__fu_stall_out;

acl_pop local_bb4_t_34_pop31__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_177to178_bb4_forked_and_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(32'h0),
	.stall_out(local_bb4_t_34_pop31__fu_stall_out),
	.valid_in(SFC_3_VALID_177_178_0_NO_SHIFT_REG),
	.valid_out(local_bb4_t_34_pop31__fu_valid_out),
	.stall_in(local_bb4_t_34_pop31__stall_local),
	.data_out(local_bb4_t_34_pop31_),
	.feedback_in(feedback_data_in_31),
	.feedback_valid_in(feedback_valid_in_31),
	.feedback_stall_out(feedback_stall_out_31)
);

defparam local_bb4_t_34_pop31__feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_t_34_pop31__feedback.DATA_WIDTH = 32;
defparam local_bb4_t_34_pop31__feedback.STYLE = "REGULAR";

assign local_bb4_t_34_pop31__inputs_ready = (SFC_3_VALID_177_178_0_valid_out_1_NO_SHIFT_REG & rnode_177to178_bb4_forked_and_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_t_34_pop31__stall_local = 1'b0;
assign local_bb4_t_34_pop31__valid_out = 1'b1;
assign SFC_3_VALID_177_178_0_stall_in_1 = 1'b0;
assign rnode_177to178_bb4_forked_and_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond546_push48_notexitcond546_pop48_NO_SHIFT_REG),
	.data_out(rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_fifo.DATA_WIDTH = 1;
defparam rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond546_push48_notexitcond546_pop48_stall_in = 1'b0;
assign rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG = rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 8
//  * capacity = 8
 logic rnode_178to186_bb4_notexitcond_or_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to186_bb4_notexitcond_or_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to186_bb4_notexitcond_or_0_NO_SHIFT_REG;
 logic rnode_178to186_bb4_notexitcond_or_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to186_bb4_notexitcond_or_0_reg_186_NO_SHIFT_REG;
 logic rnode_178to186_bb4_notexitcond_or_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_178to186_bb4_notexitcond_or_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_178to186_bb4_notexitcond_or_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_178to186_bb4_notexitcond_or_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to186_bb4_notexitcond_or_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to186_bb4_notexitcond_or_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_178to186_bb4_notexitcond_or_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_178to186_bb4_notexitcond_or_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_notexitcond_or_0_NO_SHIFT_REG),
	.data_out(rnode_178to186_bb4_notexitcond_or_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_178to186_bb4_notexitcond_or_0_reg_186_fifo.DEPTH = 8;
defparam rnode_178to186_bb4_notexitcond_or_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_178to186_bb4_notexitcond_or_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to186_bb4_notexitcond_or_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_178to186_bb4_notexitcond_or_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_notexitcond_or_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to186_bb4_notexitcond_or_0_NO_SHIFT_REG = rnode_178to186_bb4_notexitcond_or_0_reg_186_NO_SHIFT_REG;
assign rnode_178to186_bb4_notexitcond_or_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_178to186_bb4_notexitcond_or_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i_stall_local;
wire local_bb4_cmp_i;

assign local_bb4_cmp_i = ((local_bb4_shr_i & 32'h7FFF) > (local_bb4_shr3_i & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i_stall_local;
wire local_bb4_cmp8_i;

assign local_bb4_cmp8_i = ((local_bb4_shr_i & 32'h7FFF) == (local_bb4_shr3_i & 32'h7FFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_179_180_0_inputs_ready;
 reg SFC_3_VALID_179_180_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_179_180_0_stall_in;
wire SFC_3_VALID_179_180_0_output_regs_ready;
 reg SFC_3_VALID_179_180_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_179_180_0_causedstall;

assign SFC_3_VALID_179_180_0_inputs_ready = 1'b1;
assign SFC_3_VALID_179_180_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_178_179_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_179_180_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_179_180_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_179_180_0_output_regs_ready)
		begin
			SFC_3_VALID_179_180_0_NO_SHIFT_REG <= SFC_3_VALID_178_179_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_sum_33_pop32__stall_local;
wire [31:0] local_bb4_sum_33_pop32_;
wire local_bb4_sum_33_pop32__fu_valid_out;
wire local_bb4_sum_33_pop32__fu_stall_out;

acl_pop local_bb4_sum_33_pop32__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_178to179_bb4_forked_and_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(32'h0),
	.stall_out(local_bb4_sum_33_pop32__fu_stall_out),
	.valid_in(SFC_3_VALID_178_179_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sum_33_pop32__fu_valid_out),
	.stall_in(local_bb4_sum_33_pop32__stall_local),
	.data_out(local_bb4_sum_33_pop32_),
	.feedback_in(feedback_data_in_32),
	.feedback_valid_in(feedback_valid_in_32),
	.feedback_stall_out(feedback_stall_out_32)
);

defparam local_bb4_sum_33_pop32__feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_sum_33_pop32__feedback.DATA_WIDTH = 32;
defparam local_bb4_sum_33_pop32__feedback.STYLE = "REGULAR";

assign local_bb4_sum_33_pop32__stall_local = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_t_34_pop31__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_t_34_pop31__0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_t_34_pop31__0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_t_34_pop31__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_t_34_pop31__0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_t_34_pop31__1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_t_34_pop31__0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_t_34_pop31__0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_t_34_pop31__0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_t_34_pop31__0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_t_34_pop31__0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_t_34_pop31__0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_t_34_pop31__0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_t_34_pop31__0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_t_34_pop31__0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_t_34_pop31__0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4_t_34_pop31_),
	.data_out(rnode_178to179_bb4_t_34_pop31__0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_t_34_pop31__0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4_t_34_pop31__0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb4_t_34_pop31__0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4_t_34_pop31__0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4_t_34_pop31__0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_t_34_pop31__stall_in = 1'b0;
assign rnode_178to179_bb4_t_34_pop31__0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_t_34_pop31__0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_t_34_pop31__0_NO_SHIFT_REG = rnode_178to179_bb4_t_34_pop31__0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_t_34_pop31__0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_t_34_pop31__1_NO_SHIFT_REG = rnode_178to179_bb4_t_34_pop31__0_reg_179_NO_SHIFT_REG;

// Register node:
//  * latency = 8
//  * capacity = 8
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_NO_SHIFT_REG;
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG;
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_NO_SHIFT_REG;
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG),
	.data_out(rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_fifo.DEPTH = 8;
defparam rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_fifo.DATA_WIDTH = 1;
defparam rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG = rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_187_NO_SHIFT_REG;
assign rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb4_notexitcond_or_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_1_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_notexitcond_or_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb4_notexitcond_or_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb4_notexitcond_or_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb4_notexitcond_or_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb4_notexitcond_or_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb4_notexitcond_or_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(rnode_178to186_bb4_notexitcond_or_0_NO_SHIFT_REG),
	.data_out(rnode_186to187_bb4_notexitcond_or_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb4_notexitcond_or_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb4_notexitcond_or_0_reg_187_fifo.DATA_WIDTH = 1;
defparam rnode_186to187_bb4_notexitcond_or_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb4_notexitcond_or_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb4_notexitcond_or_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to186_bb4_notexitcond_or_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_notexitcond_or_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_notexitcond_or_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb4_notexitcond_or_0_NO_SHIFT_REG = rnode_186to187_bb4_notexitcond_or_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb4_notexitcond_or_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb4_notexitcond_or_1_NO_SHIFT_REG = rnode_186to187_bb4_notexitcond_or_0_reg_187_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4___i_stall_local;
wire local_bb4___i;

assign local_bb4___i = (local_bb4_cmp8_i & local_bb4_cmp13_i);

// This section implements a registered operation.
// 
wire SFC_3_VALID_180_181_0_inputs_ready;
 reg SFC_3_VALID_180_181_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_180_181_0_stall_in;
wire SFC_3_VALID_180_181_0_output_regs_ready;
 reg SFC_3_VALID_180_181_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_180_181_0_causedstall;

assign SFC_3_VALID_180_181_0_inputs_ready = 1'b1;
assign SFC_3_VALID_180_181_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_179_180_0_stall_in = 1'b0;
assign SFC_3_VALID_180_181_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_180_181_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_180_181_0_output_regs_ready)
		begin
			SFC_3_VALID_180_181_0_NO_SHIFT_REG <= SFC_3_VALID_179_180_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u26_stall_local;
wire [31:0] local_bb4_var__u26;

assign local_bb4_var__u26 = local_bb4_sum_33_pop32_;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u27_stall_local;
wire [31:0] local_bb4_var__u27;

assign local_bb4_var__u27 = rnode_178to179_bb4_t_34_pop31__0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_t_34_pop31__0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_t_34_pop31__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_t_34_pop31__0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_t_34_pop31__0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_t_34_pop31__0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_t_34_pop31__0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_t_34_pop31__0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_t_34_pop31__0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_t_34_pop31__0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_t_34_pop31__0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_t_34_pop31__0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_t_34_pop31__0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_t_34_pop31__0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(rnode_178to179_bb4_t_34_pop31__1_NO_SHIFT_REG),
	.data_out(rnode_179to180_bb4_t_34_pop31__0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_t_34_pop31__0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_t_34_pop31__0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_t_34_pop31__0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_t_34_pop31__0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_t_34_pop31__0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_t_34_pop31__0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_t_34_pop31__0_NO_SHIFT_REG = rnode_179to180_bb4_t_34_pop31__0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_t_34_pop31__0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_t_34_pop31__0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_NO_SHIFT_REG;
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG;
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG),
	.data_out(rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_fifo.DATA_WIDTH = 1;
defparam rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to187_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_NO_SHIFT_REG = rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene3_valid_out_1;
wire local_bb4_c1_ene3_stall_in_1;
wire local_bb4_var__u24_valid_out_2;
wire local_bb4_var__u24_stall_in_2;
wire local_bb4_xor_i_valid_out_2;
wire local_bb4_xor_i_stall_in_2;
wire local_bb4__21_i_valid_out;
wire local_bb4__21_i_stall_in;
wire local_bb4__21_i_inputs_ready;
wire local_bb4__21_i_stall_local;
wire local_bb4__21_i;

assign local_bb4__21_i_inputs_ready = (local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG);
assign local_bb4__21_i = (local_bb4_cmp_i | local_bb4___i);
assign local_bb4_c1_ene3_valid_out_1 = 1'b1;
assign local_bb4_var__u24_valid_out_2 = 1'b1;
assign local_bb4_xor_i_valid_out_2 = 1'b1;
assign local_bb4__21_i_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_2 = 1'b0;
assign local_bb4_c1_enter_c1_eni6_stall_in_3 = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_181_182_0_inputs_ready;
 reg SFC_3_VALID_181_182_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_181_182_0_stall_in;
wire SFC_3_VALID_181_182_0_output_regs_ready;
 reg SFC_3_VALID_181_182_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_181_182_0_causedstall;

assign SFC_3_VALID_181_182_0_inputs_ready = 1'b1;
assign SFC_3_VALID_181_182_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_180_181_0_stall_in = 1'b0;
assign SFC_3_VALID_181_182_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_181_182_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_181_182_0_output_regs_ready)
		begin
			SFC_3_VALID_181_182_0_NO_SHIFT_REG <= SFC_3_VALID_180_181_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i99_stall_local;
wire [31:0] local_bb4_shr3_i99;

assign local_bb4_shr3_i99 = (local_bb4_var__u26 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and2_i4_stall_local;
wire [31:0] local_bb4_and2_i4;

assign local_bb4_and2_i4 = (local_bb4_var__u27 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i9_stall_local;
wire [31:0] local_bb4_and12_i9;

assign local_bb4_and12_i9 = (local_bb4_var__u27 & 32'hFFFF);

// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_180to186_bb4_t_34_pop31__0_valid_out_NO_SHIFT_REG;
 logic rnode_180to186_bb4_t_34_pop31__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to186_bb4_t_34_pop31__0_NO_SHIFT_REG;
 logic rnode_180to186_bb4_t_34_pop31__0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to186_bb4_t_34_pop31__0_reg_186_NO_SHIFT_REG;
 logic rnode_180to186_bb4_t_34_pop31__0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_180to186_bb4_t_34_pop31__0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_180to186_bb4_t_34_pop31__0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_180to186_bb4_t_34_pop31__0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to186_bb4_t_34_pop31__0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to186_bb4_t_34_pop31__0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_180to186_bb4_t_34_pop31__0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_180to186_bb4_t_34_pop31__0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_179to180_bb4_t_34_pop31__0_NO_SHIFT_REG),
	.data_out(rnode_180to186_bb4_t_34_pop31__0_reg_186_NO_SHIFT_REG)
);

defparam rnode_180to186_bb4_t_34_pop31__0_reg_186_fifo.DEPTH = 6;
defparam rnode_180to186_bb4_t_34_pop31__0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_180to186_bb4_t_34_pop31__0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to186_bb4_t_34_pop31__0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_180to186_bb4_t_34_pop31__0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_t_34_pop31__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to186_bb4_t_34_pop31__0_NO_SHIFT_REG = rnode_180to186_bb4_t_34_pop31__0_reg_186_NO_SHIFT_REG;
assign rnode_180to186_bb4_t_34_pop31__0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_180to186_bb4_t_34_pop31__0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_177to179_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to179_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to179_bb4_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_177to179_bb4_c1_ene3_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to179_bb4_c1_ene3_0_reg_179_NO_SHIFT_REG;
 logic rnode_177to179_bb4_c1_ene3_0_valid_out_reg_179_NO_SHIFT_REG;
 logic rnode_177to179_bb4_c1_ene3_0_stall_in_reg_179_NO_SHIFT_REG;
 logic rnode_177to179_bb4_c1_ene3_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_177to179_bb4_c1_ene3_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to179_bb4_c1_ene3_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to179_bb4_c1_ene3_0_stall_in_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_177to179_bb4_c1_ene3_0_valid_out_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_177to179_bb4_c1_ene3_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene3),
	.data_out(rnode_177to179_bb4_c1_ene3_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_177to179_bb4_c1_ene3_0_reg_179_fifo.DEPTH = 2;
defparam rnode_177to179_bb4_c1_ene3_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_177to179_bb4_c1_ene3_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to179_bb4_c1_ene3_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_177to179_bb4_c1_ene3_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene3_stall_in_1 = 1'b0;
assign rnode_177to179_bb4_c1_ene3_0_NO_SHIFT_REG = rnode_177to179_bb4_c1_ene3_0_reg_179_NO_SHIFT_REG;
assign rnode_177to179_bb4_c1_ene3_0_stall_in_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_177to179_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_var__u24_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u24_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_var__u24_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u24_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u24_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_var__u24_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u24_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_var__u24_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u24_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u24_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u24_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_var__u24_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_var__u24_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_var__u24_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_var__u24_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_var__u24_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_var__u24),
	.data_out(rnode_177to178_bb4_var__u24_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_var__u24_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_var__u24_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_var__u24_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_var__u24_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_var__u24_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u24_stall_in_2 = 1'b0;
assign rnode_177to178_bb4_var__u24_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_var__u24_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_var__u24_0_NO_SHIFT_REG = rnode_177to178_bb4_var__u24_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_var__u24_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_var__u24_1_NO_SHIFT_REG = rnode_177to178_bb4_var__u24_0_reg_178_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_xor_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_xor_i_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_xor_i_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_xor_i_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_xor_i_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_xor_i_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_xor_i_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_xor_i_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_xor_i_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i),
	.data_out(rnode_177to178_bb4_xor_i_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_xor_i_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_xor_i_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_xor_i_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_xor_i_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_xor_i_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i_stall_in_2 = 1'b0;
assign rnode_177to178_bb4_xor_i_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_xor_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_xor_i_0_NO_SHIFT_REG = rnode_177to178_bb4_xor_i_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_xor_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_xor_i_1_NO_SHIFT_REG = rnode_177to178_bb4_xor_i_0_reg_178_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4__21_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4__21_i_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4__21_i_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4__21_i_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4__21_i_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4__21_i_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4__21_i),
	.data_out(rnode_177to178_bb4__21_i_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4__21_i_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4__21_i_0_reg_178_fifo.DATA_WIDTH = 1;
defparam rnode_177to178_bb4__21_i_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4__21_i_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4__21_i_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i_stall_in = 1'b0;
assign rnode_177to178_bb4__21_i_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4__21_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4__21_i_0_NO_SHIFT_REG = rnode_177to178_bb4__21_i_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4__21_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4__21_i_1_NO_SHIFT_REG = rnode_177to178_bb4__21_i_0_reg_178_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_182_183_0_inputs_ready;
 reg SFC_3_VALID_182_183_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_182_183_0_stall_in;
wire SFC_3_VALID_182_183_0_output_regs_ready;
 reg SFC_3_VALID_182_183_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_182_183_0_causedstall;

assign SFC_3_VALID_182_183_0_inputs_ready = 1'b1;
assign SFC_3_VALID_182_183_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_181_182_0_stall_in = 1'b0;
assign SFC_3_VALID_182_183_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_182_183_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_182_183_0_output_regs_ready)
		begin
			SFC_3_VALID_182_183_0_NO_SHIFT_REG <= SFC_3_VALID_181_182_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_sum_33_pop32__valid_out_1;
wire local_bb4_sum_33_pop32__stall_in_1;
wire local_bb4_var__u26_valid_out_1;
wire local_bb4_var__u26_stall_in_1;
wire local_bb4_cmp_i100_valid_out;
wire local_bb4_cmp_i100_stall_in;
wire local_bb4_cmp_i100_inputs_ready;
wire local_bb4_cmp_i100_stall_local;
wire local_bb4_cmp_i100;

assign local_bb4_cmp_i100_inputs_ready = (SFC_3_VALID_178_179_0_valid_out_1_NO_SHIFT_REG & rnode_178to179_bb4_forked_and_0_valid_out_NO_SHIFT_REG);
assign local_bb4_cmp_i100 = ((local_bb4_shr3_i99 & 32'h7F800000) < 32'h3F800000);
assign local_bb4_sum_33_pop32__valid_out_1 = 1'b1;
assign local_bb4_var__u26_valid_out_1 = 1'b1;
assign local_bb4_cmp_i100_valid_out = 1'b1;
assign SFC_3_VALID_178_179_0_stall_in_1 = 1'b0;
assign rnode_178to179_bb4_forked_and_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i5_stall_local;
wire [31:0] local_bb4_shr3_i5;

assign local_bb4_shr3_i5 = ((local_bb4_and2_i4 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb4_t_34_pop31__0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb4_t_34_pop31__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_t_34_pop31__0_NO_SHIFT_REG;
 logic rnode_186to187_bb4_t_34_pop31__0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_t_34_pop31__0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_t_34_pop31__0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_t_34_pop31__0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_t_34_pop31__0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb4_t_34_pop31__0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb4_t_34_pop31__0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb4_t_34_pop31__0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb4_t_34_pop31__0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb4_t_34_pop31__0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(rnode_180to186_bb4_t_34_pop31__0_NO_SHIFT_REG),
	.data_out(rnode_186to187_bb4_t_34_pop31__0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb4_t_34_pop31__0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb4_t_34_pop31__0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb4_t_34_pop31__0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb4_t_34_pop31__0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb4_t_34_pop31__0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to186_bb4_t_34_pop31__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_t_34_pop31__0_NO_SHIFT_REG = rnode_186to187_bb4_t_34_pop31__0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb4_t_34_pop31__0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_t_34_pop31__0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u28_stall_local;
wire [31:0] local_bb4_var__u28;

assign local_bb4_var__u28 = rnode_177to179_bb4_c1_ene3_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__22_i_stall_local;
wire [31:0] local_bb4__22_i;

assign local_bb4__22_i = (rnode_177to178_bb4__21_i_0_NO_SHIFT_REG ? rnode_177to178_bb4_var__u24_0_NO_SHIFT_REG : rnode_177to178_bb4_xor_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i_stall_local;
wire [31:0] local_bb4__23_i;

assign local_bb4__23_i = (rnode_177to178_bb4__21_i_1_NO_SHIFT_REG ? rnode_177to178_bb4_xor_i_1_NO_SHIFT_REG : rnode_177to178_bb4_var__u24_1_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_3_VALID_183_184_0_inputs_ready;
 reg SFC_3_VALID_183_184_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_183_184_0_stall_in;
wire SFC_3_VALID_183_184_0_output_regs_ready;
 reg SFC_3_VALID_183_184_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_183_184_0_causedstall;

assign SFC_3_VALID_183_184_0_inputs_ready = 1'b1;
assign SFC_3_VALID_183_184_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_182_183_0_stall_in = 1'b0;
assign SFC_3_VALID_183_184_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_183_184_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_183_184_0_output_regs_ready)
		begin
			SFC_3_VALID_183_184_0_NO_SHIFT_REG <= SFC_3_VALID_182_183_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_sum_33_pop32__0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_sum_33_pop32__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_sum_33_pop32__0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_sum_33_pop32__0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_sum_33_pop32__0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_sum_33_pop32__0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_sum_33_pop32__0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_sum_33_pop32__0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_sum_33_pop32__0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_sum_33_pop32__0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_sum_33_pop32__0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_sum_33_pop32__0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_sum_33_pop32__0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_sum_33_pop32_),
	.data_out(rnode_179to180_bb4_sum_33_pop32__0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_sum_33_pop32__0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_sum_33_pop32__0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_sum_33_pop32__0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_sum_33_pop32__0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_sum_33_pop32__0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_sum_33_pop32__stall_in_1 = 1'b0;
assign rnode_179to180_bb4_sum_33_pop32__0_NO_SHIFT_REG = rnode_179to180_bb4_sum_33_pop32__0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_sum_33_pop32__0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_sum_33_pop32__0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_var__u26_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u26_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u26_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u26_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u26_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u26_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u26_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u26_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u26_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u26_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u26_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_var__u26_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_var__u26_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_var__u26_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_var__u26_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_var__u26_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_var__u26),
	.data_out(rnode_179to180_bb4_var__u26_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_var__u26_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_var__u26_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_var__u26_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_var__u26_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_var__u26_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u26_stall_in_1 = 1'b0;
assign rnode_179to180_bb4_var__u26_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u26_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_var__u26_0_NO_SHIFT_REG = rnode_179to180_bb4_var__u26_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_var__u26_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_var__u26_1_NO_SHIFT_REG = rnode_179to180_bb4_var__u26_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_cmp_i100_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp_i100_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_cmp_i100_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_cmp_i100_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_cmp_i100_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_cmp_i100_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_cmp_i100_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_cmp_i100),
	.data_out(rnode_179to180_bb4_cmp_i100_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_cmp_i100_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_cmp_i100_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb4_cmp_i100_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_cmp_i100_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_cmp_i100_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp_i100_stall_in = 1'b0;
assign rnode_179to180_bb4_cmp_i100_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_cmp_i100_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp_i100_0_NO_SHIFT_REG = rnode_179to180_bb4_cmp_i100_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_cmp_i100_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp_i100_1_NO_SHIFT_REG = rnode_179to180_bb4_cmp_i100_0_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i2_stall_local;
wire [31:0] local_bb4_and_i2;

assign local_bb4_and_i2 = (local_bb4_var__u28 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i8_stall_local;
wire [31:0] local_bb4_and10_i8;

assign local_bb4_and10_i8 = (local_bb4_var__u28 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i_stall_local;
wire [31:0] local_bb4_shr18_i;

assign local_bb4_shr18_i = (local_bb4__22_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i_stall_local;
wire [31:0] local_bb4_shr16_i;

assign local_bb4_shr16_i = (local_bb4__23_i >> 32'h17);

// This section implements a registered operation.
// 
wire SFC_3_VALID_184_185_0_inputs_ready;
 reg SFC_3_VALID_184_185_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_184_185_0_stall_in;
wire SFC_3_VALID_184_185_0_output_regs_ready;
 reg SFC_3_VALID_184_185_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_184_185_0_causedstall;

assign SFC_3_VALID_184_185_0_inputs_ready = 1'b1;
assign SFC_3_VALID_184_185_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_183_184_0_stall_in = 1'b0;
assign SFC_3_VALID_184_185_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_184_185_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_184_185_0_output_regs_ready)
		begin
			SFC_3_VALID_184_185_0_NO_SHIFT_REG <= SFC_3_VALID_183_184_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_180to186_bb4_sum_33_pop32__0_valid_out_NO_SHIFT_REG;
 logic rnode_180to186_bb4_sum_33_pop32__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to186_bb4_sum_33_pop32__0_NO_SHIFT_REG;
 logic rnode_180to186_bb4_sum_33_pop32__0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to186_bb4_sum_33_pop32__0_reg_186_NO_SHIFT_REG;
 logic rnode_180to186_bb4_sum_33_pop32__0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_180to186_bb4_sum_33_pop32__0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_180to186_bb4_sum_33_pop32__0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_180to186_bb4_sum_33_pop32__0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to186_bb4_sum_33_pop32__0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to186_bb4_sum_33_pop32__0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_180to186_bb4_sum_33_pop32__0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_180to186_bb4_sum_33_pop32__0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_179to180_bb4_sum_33_pop32__0_NO_SHIFT_REG),
	.data_out(rnode_180to186_bb4_sum_33_pop32__0_reg_186_NO_SHIFT_REG)
);

defparam rnode_180to186_bb4_sum_33_pop32__0_reg_186_fifo.DEPTH = 6;
defparam rnode_180to186_bb4_sum_33_pop32__0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_180to186_bb4_sum_33_pop32__0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to186_bb4_sum_33_pop32__0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_180to186_bb4_sum_33_pop32__0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_sum_33_pop32__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to186_bb4_sum_33_pop32__0_NO_SHIFT_REG = rnode_180to186_bb4_sum_33_pop32__0_reg_186_NO_SHIFT_REG;
assign rnode_180to186_bb4_sum_33_pop32__0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_180to186_bb4_sum_33_pop32__0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__22_i106_stall_local;
wire [31:0] local_bb4__22_i106;

assign local_bb4__22_i106 = (rnode_179to180_bb4_cmp_i100_0_NO_SHIFT_REG ? rnode_179to180_bb4_var__u26_0_NO_SHIFT_REG : 32'h3F800000);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i107_stall_local;
wire [31:0] local_bb4__23_i107;

assign local_bb4__23_i107 = (rnode_179to180_bb4_cmp_i100_1_NO_SHIFT_REG ? 32'h3F800000 : rnode_179to180_bb4_var__u26_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i3_stall_local;
wire [31:0] local_bb4_shr_i3;

assign local_bb4_shr_i3 = ((local_bb4_and_i2 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i10_stall_local;
wire local_bb4_cmp13_i10;

assign local_bb4_cmp13_i10 = ((local_bb4_and10_i8 & 32'hFFFF) > (local_bb4_and12_i9 & 32'hFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i_stall_local;
wire [31:0] local_bb4_and19_i;

assign local_bb4_and19_i = ((local_bb4_shr18_i & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i_stall_local;
wire [31:0] local_bb4_sub_i;

assign local_bb4_sub_i = ((local_bb4_shr16_i & 32'h1FF) - (local_bb4_shr18_i & 32'h1FF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_185_186_0_inputs_ready;
 reg SFC_3_VALID_185_186_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_185_186_0_stall_in;
wire SFC_3_VALID_185_186_0_output_regs_ready;
 reg SFC_3_VALID_185_186_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_185_186_0_causedstall;

assign SFC_3_VALID_185_186_0_inputs_ready = 1'b1;
assign SFC_3_VALID_185_186_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_184_185_0_stall_in = 1'b0;
assign SFC_3_VALID_185_186_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_185_186_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_185_186_0_output_regs_ready)
		begin
			SFC_3_VALID_185_186_0_NO_SHIFT_REG <= SFC_3_VALID_184_185_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb4_sum_33_pop32__0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb4_sum_33_pop32__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_sum_33_pop32__0_NO_SHIFT_REG;
 logic rnode_186to187_bb4_sum_33_pop32__0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_sum_33_pop32__0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_sum_33_pop32__0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_sum_33_pop32__0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_sum_33_pop32__0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb4_sum_33_pop32__0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb4_sum_33_pop32__0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb4_sum_33_pop32__0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb4_sum_33_pop32__0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb4_sum_33_pop32__0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(rnode_180to186_bb4_sum_33_pop32__0_NO_SHIFT_REG),
	.data_out(rnode_186to187_bb4_sum_33_pop32__0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb4_sum_33_pop32__0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb4_sum_33_pop32__0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb4_sum_33_pop32__0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb4_sum_33_pop32__0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb4_sum_33_pop32__0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to186_bb4_sum_33_pop32__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_sum_33_pop32__0_NO_SHIFT_REG = rnode_186to187_bb4_sum_33_pop32__0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb4_sum_33_pop32__0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_sum_33_pop32__0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i110_stall_local;
wire [31:0] local_bb4_shr18_i110;

assign local_bb4_shr18_i110 = (local_bb4__22_i106 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i108_stall_local;
wire [31:0] local_bb4_shr16_i108;

assign local_bb4_shr16_i108 = (local_bb4__23_i107 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i6_stall_local;
wire local_bb4_cmp_i6;

assign local_bb4_cmp_i6 = ((local_bb4_shr_i3 & 32'h7FFF) > (local_bb4_shr3_i5 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i7_stall_local;
wire local_bb4_cmp8_i7;

assign local_bb4_cmp8_i7 = ((local_bb4_shr_i3 & 32'h7FFF) == (local_bb4_shr3_i5 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i_stall_local;
wire local_bb4_lnot23_i;

assign local_bb4_lnot23_i = ((local_bb4_and19_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i_stall_local;
wire local_bb4_cmp27_i;

assign local_bb4_cmp27_i = ((local_bb4_and19_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and69_i_stall_local;
wire [31:0] local_bb4_and69_i;

assign local_bb4_and69_i = (local_bb4_sub_i & 32'hFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_186_187_0_inputs_ready;
 reg SFC_3_VALID_186_187_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_186_187_0_stall_in_0;
 reg SFC_3_VALID_186_187_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_186_187_0_stall_in_1;
 reg SFC_3_VALID_186_187_0_valid_out_2_NO_SHIFT_REG;
wire SFC_3_VALID_186_187_0_stall_in_2;
wire SFC_3_VALID_186_187_0_output_regs_ready;
 reg SFC_3_VALID_186_187_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_186_187_0_causedstall;

assign SFC_3_VALID_186_187_0_inputs_ready = 1'b1;
assign SFC_3_VALID_186_187_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_185_186_0_stall_in = 1'b0;
assign SFC_3_VALID_186_187_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_186_187_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_186_187_0_output_regs_ready)
		begin
			SFC_3_VALID_186_187_0_NO_SHIFT_REG <= SFC_3_VALID_185_186_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and19_i111_stall_local;
wire [31:0] local_bb4_and19_i111;

assign local_bb4_and19_i111 = ((local_bb4_shr18_i110 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i140_stall_local;
wire [31:0] local_bb4_sub_i140;

assign local_bb4_sub_i140 = ((local_bb4_shr16_i108 & 32'h1FF) - (local_bb4_shr18_i110 & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4___i11_stall_local;
wire local_bb4___i11;

assign local_bb4___i11 = (local_bb4_cmp8_i7 & local_bb4_cmp13_i10);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp70_i_stall_local;
wire local_bb4_cmp70_i;

assign local_bb4_cmp70_i = ((local_bb4_and69_i & 32'hFF) > 32'h1F);

// This section implements a registered operation.
// 
wire SFC_3_VALID_187_188_0_inputs_ready;
 reg SFC_3_VALID_187_188_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_187_188_0_stall_in;
wire SFC_3_VALID_187_188_0_output_regs_ready;
 reg SFC_3_VALID_187_188_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_187_188_0_causedstall;

assign SFC_3_VALID_187_188_0_inputs_ready = 1'b1;
assign SFC_3_VALID_187_188_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_186_187_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_187_188_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_187_188_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_187_188_0_output_regs_ready)
		begin
			SFC_3_VALID_187_188_0_NO_SHIFT_REG <= SFC_3_VALID_186_187_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i115_stall_local;
wire local_bb4_lnot23_i115;

assign local_bb4_lnot23_i115 = ((local_bb4_and19_i111 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i117_stall_local;
wire local_bb4_cmp27_i117;

assign local_bb4_cmp27_i117 = ((local_bb4_and19_i111 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and68_i141_stall_local;
wire [31:0] local_bb4_and68_i141;

assign local_bb4_and68_i141 = (local_bb4_sub_i140 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u28_valid_out_2;
wire local_bb4_var__u28_stall_in_2;
wire local_bb4__21_i12_valid_out;
wire local_bb4__21_i12_stall_in;
wire local_bb4_var__u27_valid_out_2;
wire local_bb4_var__u27_stall_in_2;
wire local_bb4__21_i12_inputs_ready;
wire local_bb4__21_i12_stall_local;
wire local_bb4__21_i12;

assign local_bb4__21_i12_inputs_ready = (rnode_177to179_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG & rnode_178to179_bb4_t_34_pop31__0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__21_i12 = (local_bb4_cmp_i6 | local_bb4___i11);
assign local_bb4_var__u28_valid_out_2 = 1'b1;
assign local_bb4__21_i12_valid_out = 1'b1;
assign local_bb4_var__u27_valid_out_2 = 1'b1;
assign rnode_177to179_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_t_34_pop31__0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__22_i_valid_out_1;
wire local_bb4__22_i_stall_in_1;
wire local_bb4__23_i_valid_out_1;
wire local_bb4__23_i_stall_in_1;
wire local_bb4_shr16_i_valid_out_1;
wire local_bb4_shr16_i_stall_in_1;
wire local_bb4_lnot23_i_valid_out;
wire local_bb4_lnot23_i_stall_in;
wire local_bb4_cmp27_i_valid_out;
wire local_bb4_cmp27_i_stall_in;
wire local_bb4_align_0_i_valid_out;
wire local_bb4_align_0_i_stall_in;
wire local_bb4_align_0_i_inputs_ready;
wire local_bb4_align_0_i_stall_local;
wire [31:0] local_bb4_align_0_i;

assign local_bb4_align_0_i_inputs_ready = (rnode_177to178_bb4__21_i_0_valid_out_0_NO_SHIFT_REG & rnode_177to178_bb4_var__u24_0_valid_out_0_NO_SHIFT_REG & rnode_177to178_bb4_xor_i_0_valid_out_0_NO_SHIFT_REG & rnode_177to178_bb4__21_i_0_valid_out_1_NO_SHIFT_REG & rnode_177to178_bb4_xor_i_0_valid_out_1_NO_SHIFT_REG & rnode_177to178_bb4_var__u24_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_align_0_i = (local_bb4_cmp70_i ? 32'h1F : (local_bb4_and69_i & 32'hFF));
assign local_bb4__22_i_valid_out_1 = 1'b1;
assign local_bb4__23_i_valid_out_1 = 1'b1;
assign local_bb4_shr16_i_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i_valid_out = 1'b1;
assign local_bb4_cmp27_i_valid_out = 1'b1;
assign local_bb4_align_0_i_valid_out = 1'b1;
assign rnode_177to178_bb4__21_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_var__u24_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_xor_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4__21_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_xor_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_var__u24_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp69_i142_stall_local;
wire local_bb4_cmp69_i142;

assign local_bb4_cmp69_i142 = ((local_bb4_and68_i141 & 32'hFF) > 32'h1F);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_var__u28_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u28_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u28_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u28_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u28_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u28_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u28_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u28_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u28_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u28_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u28_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_var__u28_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_var__u28_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_var__u28_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_var__u28_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_var__u28_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_var__u28),
	.data_out(rnode_179to180_bb4_var__u28_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_var__u28_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_var__u28_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_var__u28_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_var__u28_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_var__u28_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u28_stall_in_2 = 1'b0;
assign rnode_179to180_bb4_var__u28_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u28_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_var__u28_0_NO_SHIFT_REG = rnode_179to180_bb4_var__u28_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_var__u28_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_var__u28_1_NO_SHIFT_REG = rnode_179to180_bb4_var__u28_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4__21_i12_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4__21_i12_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4__21_i12_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4__21_i12_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4__21_i12_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4__21_i12_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4__21_i12_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4__21_i12),
	.data_out(rnode_179to180_bb4__21_i12_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4__21_i12_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4__21_i12_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb4__21_i12_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4__21_i12_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4__21_i12_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i12_stall_in = 1'b0;
assign rnode_179to180_bb4__21_i12_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4__21_i12_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4__21_i12_0_NO_SHIFT_REG = rnode_179to180_bb4__21_i12_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4__21_i12_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4__21_i12_1_NO_SHIFT_REG = rnode_179to180_bb4__21_i12_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_var__u27_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u27_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u27_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u27_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u27_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u27_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u27_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_var__u27_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u27_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u27_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_var__u27_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_var__u27_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_var__u27_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_var__u27_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_var__u27_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_var__u27_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_var__u27),
	.data_out(rnode_179to180_bb4_var__u27_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_var__u27_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_var__u27_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_var__u27_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_var__u27_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_var__u27_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u27_stall_in_2 = 1'b0;
assign rnode_179to180_bb4_var__u27_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u27_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_var__u27_0_NO_SHIFT_REG = rnode_179to180_bb4_var__u27_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_var__u27_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_var__u27_1_NO_SHIFT_REG = rnode_179to180_bb4_var__u27_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4__22_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__22_i_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__22_i_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__22_i_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4__22_i_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4__22_i_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4__22_i_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4__22_i_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4__22_i_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4__22_i),
	.data_out(rnode_178to179_bb4__22_i_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4__22_i_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4__22_i_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb4__22_i_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4__22_i_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4__22_i_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i_stall_in_1 = 1'b0;
assign rnode_178to179_bb4__22_i_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__22_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__22_i_0_NO_SHIFT_REG = rnode_178to179_bb4__22_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4__22_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__22_i_1_NO_SHIFT_REG = rnode_178to179_bb4__22_i_0_reg_179_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4__23_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4__23_i_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4__23_i_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4__23_i_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4__23_i_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4__23_i_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4__23_i),
	.data_out(rnode_178to179_bb4__23_i_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4__23_i_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4__23_i_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb4__23_i_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4__23_i_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4__23_i_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i_stall_in_1 = 1'b0;
assign rnode_178to179_bb4__23_i_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__23_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__23_i_0_NO_SHIFT_REG = rnode_178to179_bb4__23_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4__23_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__23_i_1_NO_SHIFT_REG = rnode_178to179_bb4__23_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4__23_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__23_i_2_NO_SHIFT_REG = rnode_178to179_bb4__23_i_0_reg_179_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_178to180_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to180_bb4_shr16_i_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to180_bb4_shr16_i_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to180_bb4_shr16_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_178to180_bb4_shr16_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to180_bb4_shr16_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to180_bb4_shr16_i_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_178to180_bb4_shr16_i_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_178to180_bb4_shr16_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i & 32'h1FF)),
	.data_out(rnode_178to180_bb4_shr16_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_178to180_bb4_shr16_i_0_reg_180_fifo.DEPTH = 2;
defparam rnode_178to180_bb4_shr16_i_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_178to180_bb4_shr16_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to180_bb4_shr16_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_178to180_bb4_shr16_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i_stall_in_1 = 1'b0;
assign rnode_178to180_bb4_shr16_i_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_shr16_i_0_NO_SHIFT_REG = rnode_178to180_bb4_shr16_i_0_reg_180_NO_SHIFT_REG;
assign rnode_178to180_bb4_shr16_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_shr16_i_1_NO_SHIFT_REG = rnode_178to180_bb4_shr16_i_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i_0_valid_out_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i_0_stall_in_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_lnot23_i_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_lnot23_i_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_lnot23_i_0_stall_in_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_lnot23_i_0_valid_out_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_lnot23_i_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i),
	.data_out(rnode_178to179_bb4_lnot23_i_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_lnot23_i_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4_lnot23_i_0_reg_179_fifo.DATA_WIDTH = 1;
defparam rnode_178to179_bb4_lnot23_i_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4_lnot23_i_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4_lnot23_i_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i_stall_in = 1'b0;
assign rnode_178to179_bb4_lnot23_i_0_NO_SHIFT_REG = rnode_178to179_bb4_lnot23_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_lnot23_i_0_stall_in_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_178to180_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_2_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_178to180_bb4_cmp27_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to180_bb4_cmp27_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to180_bb4_cmp27_i_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_178to180_bb4_cmp27_i_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_178to180_bb4_cmp27_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i),
	.data_out(rnode_178to180_bb4_cmp27_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_178to180_bb4_cmp27_i_0_reg_180_fifo.DEPTH = 2;
defparam rnode_178to180_bb4_cmp27_i_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_178to180_bb4_cmp27_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to180_bb4_cmp27_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_178to180_bb4_cmp27_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i_stall_in = 1'b0;
assign rnode_178to180_bb4_cmp27_i_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_cmp27_i_0_NO_SHIFT_REG = rnode_178to180_bb4_cmp27_i_0_reg_180_NO_SHIFT_REG;
assign rnode_178to180_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_cmp27_i_1_NO_SHIFT_REG = rnode_178to180_bb4_cmp27_i_0_reg_180_NO_SHIFT_REG;
assign rnode_178to180_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_cmp27_i_2_NO_SHIFT_REG = rnode_178to180_bb4_cmp27_i_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_align_0_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i_3_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i_4_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_align_0_i_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_align_0_i_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_align_0_i_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_align_0_i_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_align_0_i_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in((local_bb4_align_0_i & 32'hFF)),
	.data_out(rnode_178to179_bb4_align_0_i_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_align_0_i_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4_align_0_i_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb4_align_0_i_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4_align_0_i_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4_align_0_i_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_align_0_i_stall_in = 1'b0;
assign rnode_178to179_bb4_align_0_i_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i_0_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i_1_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i_2_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i_3_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i_4_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i_0_reg_179_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_align_0_i143_stall_local;
wire [31:0] local_bb4_align_0_i143;

assign local_bb4_align_0_i143 = (local_bb4_cmp69_i142 ? 32'h1F : (local_bb4_and68_i141 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4__22_i13_stall_local;
wire [31:0] local_bb4__22_i13;

assign local_bb4__22_i13 = (rnode_179to180_bb4__21_i12_0_NO_SHIFT_REG ? rnode_179to180_bb4_var__u27_0_NO_SHIFT_REG : rnode_179to180_bb4_var__u28_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i14_stall_local;
wire [31:0] local_bb4__23_i14;

assign local_bb4__23_i14 = (rnode_179to180_bb4__21_i12_1_NO_SHIFT_REG ? rnode_179to180_bb4_var__u28_1_NO_SHIFT_REG : rnode_179to180_bb4_var__u27_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i_stall_local;
wire [31:0] local_bb4_and21_i;

assign local_bb4_and21_i = (rnode_178to179_bb4__22_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i_valid_out;
wire local_bb4_and20_i_stall_in;
wire local_bb4_and20_i_inputs_ready;
wire local_bb4_and20_i_stall_local;
wire [31:0] local_bb4_and20_i;

assign local_bb4_and20_i_inputs_ready = rnode_178to179_bb4__23_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i = (rnode_178to179_bb4__23_i_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i_valid_out = 1'b1;
assign rnode_178to179_bb4__23_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i_valid_out;
wire local_bb4_and35_i_stall_in;
wire local_bb4_and35_i_inputs_ready;
wire local_bb4_and35_i_stall_local;
wire [31:0] local_bb4_and35_i;

assign local_bb4_and35_i_inputs_ready = rnode_178to179_bb4__23_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i = (rnode_178to179_bb4__23_i_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i_valid_out = 1'b1;
assign rnode_178to179_bb4__23_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor36_i_stall_local;
wire [31:0] local_bb4_xor36_i;

assign local_bb4_xor36_i = (rnode_178to179_bb4__23_i_2_NO_SHIFT_REG ^ rnode_178to179_bb4__22_i_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i_stall_local;
wire [31:0] local_bb4_and17_i;

assign local_bb4_and17_i = ((rnode_178to180_bb4_shr16_i_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_shr16_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_shr16_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_shr16_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_shr16_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_shr16_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_shr16_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((rnode_178to180_bb4_shr16_i_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_180to182_bb4_shr16_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_shr16_i_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_shr16_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_shr16_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_shr16_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_shr16_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_shr16_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_shr16_i_0_NO_SHIFT_REG = rnode_180to182_bb4_shr16_i_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_shr16_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_shr16_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and94_i_stall_local;
wire [31:0] local_bb4_and94_i;

assign local_bb4_and94_i = ((rnode_178to179_bb4_align_0_i_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and96_i_stall_local;
wire [31:0] local_bb4_and96_i;

assign local_bb4_and96_i = ((rnode_178to179_bb4_align_0_i_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and116_i_stall_local;
wire [31:0] local_bb4_and116_i;

assign local_bb4_and116_i = ((rnode_178to179_bb4_align_0_i_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and131_i_stall_local;
wire [31:0] local_bb4_and131_i;

assign local_bb4_and131_i = ((rnode_178to179_bb4_align_0_i_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and150_i_stall_local;
wire [31:0] local_bb4_and150_i;

assign local_bb4_and150_i = ((rnode_178to179_bb4_align_0_i_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and93_i151_stall_local;
wire [31:0] local_bb4_and93_i151;

assign local_bb4_and93_i151 = ((local_bb4_align_0_i143 & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and95_i153_stall_local;
wire [31:0] local_bb4_and95_i153;

assign local_bb4_and95_i153 = ((local_bb4_align_0_i143 & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and115_i169_stall_local;
wire [31:0] local_bb4_and115_i169;

assign local_bb4_and115_i169 = ((local_bb4_align_0_i143 & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and130_i175_stall_local;
wire [31:0] local_bb4_and130_i175;

assign local_bb4_and130_i175 = ((local_bb4_align_0_i143 & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i106_valid_out_1;
wire local_bb4__22_i106_stall_in_1;
wire local_bb4__23_i107_valid_out_1;
wire local_bb4__23_i107_stall_in_1;
wire local_bb4_shr16_i108_valid_out_1;
wire local_bb4_shr16_i108_stall_in_1;
wire local_bb4_lnot23_i115_valid_out;
wire local_bb4_lnot23_i115_stall_in;
wire local_bb4_cmp27_i117_valid_out;
wire local_bb4_cmp27_i117_stall_in;
wire local_bb4_and93_i151_valid_out;
wire local_bb4_and93_i151_stall_in;
wire local_bb4_and95_i153_valid_out;
wire local_bb4_and95_i153_stall_in;
wire local_bb4_and115_i169_valid_out;
wire local_bb4_and115_i169_stall_in;
wire local_bb4_and130_i175_valid_out;
wire local_bb4_and130_i175_stall_in;
wire local_bb4_and149_i180_valid_out;
wire local_bb4_and149_i180_stall_in;
wire local_bb4_and149_i180_inputs_ready;
wire local_bb4_and149_i180_stall_local;
wire [31:0] local_bb4_and149_i180;

assign local_bb4_and149_i180_inputs_ready = (rnode_179to180_bb4_cmp_i100_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb4_var__u26_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb4_cmp_i100_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb4_var__u26_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_and149_i180 = ((local_bb4_align_0_i143 & 32'hFF) & 32'h3);
assign local_bb4__22_i106_valid_out_1 = 1'b1;
assign local_bb4__23_i107_valid_out_1 = 1'b1;
assign local_bb4_shr16_i108_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i115_valid_out = 1'b1;
assign local_bb4_cmp27_i117_valid_out = 1'b1;
assign local_bb4_and93_i151_valid_out = 1'b1;
assign local_bb4_and95_i153_valid_out = 1'b1;
assign local_bb4_and115_i169_valid_out = 1'b1;
assign local_bb4_and130_i175_valid_out = 1'b1;
assign local_bb4_and149_i180_valid_out = 1'b1;
assign rnode_179to180_bb4_cmp_i100_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u26_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_cmp_i100_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u26_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i17_stall_local;
wire [31:0] local_bb4_shr18_i17;

assign local_bb4_shr18_i17 = (local_bb4__22_i13 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i15_stall_local;
wire [31:0] local_bb4_shr16_i15;

assign local_bb4_shr16_i15 = (local_bb4__23_i14 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i_stall_local;
wire local_bb4_lnot33_not_i;

assign local_bb4_lnot33_not_i = ((local_bb4_and21_i & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or65_i_stall_local;
wire [31:0] local_bb4_or65_i;

assign local_bb4_or65_i = ((local_bb4_and21_i & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and20_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and20_i_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and20_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_and20_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_and20_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_and20_i_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_and20_i_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_and20_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i & 32'h7FFFFF)),
	.data_out(rnode_179to180_bb4_and20_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_and20_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_and20_i_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_and20_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_and20_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_and20_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i_stall_in = 1'b0;
assign rnode_179to180_bb4_and20_i_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_and20_i_0_NO_SHIFT_REG = rnode_179to180_bb4_and20_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_and20_i_1_NO_SHIFT_REG = rnode_179to180_bb4_and20_i_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and35_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_and35_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_and35_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_and35_i_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_and35_i_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_and35_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i & 32'h80000000)),
	.data_out(rnode_179to180_bb4_and35_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_and35_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_and35_i_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_and35_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_and35_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_and35_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i_stall_in = 1'b0;
assign rnode_179to180_bb4_and35_i_0_NO_SHIFT_REG = rnode_179to180_bb4_and35_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_and35_i_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp38_i_stall_local;
wire local_bb4_cmp38_i;

assign local_bb4_cmp38_i = ($signed(local_bb4_xor36_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor36_lobit_i_stall_local;
wire [31:0] local_bb4_xor36_lobit_i;

assign local_bb4_xor36_lobit_i = ($signed(local_bb4_xor36_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and37_lobit_i_stall_local;
wire [31:0] local_bb4_and37_lobit_i;

assign local_bb4_and37_lobit_i = (local_bb4_xor36_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i_stall_local;
wire local_bb4_lnot_i;

assign local_bb4_lnot_i = ((local_bb4_and17_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i_stall_local;
wire local_bb4_cmp25_i;

assign local_bb4_cmp25_i = ((local_bb4_and17_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp97_i_stall_local;
wire local_bb4_cmp97_i;

assign local_bb4_cmp97_i = ((local_bb4_and96_i & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp117_i_stall_local;
wire local_bb4_cmp117_i;

assign local_bb4_cmp117_i = ((local_bb4_and116_i & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp132_not_i_stall_local;
wire local_bb4_cmp132_not_i;

assign local_bb4_cmp132_not_i = ((local_bb4_and131_i & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i_stall_local;
wire local_bb4_Pivot20_i;

assign local_bb4_Pivot20_i = ((local_bb4_and150_i & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i_stall_local;
wire local_bb4_SwitchLeaf_i;

assign local_bb4_SwitchLeaf_i = ((local_bb4_and150_i & 32'h3) == 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4__22_i106_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i106_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__22_i106_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i106_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i106_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__22_i106_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i106_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__22_i106_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i106_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i106_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i106_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4__22_i106_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4__22_i106_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4__22_i106_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4__22_i106_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4__22_i106_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4__22_i106),
	.data_out(rnode_180to181_bb4__22_i106_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4__22_i106_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4__22_i106_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4__22_i106_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4__22_i106_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4__22_i106_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i106_stall_in_1 = 1'b0;
assign rnode_180to181_bb4__22_i106_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__22_i106_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__22_i106_0_NO_SHIFT_REG = rnode_180to181_bb4__22_i106_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__22_i106_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__22_i106_1_NO_SHIFT_REG = rnode_180to181_bb4__22_i106_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4__23_i107_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i107_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i107_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i107_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i107_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i107_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4__23_i107_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4__23_i107_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4__23_i107_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4__23_i107_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4__23_i107_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4__23_i107),
	.data_out(rnode_180to181_bb4__23_i107_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4__23_i107_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4__23_i107_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4__23_i107_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4__23_i107_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4__23_i107_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i107_stall_in_1 = 1'b0;
assign rnode_180to181_bb4__23_i107_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__23_i107_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__23_i107_0_NO_SHIFT_REG = rnode_180to181_bb4__23_i107_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__23_i107_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__23_i107_1_NO_SHIFT_REG = rnode_180to181_bb4__23_i107_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__23_i107_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__23_i107_2_NO_SHIFT_REG = rnode_180to181_bb4__23_i107_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_shr16_i108_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i108_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i108_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i108_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i108_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i108_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i108_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i108_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i108_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i108_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i108_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_shr16_i108_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_shr16_i108_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_shr16_i108_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_shr16_i108_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_shr16_i108_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i108 & 32'h1FF)),
	.data_out(rnode_180to182_bb4_shr16_i108_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_shr16_i108_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_shr16_i108_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_shr16_i108_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_shr16_i108_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_shr16_i108_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i108_stall_in_1 = 1'b0;
assign rnode_180to182_bb4_shr16_i108_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_shr16_i108_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_shr16_i108_0_NO_SHIFT_REG = rnode_180to182_bb4_shr16_i108_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_shr16_i108_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_shr16_i108_1_NO_SHIFT_REG = rnode_180to182_bb4_shr16_i108_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_lnot23_i115_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i115_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i115_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i115_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i115_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i115_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i115_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i115_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_lnot23_i115_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_lnot23_i115_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_lnot23_i115_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_lnot23_i115_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_lnot23_i115_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i115),
	.data_out(rnode_180to181_bb4_lnot23_i115_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_lnot23_i115_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_lnot23_i115_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb4_lnot23_i115_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_lnot23_i115_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_lnot23_i115_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i115_stall_in = 1'b0;
assign rnode_180to181_bb4_lnot23_i115_0_NO_SHIFT_REG = rnode_180to181_bb4_lnot23_i115_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_lnot23_i115_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_lnot23_i115_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_cmp27_i117_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i117_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_cmp27_i117_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_cmp27_i117_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_cmp27_i117_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_cmp27_i117_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_cmp27_i117_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i117),
	.data_out(rnode_180to182_bb4_cmp27_i117_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_cmp27_i117_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_cmp27_i117_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_180to182_bb4_cmp27_i117_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_cmp27_i117_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_cmp27_i117_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i117_stall_in = 1'b0;
assign rnode_180to182_bb4_cmp27_i117_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i117_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp27_i117_0_NO_SHIFT_REG = rnode_180to182_bb4_cmp27_i117_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp27_i117_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp27_i117_1_NO_SHIFT_REG = rnode_180to182_bb4_cmp27_i117_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp27_i117_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp27_i117_2_NO_SHIFT_REG = rnode_180to182_bb4_cmp27_i117_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_and93_i151_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and93_i151_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and93_i151_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and93_i151_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and93_i151_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and93_i151_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and93_i151_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and93_i151_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_and93_i151_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_and93_i151_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_and93_i151_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_and93_i151_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_and93_i151_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in((local_bb4_and93_i151 & 32'h1C)),
	.data_out(rnode_180to181_bb4_and93_i151_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_and93_i151_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_and93_i151_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_and93_i151_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_and93_i151_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_and93_i151_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and93_i151_stall_in = 1'b0;
assign rnode_180to181_bb4_and93_i151_0_NO_SHIFT_REG = rnode_180to181_bb4_and93_i151_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_and93_i151_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and93_i151_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_and95_i153_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and95_i153_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and95_i153_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and95_i153_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and95_i153_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and95_i153_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and95_i153_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and95_i153_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_and95_i153_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_and95_i153_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_and95_i153_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_and95_i153_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_and95_i153_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in((local_bb4_and95_i153 & 32'h10)),
	.data_out(rnode_180to181_bb4_and95_i153_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_and95_i153_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_and95_i153_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_and95_i153_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_and95_i153_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_and95_i153_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and95_i153_stall_in = 1'b0;
assign rnode_180to181_bb4_and95_i153_0_NO_SHIFT_REG = rnode_180to181_bb4_and95_i153_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_and95_i153_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and95_i153_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_and115_i169_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and115_i169_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and115_i169_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and115_i169_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and115_i169_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and115_i169_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and115_i169_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and115_i169_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_and115_i169_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_and115_i169_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_and115_i169_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_and115_i169_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_and115_i169_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in((local_bb4_and115_i169 & 32'h8)),
	.data_out(rnode_180to181_bb4_and115_i169_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_and115_i169_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_and115_i169_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_and115_i169_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_and115_i169_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_and115_i169_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and115_i169_stall_in = 1'b0;
assign rnode_180to181_bb4_and115_i169_0_NO_SHIFT_REG = rnode_180to181_bb4_and115_i169_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_and115_i169_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and115_i169_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_and130_i175_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and130_i175_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and130_i175_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and130_i175_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and130_i175_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and130_i175_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and130_i175_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and130_i175_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_and130_i175_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_and130_i175_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_and130_i175_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_and130_i175_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_and130_i175_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in((local_bb4_and130_i175 & 32'h4)),
	.data_out(rnode_180to181_bb4_and130_i175_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_and130_i175_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_and130_i175_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_and130_i175_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_and130_i175_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_and130_i175_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and130_i175_stall_in = 1'b0;
assign rnode_180to181_bb4_and130_i175_0_NO_SHIFT_REG = rnode_180to181_bb4_and130_i175_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_and130_i175_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and130_i175_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_and149_i180_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and149_i180_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and149_i180_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and149_i180_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_and149_i180_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_and149_i180_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_and149_i180_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_and149_i180_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_and149_i180_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_and149_i180_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_and149_i180_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in((local_bb4_and149_i180 & 32'h3)),
	.data_out(rnode_180to181_bb4_and149_i180_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_and149_i180_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_and149_i180_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_and149_i180_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_and149_i180_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_and149_i180_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and149_i180_stall_in = 1'b0;
assign rnode_180to181_bb4_and149_i180_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and149_i180_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_and149_i180_0_NO_SHIFT_REG = rnode_180to181_bb4_and149_i180_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_and149_i180_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_and149_i180_1_NO_SHIFT_REG = rnode_180to181_bb4_and149_i180_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_and149_i180_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_and149_i180_2_NO_SHIFT_REG = rnode_180to181_bb4_and149_i180_0_reg_181_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i18_stall_local;
wire [31:0] local_bb4_and19_i18;

assign local_bb4_and19_i18 = ((local_bb4_shr18_i17 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i44_stall_local;
wire [31:0] local_bb4_sub_i44;

assign local_bb4_sub_i44 = ((local_bb4_shr16_i15 & 32'h1FF) - (local_bb4_shr18_i17 & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl66_i_stall_local;
wire [31:0] local_bb4_shl66_i;

assign local_bb4_shl66_i = ((local_bb4_or65_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i_stall_local;
wire local_bb4_lnot30_i;

assign local_bb4_lnot30_i = ((rnode_179to180_bb4_and20_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_stall_local;
wire [31:0] local_bb4_or_i;

assign local_bb4_or_i = ((rnode_179to180_bb4_and20_i_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and35_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_and35_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_and35_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_and35_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_and35_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_and35_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((rnode_179to180_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_180to182_bb4_and35_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_and35_i_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_and35_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_and35_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_and35_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_and35_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and35_i_0_NO_SHIFT_REG = rnode_180to182_bb4_and35_i_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_and35_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i_stall_local;
wire local_bb4_cmp25_not_i;

assign local_bb4_cmp25_not_i = (local_bb4_cmp25_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u29_stall_local;
wire local_bb4_var__u29;

assign local_bb4_var__u29 = (local_bb4_cmp25_i | rnode_178to180_bb4_cmp27_i_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i113_stall_local;
wire [31:0] local_bb4_and21_i113;

assign local_bb4_and21_i113 = (rnode_180to181_bb4__22_i106_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i112_valid_out;
wire local_bb4_and20_i112_stall_in;
wire local_bb4_and20_i112_inputs_ready;
wire local_bb4_and20_i112_stall_local;
wire [31:0] local_bb4_and20_i112;

assign local_bb4_and20_i112_inputs_ready = rnode_180to181_bb4__23_i107_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i112 = (rnode_180to181_bb4__23_i107_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i112_valid_out = 1'b1;
assign rnode_180to181_bb4__23_i107_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i118_valid_out;
wire local_bb4_and35_i118_stall_in;
wire local_bb4_and35_i118_inputs_ready;
wire local_bb4_and35_i118_stall_local;
wire [31:0] local_bb4_and35_i118;

assign local_bb4_and35_i118_inputs_ready = rnode_180to181_bb4__23_i107_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i118 = (rnode_180to181_bb4__23_i107_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i118_valid_out = 1'b1;
assign rnode_180to181_bb4__23_i107_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i119_stall_local;
wire [31:0] local_bb4_xor_i119;

assign local_bb4_xor_i119 = (rnode_180to181_bb4__23_i107_2_NO_SHIFT_REG ^ rnode_180to181_bb4__22_i106_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i109_stall_local;
wire [31:0] local_bb4_and17_i109;

assign local_bb4_and17_i109 = ((rnode_180to182_bb4_shr16_i108_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_shr16_i108_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i108_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_shr16_i108_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i108_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_shr16_i108_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i108_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i108_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i108_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_shr16_i108_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_shr16_i108_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_shr16_i108_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_shr16_i108_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_shr16_i108_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((rnode_180to182_bb4_shr16_i108_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_182to184_bb4_shr16_i108_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_shr16_i108_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_shr16_i108_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_shr16_i108_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_shr16_i108_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_shr16_i108_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_shr16_i108_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_shr16_i108_0_NO_SHIFT_REG = rnode_182to184_bb4_shr16_i108_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_shr16_i108_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_shr16_i108_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp96_i154_stall_local;
wire local_bb4_cmp96_i154;

assign local_bb4_cmp96_i154 = ((rnode_180to181_bb4_and95_i153_0_NO_SHIFT_REG & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp116_i170_stall_local;
wire local_bb4_cmp116_i170;

assign local_bb4_cmp116_i170 = ((rnode_180to181_bb4_and115_i169_0_NO_SHIFT_REG & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp131_not_i177_stall_local;
wire local_bb4_cmp131_not_i177;

assign local_bb4_cmp131_not_i177 = ((rnode_180to181_bb4_and130_i175_0_NO_SHIFT_REG & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i182_stall_local;
wire local_bb4_Pivot20_i182;

assign local_bb4_Pivot20_i182 = ((rnode_180to181_bb4_and149_i180_1_NO_SHIFT_REG & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i183_stall_local;
wire local_bb4_SwitchLeaf_i183;

assign local_bb4_SwitchLeaf_i183 = ((rnode_180to181_bb4_and149_i180_2_NO_SHIFT_REG & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i22_stall_local;
wire local_bb4_lnot23_i22;

assign local_bb4_lnot23_i22 = ((local_bb4_and19_i18 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i24_stall_local;
wire local_bb4_cmp27_i24;

assign local_bb4_cmp27_i24 = ((local_bb4_and19_i18 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and68_i_stall_local;
wire [31:0] local_bb4_and68_i;

assign local_bb4_and68_i = (local_bb4_sub_i44 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i_stall_local;
wire [31:0] local_bb4__28_i;

assign local_bb4__28_i = (rnode_178to179_bb4_lnot23_i_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl66_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i_stall_local;
wire local_bb4_lnot30_not_i;

assign local_bb4_lnot30_not_i = (local_bb4_lnot30_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_stall_local;
wire [31:0] local_bb4_shl_i;

assign local_bb4_shl_i = ((local_bb4_or_i & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and35_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_and35_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_and35_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_and35_i_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_and35_i_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_and35_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in((rnode_180to182_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_182to183_bb4_and35_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_and35_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_and35_i_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_and35_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_and35_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_and35_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and35_i_0_NO_SHIFT_REG = rnode_182to183_bb4_and35_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_and35_i_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i_stall_local;
wire local_bb4_or_cond_i;

assign local_bb4_or_cond_i = (local_bb4_lnot30_i | local_bb4_cmp25_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i124_stall_local;
wire local_bb4_lnot33_not_i124;

assign local_bb4_lnot33_not_i124 = ((local_bb4_and21_i113 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or64_i137_stall_local;
wire [31:0] local_bb4_or64_i137;

assign local_bb4_or64_i137 = ((local_bb4_and21_i113 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and20_i112_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i112_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and20_i112_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i112_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i112_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and20_i112_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i112_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and20_i112_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i112_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i112_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i112_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and20_i112_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and20_i112_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and20_i112_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and20_i112_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and20_i112_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i112 & 32'h7FFFFF)),
	.data_out(rnode_181to182_bb4_and20_i112_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and20_i112_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and20_i112_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and20_i112_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and20_i112_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and20_i112_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i112_stall_in = 1'b0;
assign rnode_181to182_bb4_and20_i112_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and20_i112_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and20_i112_0_NO_SHIFT_REG = rnode_181to182_bb4_and20_i112_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and20_i112_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and20_i112_1_NO_SHIFT_REG = rnode_181to182_bb4_and20_i112_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and35_i118_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i118_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and35_i118_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i118_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and35_i118_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i118_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i118_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i118_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and35_i118_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and35_i118_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and35_i118_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and35_i118_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and35_i118_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i118 & 32'h80000000)),
	.data_out(rnode_181to182_bb4_and35_i118_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and35_i118_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and35_i118_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and35_i118_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and35_i118_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and35_i118_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i118_stall_in = 1'b0;
assign rnode_181to182_bb4_and35_i118_0_NO_SHIFT_REG = rnode_181to182_bb4_and35_i118_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and35_i118_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and35_i118_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp37_i120_stall_local;
wire local_bb4_cmp37_i120;

assign local_bb4_cmp37_i120 = ($signed(local_bb4_xor_i119) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor_lobit_i193_stall_local;
wire [31:0] local_bb4_xor_lobit_i193;

assign local_bb4_xor_lobit_i193 = ($signed(local_bb4_xor_i119) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and36_lobit_i195_stall_local;
wire [31:0] local_bb4_and36_lobit_i195;

assign local_bb4_and36_lobit_i195 = (local_bb4_xor_i119 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i114_stall_local;
wire local_bb4_lnot_i114;

assign local_bb4_lnot_i114 = ((local_bb4_and17_i109 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i116_stall_local;
wire local_bb4_cmp25_i116;

assign local_bb4_cmp25_i116 = ((local_bb4_and17_i109 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp69_i_stall_local;
wire local_bb4_cmp69_i;

assign local_bb4_cmp69_i = ((local_bb4_and68_i & 32'hFF) > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and73_i_stall_local;
wire [31:0] local_bb4_and73_i;

assign local_bb4_and73_i = ((local_bb4__28_i & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and76_i_stall_local;
wire [31:0] local_bb4_and76_i;

assign local_bb4_and76_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and79_i_stall_local;
wire [31:0] local_bb4_and79_i;

assign local_bb4_and79_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr95_i_stall_local;
wire [31:0] local_bb4_shr95_i;

assign local_bb4_shr95_i = ((local_bb4__28_i & 32'h7FFFFF8) >> (local_bb4_and94_i & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and91_i_stall_local;
wire [31:0] local_bb4_and91_i;

assign local_bb4_and91_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i_stall_local;
wire [31:0] local_bb4_and88_i;

assign local_bb4_and88_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and85_i_stall_local;
wire [31:0] local_bb4_and85_i;

assign local_bb4_and85_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u30_stall_local;
wire [31:0] local_bb4_var__u30;

assign local_bb4_var__u30 = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i_stall_local;
wire local_bb4_or_cond_not_i;

assign local_bb4_or_cond_not_i = (local_bb4_cmp25_i & local_bb4_lnot30_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i_stall_local;
wire [31:0] local_bb4__27_i;

assign local_bb4__27_i = (local_bb4_lnot_i ? 32'h0 : ((local_bb4_shl_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i_stall_local;
wire local_bb4_reduction_8_i;

assign local_bb4_reduction_8_i = (rnode_178to180_bb4_cmp27_i_1_NO_SHIFT_REG & local_bb4_or_cond_i);

// This section implements an unregistered operation.
// 
wire local_bb4_shl65_i138_stall_local;
wire [31:0] local_bb4_shl65_i138;

assign local_bb4_shl65_i138 = ((local_bb4_or64_i137 & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i122_stall_local;
wire local_bb4_lnot30_i122;

assign local_bb4_lnot30_i122 = ((rnode_181to182_bb4_and20_i112_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i134_stall_local;
wire [31:0] local_bb4_or_i134;

assign local_bb4_or_i134 = ((rnode_181to182_bb4_and20_i112_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_and35_i118_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i118_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and35_i118_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i118_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and35_i118_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i118_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i118_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i118_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_and35_i118_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_and35_i118_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_and35_i118_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_and35_i118_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_and35_i118_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((rnode_181to182_bb4_and35_i118_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_182to184_bb4_and35_i118_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_and35_i118_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_and35_i118_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_and35_i118_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_and35_i118_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_and35_i118_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and35_i118_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and35_i118_0_NO_SHIFT_REG = rnode_182to184_bb4_and35_i118_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_and35_i118_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and35_i118_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i121_stall_local;
wire local_bb4_cmp25_not_i121;

assign local_bb4_cmp25_not_i121 = (local_bb4_cmp25_i116 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u31_stall_local;
wire local_bb4_var__u31;

assign local_bb4_var__u31 = (local_bb4_cmp25_i116 | rnode_180to182_bb4_cmp27_i117_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i13_valid_out_1;
wire local_bb4__22_i13_stall_in_1;
wire local_bb4__23_i14_valid_out_1;
wire local_bb4__23_i14_stall_in_1;
wire local_bb4_shr16_i15_valid_out_1;
wire local_bb4_shr16_i15_stall_in_1;
wire local_bb4_lnot23_i22_valid_out;
wire local_bb4_lnot23_i22_stall_in;
wire local_bb4_cmp27_i24_valid_out;
wire local_bb4_cmp27_i24_stall_in;
wire local_bb4_align_0_i45_valid_out;
wire local_bb4_align_0_i45_stall_in;
wire local_bb4_align_0_i45_inputs_ready;
wire local_bb4_align_0_i45_stall_local;
wire [31:0] local_bb4_align_0_i45;

assign local_bb4_align_0_i45_inputs_ready = (rnode_179to180_bb4__21_i12_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb4_var__u27_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb4_var__u28_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb4__21_i12_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb4_var__u28_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb4_var__u27_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_align_0_i45 = (local_bb4_cmp69_i ? 32'h1F : (local_bb4_and68_i & 32'hFF));
assign local_bb4__22_i13_valid_out_1 = 1'b1;
assign local_bb4__23_i14_valid_out_1 = 1'b1;
assign local_bb4_shr16_i15_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i22_valid_out = 1'b1;
assign local_bb4_cmp27_i24_valid_out = 1'b1;
assign local_bb4_align_0_i45_valid_out = 1'b1;
assign rnode_179to180_bb4__21_i12_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u27_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u28_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4__21_i12_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u28_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_var__u27_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and73_tr_i_stall_local;
wire [7:0] local_bb4_and73_tr_i;
wire [31:0] local_bb4_and73_tr_i$ps;

assign local_bb4_and73_tr_i$ps = (local_bb4_and73_i & 32'hFFFFFF);
assign local_bb4_and73_tr_i = local_bb4_and73_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i_stall_local;
wire local_bb4_cmp77_i;

assign local_bb4_cmp77_i = ((local_bb4_and76_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp80_i_stall_local;
wire local_bb4_cmp80_i;

assign local_bb4_cmp80_i = ((local_bb4_and79_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and143_i_stall_local;
wire [31:0] local_bb4_and143_i;

assign local_bb4_and143_i = (local_bb4_shr95_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr151_i_stall_local;
wire [31:0] local_bb4_shr151_i;

assign local_bb4_shr151_i = (local_bb4_shr95_i >> (local_bb4_and150_i & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u32_stall_local;
wire [31:0] local_bb4_var__u32;

assign local_bb4_var__u32 = (local_bb4_shr95_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and147_i_stall_local;
wire [31:0] local_bb4_and147_i;

assign local_bb4_and147_i = (local_bb4_shr95_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp92_i_stall_local;
wire local_bb4_cmp92_i;

assign local_bb4_cmp92_i = ((local_bb4_and91_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp89_i_stall_local;
wire local_bb4_cmp89_i;

assign local_bb4_cmp89_i = ((local_bb4_and88_i & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp86_i_stall_local;
wire local_bb4_cmp86_i;

assign local_bb4_cmp86_i = ((local_bb4_and85_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u33_stall_local;
wire local_bb4_var__u33;

assign local_bb4_var__u33 = ((local_bb4_var__u30 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i139_stall_local;
wire [31:0] local_bb4__28_i139;

assign local_bb4__28_i139 = (rnode_180to181_bb4_lnot23_i115_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl65_i138 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i126_stall_local;
wire local_bb4_lnot30_not_i126;

assign local_bb4_lnot30_not_i126 = (local_bb4_lnot30_i122 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i135_stall_local;
wire [31:0] local_bb4_shl_i135;

assign local_bb4_shl_i135 = ((local_bb4_or_i134 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_and35_i118_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i118_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and35_i118_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i118_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and35_i118_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i118_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i118_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i118_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_and35_i118_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_and35_i118_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_and35_i118_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_and35_i118_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_and35_i118_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in((rnode_182to184_bb4_and35_i118_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_184to185_bb4_and35_i118_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_and35_i118_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_and35_i118_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4_and35_i118_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_and35_i118_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_and35_i118_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_and35_i118_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and35_i118_0_NO_SHIFT_REG = rnode_184to185_bb4_and35_i118_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_and35_i118_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and35_i118_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i123_stall_local;
wire local_bb4_or_cond_i123;

assign local_bb4_or_cond_i123 = (local_bb4_lnot30_i122 | local_bb4_cmp25_not_i121);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4__22_i13_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i13_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__22_i13_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i13_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i13_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__22_i13_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i13_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__22_i13_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i13_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i13_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__22_i13_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4__22_i13_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4__22_i13_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4__22_i13_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4__22_i13_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4__22_i13_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4__22_i13),
	.data_out(rnode_180to181_bb4__22_i13_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4__22_i13_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4__22_i13_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4__22_i13_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4__22_i13_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4__22_i13_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i13_stall_in_1 = 1'b0;
assign rnode_180to181_bb4__22_i13_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__22_i13_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__22_i13_0_NO_SHIFT_REG = rnode_180to181_bb4__22_i13_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__22_i13_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__22_i13_1_NO_SHIFT_REG = rnode_180to181_bb4__22_i13_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4__23_i14_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i14_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i14_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i14_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4__23_i14_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__23_i14_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4__23_i14_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4__23_i14_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4__23_i14_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4__23_i14_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4__23_i14_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4__23_i14),
	.data_out(rnode_180to181_bb4__23_i14_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4__23_i14_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4__23_i14_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4__23_i14_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4__23_i14_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4__23_i14_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i14_stall_in_1 = 1'b0;
assign rnode_180to181_bb4__23_i14_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__23_i14_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__23_i14_0_NO_SHIFT_REG = rnode_180to181_bb4__23_i14_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__23_i14_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__23_i14_1_NO_SHIFT_REG = rnode_180to181_bb4__23_i14_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__23_i14_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__23_i14_2_NO_SHIFT_REG = rnode_180to181_bb4__23_i14_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_shr16_i15_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i15_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i15_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i15_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i15_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i15_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i15_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i15_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i15_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i15_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i15_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_shr16_i15_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_shr16_i15_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_shr16_i15_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_shr16_i15_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_shr16_i15_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i15 & 32'h1FF)),
	.data_out(rnode_180to182_bb4_shr16_i15_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_shr16_i15_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_shr16_i15_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_shr16_i15_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_shr16_i15_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_shr16_i15_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i15_stall_in_1 = 1'b0;
assign rnode_180to182_bb4_shr16_i15_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_shr16_i15_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_shr16_i15_0_NO_SHIFT_REG = rnode_180to182_bb4_shr16_i15_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_shr16_i15_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_shr16_i15_1_NO_SHIFT_REG = rnode_180to182_bb4_shr16_i15_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_lnot23_i22_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i22_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i22_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i22_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i22_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i22_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i22_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_lnot23_i22_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_lnot23_i22_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_lnot23_i22_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_lnot23_i22_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_lnot23_i22_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_lnot23_i22_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i22),
	.data_out(rnode_180to181_bb4_lnot23_i22_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_lnot23_i22_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_lnot23_i22_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb4_lnot23_i22_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_lnot23_i22_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_lnot23_i22_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i22_stall_in = 1'b0;
assign rnode_180to181_bb4_lnot23_i22_0_NO_SHIFT_REG = rnode_180to181_bb4_lnot23_i22_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_lnot23_i22_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_lnot23_i22_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_cmp27_i24_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp27_i24_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_cmp27_i24_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_cmp27_i24_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_cmp27_i24_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_cmp27_i24_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_cmp27_i24_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i24),
	.data_out(rnode_180to182_bb4_cmp27_i24_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_cmp27_i24_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_cmp27_i24_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_180to182_bb4_cmp27_i24_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_cmp27_i24_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_cmp27_i24_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i24_stall_in = 1'b0;
assign rnode_180to182_bb4_cmp27_i24_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i24_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp27_i24_0_NO_SHIFT_REG = rnode_180to182_bb4_cmp27_i24_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp27_i24_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp27_i24_1_NO_SHIFT_REG = rnode_180to182_bb4_cmp27_i24_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp27_i24_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp27_i24_2_NO_SHIFT_REG = rnode_180to182_bb4_cmp27_i24_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_align_0_i45_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_align_0_i45_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_align_0_i45_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_align_0_i45_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_align_0_i45_3_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_align_0_i45_4_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_align_0_i45_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_align_0_i45_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_align_0_i45_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_align_0_i45_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_align_0_i45_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_align_0_i45_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_align_0_i45_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in((local_bb4_align_0_i45 & 32'hFF)),
	.data_out(rnode_180to181_bb4_align_0_i45_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_align_0_i45_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_align_0_i45_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_align_0_i45_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_align_0_i45_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_align_0_i45_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_align_0_i45_stall_in = 1'b0;
assign rnode_180to181_bb4_align_0_i45_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_align_0_i45_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_align_0_i45_0_NO_SHIFT_REG = rnode_180to181_bb4_align_0_i45_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_align_0_i45_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_align_0_i45_1_NO_SHIFT_REG = rnode_180to181_bb4_align_0_i45_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_align_0_i45_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_align_0_i45_2_NO_SHIFT_REG = rnode_180to181_bb4_align_0_i45_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_align_0_i45_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_align_0_i45_3_NO_SHIFT_REG = rnode_180to181_bb4_align_0_i45_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_align_0_i45_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_align_0_i45_4_NO_SHIFT_REG = rnode_180to181_bb4_align_0_i45_0_reg_181_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_frombool75_i_stall_local;
wire [7:0] local_bb4_frombool75_i;

assign local_bb4_frombool75_i = (local_bb4_and73_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u34_stall_local;
wire [31:0] local_bb4_var__u34;

assign local_bb4_var__u34 = ((local_bb4_and147_i & 32'h3FFFFFFF) | local_bb4_shr95_i);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i_stall_local;
wire local_bb4__31_v_i;

assign local_bb4__31_v_i = (local_bb4_cmp97_i ? local_bb4_cmp80_i : local_bb4_cmp92_i);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i_stall_local;
wire local_bb4__30_v_i;

assign local_bb4__30_v_i = (local_bb4_cmp97_i ? local_bb4_cmp77_i : local_bb4_cmp89_i);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool110_i_stall_local;
wire [7:0] local_bb4_frombool110_i;

assign local_bb4_frombool110_i[7:1] = 7'h0;
assign local_bb4_frombool110_i[0] = local_bb4_cmp86_i;

// This section implements an unregistered operation.
// 
wire local_bb4_or108_i_stall_local;
wire [31:0] local_bb4_or108_i;

assign local_bb4_or108_i[31:1] = 31'h0;
assign local_bb4_or108_i[0] = local_bb4_var__u33;

// This section implements an unregistered operation.
// 
wire local_bb4_and72_i144_stall_local;
wire [31:0] local_bb4_and72_i144;

assign local_bb4_and72_i144 = ((local_bb4__28_i139 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i147_stall_local;
wire [31:0] local_bb4_and75_i147;

assign local_bb4_and75_i147 = ((local_bb4__28_i139 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and78_i149_stall_local;
wire [31:0] local_bb4_and78_i149;

assign local_bb4_and78_i149 = ((local_bb4__28_i139 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr94_i152_stall_local;
wire [31:0] local_bb4_shr94_i152;

assign local_bb4_shr94_i152 = ((local_bb4__28_i139 & 32'h7FFFFF8) >> (rnode_180to181_bb4_and93_i151_0_NO_SHIFT_REG & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i155_stall_local;
wire [31:0] local_bb4_and90_i155;

assign local_bb4_and90_i155 = ((local_bb4__28_i139 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and87_i156_stall_local;
wire [31:0] local_bb4_and87_i156;

assign local_bb4_and87_i156 = ((local_bb4__28_i139 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and84_i157_stall_local;
wire [31:0] local_bb4_and84_i157;

assign local_bb4_and84_i157 = ((local_bb4__28_i139 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u35_stall_local;
wire [31:0] local_bb4_var__u35;

assign local_bb4_var__u35 = ((local_bb4__28_i139 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i127_stall_local;
wire local_bb4_or_cond_not_i127;

assign local_bb4_or_cond_not_i127 = (local_bb4_cmp25_i116 & local_bb4_lnot30_not_i126);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i136_stall_local;
wire [31:0] local_bb4__27_i136;

assign local_bb4__27_i136 = (local_bb4_lnot_i114 ? 32'h0 : ((local_bb4_shl_i135 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i131_stall_local;
wire local_bb4_reduction_8_i131;

assign local_bb4_reduction_8_i131 = (rnode_180to182_bb4_cmp27_i117_1_NO_SHIFT_REG & local_bb4_or_cond_i123);

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i20_stall_local;
wire [31:0] local_bb4_and21_i20;

assign local_bb4_and21_i20 = (rnode_180to181_bb4__22_i13_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i19_valid_out;
wire local_bb4_and20_i19_stall_in;
wire local_bb4_and20_i19_inputs_ready;
wire local_bb4_and20_i19_stall_local;
wire [31:0] local_bb4_and20_i19;

assign local_bb4_and20_i19_inputs_ready = rnode_180to181_bb4__23_i14_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i19 = (rnode_180to181_bb4__23_i14_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i19_valid_out = 1'b1;
assign rnode_180to181_bb4__23_i14_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i25_valid_out;
wire local_bb4_and35_i25_stall_in;
wire local_bb4_and35_i25_inputs_ready;
wire local_bb4_and35_i25_stall_local;
wire [31:0] local_bb4_and35_i25;

assign local_bb4_and35_i25_inputs_ready = rnode_180to181_bb4__23_i14_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i25 = (rnode_180to181_bb4__23_i14_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i25_valid_out = 1'b1;
assign rnode_180to181_bb4__23_i14_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i26_stall_local;
wire [31:0] local_bb4_xor_i26;

assign local_bb4_xor_i26 = (rnode_180to181_bb4__23_i14_2_NO_SHIFT_REG ^ rnode_180to181_bb4__22_i13_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i16_stall_local;
wire [31:0] local_bb4_and17_i16;

assign local_bb4_and17_i16 = ((rnode_180to182_bb4_shr16_i15_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_shr16_i15_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i15_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_shr16_i15_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i15_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_shr16_i15_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i15_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i15_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_shr16_i15_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_shr16_i15_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_shr16_i15_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_shr16_i15_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_shr16_i15_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_shr16_i15_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((rnode_180to182_bb4_shr16_i15_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_182to184_bb4_shr16_i15_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_shr16_i15_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_shr16_i15_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_shr16_i15_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_shr16_i15_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_shr16_i15_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_shr16_i15_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_shr16_i15_0_NO_SHIFT_REG = rnode_182to184_bb4_shr16_i15_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_shr16_i15_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_shr16_i15_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and93_i_stall_local;
wire [31:0] local_bb4_and93_i;

assign local_bb4_and93_i = ((rnode_180to181_bb4_align_0_i45_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and95_i_stall_local;
wire [31:0] local_bb4_and95_i;

assign local_bb4_and95_i = ((rnode_180to181_bb4_align_0_i45_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and115_i_stall_local;
wire [31:0] local_bb4_and115_i;

assign local_bb4_and115_i = ((rnode_180to181_bb4_align_0_i45_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and130_i_stall_local;
wire [31:0] local_bb4_and130_i;

assign local_bb4_and130_i = ((rnode_180to181_bb4_align_0_i45_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and149_i_stall_local;
wire [31:0] local_bb4_and149_i;

assign local_bb4_and149_i = ((rnode_180to181_bb4_align_0_i45_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_or1606_i_stall_local;
wire [31:0] local_bb4_or1606_i;

assign local_bb4_or1606_i = (local_bb4_var__u34 | (local_bb4_and143_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i_stall_local;
wire [7:0] local_bb4__31_i;

assign local_bb4__31_i[7:1] = 7'h0;
assign local_bb4__31_i[0] = local_bb4__31_v_i;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i_stall_local;
wire [7:0] local_bb4__30_i;

assign local_bb4__30_i[7:1] = 7'h0;
assign local_bb4__30_i[0] = local_bb4__30_v_i;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i_stall_local;
wire [7:0] local_bb4__29_i;

assign local_bb4__29_i = (local_bb4_cmp97_i ? (local_bb4_frombool75_i & 8'h1) : (local_bb4_frombool110_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i_stall_local;
wire [31:0] local_bb4__32_i;

assign local_bb4__32_i = (local_bb4_cmp97_i ? 32'h0 : (local_bb4_or108_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and72_tr_i145_stall_local;
wire [7:0] local_bb4_and72_tr_i145;
wire [31:0] local_bb4_and72_tr_i145$ps;

assign local_bb4_and72_tr_i145$ps = (local_bb4_and72_i144 & 32'hFFFFFF);
assign local_bb4_and72_tr_i145 = local_bb4_and72_tr_i145$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp76_i148_stall_local;
wire local_bb4_cmp76_i148;

assign local_bb4_cmp76_i148 = ((local_bb4_and75_i147 & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp79_i150_stall_local;
wire local_bb4_cmp79_i150;

assign local_bb4_cmp79_i150 = ((local_bb4_and78_i149 & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and142_i179_stall_local;
wire [31:0] local_bb4_and142_i179;

assign local_bb4_and142_i179 = (local_bb4_shr94_i152 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr150_i181_stall_local;
wire [31:0] local_bb4_shr150_i181;

assign local_bb4_shr150_i181 = (local_bb4_shr94_i152 >> (rnode_180to181_bb4_and149_i180_0_NO_SHIFT_REG & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u36_stall_local;
wire [31:0] local_bb4_var__u36;

assign local_bb4_var__u36 = (local_bb4_shr94_i152 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and146_i184_stall_local;
wire [31:0] local_bb4_and146_i184;

assign local_bb4_and146_i184 = (local_bb4_shr94_i152 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i158_stall_local;
wire local_bb4_cmp91_i158;

assign local_bb4_cmp91_i158 = ((local_bb4_and90_i155 & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp88_i159_stall_local;
wire local_bb4_cmp88_i159;

assign local_bb4_cmp88_i159 = ((local_bb4_and87_i156 & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp85_i160_stall_local;
wire local_bb4_cmp85_i160;

assign local_bb4_cmp85_i160 = ((local_bb4_and84_i157 & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u37_stall_local;
wire local_bb4_var__u37;

assign local_bb4_var__u37 = ((local_bb4_var__u35 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i30_stall_local;
wire local_bb4_lnot33_not_i30;

assign local_bb4_lnot33_not_i30 = ((local_bb4_and21_i20 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or64_i_stall_local;
wire [31:0] local_bb4_or64_i;

assign local_bb4_or64_i = ((local_bb4_and21_i20 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and20_i19_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i19_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and20_i19_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i19_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i19_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and20_i19_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i19_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and20_i19_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i19_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i19_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and20_i19_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and20_i19_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and20_i19_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and20_i19_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and20_i19_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and20_i19_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i19 & 32'h7FFFFF)),
	.data_out(rnode_181to182_bb4_and20_i19_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and20_i19_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and20_i19_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and20_i19_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and20_i19_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and20_i19_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i19_stall_in = 1'b0;
assign rnode_181to182_bb4_and20_i19_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and20_i19_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and20_i19_0_NO_SHIFT_REG = rnode_181to182_bb4_and20_i19_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and20_i19_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and20_i19_1_NO_SHIFT_REG = rnode_181to182_bb4_and20_i19_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and35_i25_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and35_i25_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i25_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and35_i25_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i25_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i25_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and35_i25_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and35_i25_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and35_i25_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and35_i25_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and35_i25_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and35_i25_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i25 & 32'h80000000)),
	.data_out(rnode_181to182_bb4_and35_i25_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and35_i25_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and35_i25_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and35_i25_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and35_i25_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and35_i25_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i25_stall_in = 1'b0;
assign rnode_181to182_bb4_and35_i25_0_NO_SHIFT_REG = rnode_181to182_bb4_and35_i25_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and35_i25_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and35_i25_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp37_i_stall_local;
wire local_bb4_cmp37_i;

assign local_bb4_cmp37_i = ($signed(local_bb4_xor_i26) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor_lobit_i_stall_local;
wire [31:0] local_bb4_xor_lobit_i;

assign local_bb4_xor_lobit_i = ($signed(local_bb4_xor_i26) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and36_lobit_i_stall_local;
wire [31:0] local_bb4_and36_lobit_i;

assign local_bb4_and36_lobit_i = (local_bb4_xor_i26 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i21_stall_local;
wire local_bb4_lnot_i21;

assign local_bb4_lnot_i21 = ((local_bb4_and17_i16 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i23_stall_local;
wire local_bb4_cmp25_i23;

assign local_bb4_cmp25_i23 = ((local_bb4_and17_i16 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp96_i_stall_local;
wire local_bb4_cmp96_i;

assign local_bb4_cmp96_i = ((local_bb4_and95_i & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp116_i_stall_local;
wire local_bb4_cmp116_i;

assign local_bb4_cmp116_i = ((local_bb4_and115_i & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp131_not_i_stall_local;
wire local_bb4_cmp131_not_i;

assign local_bb4_cmp131_not_i = ((local_bb4_and130_i & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i54_stall_local;
wire local_bb4_Pivot20_i54;

assign local_bb4_Pivot20_i54 = ((local_bb4_and149_i & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i55_stall_local;
wire local_bb4_SwitchLeaf_i55;

assign local_bb4_SwitchLeaf_i55 = ((local_bb4_and149_i & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or163_i_stall_local;
wire [31:0] local_bb4_or163_i;

assign local_bb4_or163_i = (local_bb4_or1606_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1247_i_stall_local;
wire [7:0] local_bb4_or1247_i;

assign local_bb4_or1247_i = ((local_bb4__30_i & 8'h1) | (local_bb4__29_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i_stall_local;
wire [7:0] local_bb4__33_i;

assign local_bb4__33_i = (local_bb4_cmp117_i ? (local_bb4__29_i & 8'h1) : (local_bb4__31_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_frombool74_i146_stall_local;
wire [7:0] local_bb4_frombool74_i146;

assign local_bb4_frombool74_i146 = (local_bb4_and72_tr_i145 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u38_stall_local;
wire [31:0] local_bb4_var__u38;

assign local_bb4_var__u38 = ((local_bb4_and146_i184 & 32'h3FFFFFFF) | local_bb4_shr94_i152);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i166_stall_local;
wire local_bb4__31_v_i166;

assign local_bb4__31_v_i166 = (local_bb4_cmp96_i154 ? local_bb4_cmp79_i150 : local_bb4_cmp91_i158);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i164_stall_local;
wire local_bb4__30_v_i164;

assign local_bb4__30_v_i164 = (local_bb4_cmp96_i154 ? local_bb4_cmp76_i148 : local_bb4_cmp88_i159);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool109_i162_stall_local;
wire [7:0] local_bb4_frombool109_i162;

assign local_bb4_frombool109_i162[7:1] = 7'h0;
assign local_bb4_frombool109_i162[0] = local_bb4_cmp85_i160;

// This section implements an unregistered operation.
// 
wire local_bb4_or107_i161_stall_local;
wire [31:0] local_bb4_or107_i161;

assign local_bb4_or107_i161[31:1] = 31'h0;
assign local_bb4_or107_i161[0] = local_bb4_var__u37;

// This section implements an unregistered operation.
// 
wire local_bb4_shl65_i_stall_local;
wire [31:0] local_bb4_shl65_i;

assign local_bb4_shl65_i = ((local_bb4_or64_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i28_stall_local;
wire local_bb4_lnot30_i28;

assign local_bb4_lnot30_i28 = ((rnode_181to182_bb4_and20_i19_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i40_stall_local;
wire [31:0] local_bb4_or_i40;

assign local_bb4_or_i40 = ((rnode_181to182_bb4_and20_i19_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_and35_i25_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and35_i25_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i25_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and35_i25_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i25_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i25_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and35_i25_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_and35_i25_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_and35_i25_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_and35_i25_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_and35_i25_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_and35_i25_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((rnode_181to182_bb4_and35_i25_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_182to184_bb4_and35_i25_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_and35_i25_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_and35_i25_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_and35_i25_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_and35_i25_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_and35_i25_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and35_i25_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and35_i25_0_NO_SHIFT_REG = rnode_182to184_bb4_and35_i25_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_and35_i25_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and35_i25_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i27_stall_local;
wire local_bb4_cmp25_not_i27;

assign local_bb4_cmp25_not_i27 = (local_bb4_cmp25_i23 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u39_stall_local;
wire local_bb4_var__u39;

assign local_bb4_var__u39 = (local_bb4_cmp25_i23 | rnode_180to182_bb4_cmp27_i24_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i_stall_local;
wire [31:0] local_bb4__37_v_i;

assign local_bb4__37_v_i = (local_bb4_Pivot20_i ? 32'h0 : (local_bb4_or163_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i_stall_local;
wire [31:0] local_bb4_or124_i;

assign local_bb4_or124_i[31:8] = 24'h0;
assign local_bb4_or124_i[7:0] = (local_bb4_or1247_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u40_stall_local;
wire [7:0] local_bb4_var__u40;

assign local_bb4_var__u40 = ((local_bb4__33_i & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1596_i185_stall_local;
wire [31:0] local_bb4_or1596_i185;

assign local_bb4_or1596_i185 = (local_bb4_var__u38 | (local_bb4_and142_i179 & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i167_stall_local;
wire [7:0] local_bb4__31_i167;

assign local_bb4__31_i167[7:1] = 7'h0;
assign local_bb4__31_i167[0] = local_bb4__31_v_i166;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i165_stall_local;
wire [7:0] local_bb4__30_i165;

assign local_bb4__30_i165[7:1] = 7'h0;
assign local_bb4__30_i165[0] = local_bb4__30_v_i164;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i163_stall_local;
wire [7:0] local_bb4__29_i163;

assign local_bb4__29_i163 = (local_bb4_cmp96_i154 ? (local_bb4_frombool74_i146 & 8'h1) : (local_bb4_frombool109_i162 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i168_stall_local;
wire [31:0] local_bb4__32_i168;

assign local_bb4__32_i168 = (local_bb4_cmp96_i154 ? 32'h0 : (local_bb4_or107_i161 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__28_i43_stall_local;
wire [31:0] local_bb4__28_i43;

assign local_bb4__28_i43 = (rnode_180to181_bb4_lnot23_i22_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl65_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i32_stall_local;
wire local_bb4_lnot30_not_i32;

assign local_bb4_lnot30_not_i32 = (local_bb4_lnot30_i28 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i41_stall_local;
wire [31:0] local_bb4_shl_i41;

assign local_bb4_shl_i41 = ((local_bb4_or_i40 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_and35_i25_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and35_i25_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i25_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and35_i25_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i25_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i25_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and35_i25_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_and35_i25_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_and35_i25_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_and35_i25_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_and35_i25_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_and35_i25_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in((rnode_182to184_bb4_and35_i25_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_184to185_bb4_and35_i25_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_and35_i25_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_and35_i25_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4_and35_i25_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_and35_i25_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_and35_i25_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_and35_i25_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and35_i25_0_NO_SHIFT_REG = rnode_184to185_bb4_and35_i25_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_and35_i25_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and35_i25_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i29_stall_local;
wire local_bb4_or_cond_i29;

assign local_bb4_or_cond_i29 = (local_bb4_lnot30_i28 | local_bb4_cmp25_not_i27);

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i_stall_local;
wire [31:0] local_bb4__39_v_i;

assign local_bb4__39_v_i = (local_bb4_SwitchLeaf_i ? (local_bb4_var__u32 & 32'h1) : (local_bb4__37_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or125_i_stall_local;
wire [31:0] local_bb4_or125_i;

assign local_bb4_or125_i = (local_bb4_cmp117_i ? 32'h0 : (local_bb4_or124_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv136_i_stall_local;
wire [31:0] local_bb4_conv136_i;

assign local_bb4_conv136_i[31:8] = 24'h0;
assign local_bb4_conv136_i[7:0] = (local_bb4_var__u40 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or162_i186_stall_local;
wire [31:0] local_bb4_or162_i186;

assign local_bb4_or162_i186 = (local_bb4_or1596_i185 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1237_i171_stall_local;
wire [7:0] local_bb4_or1237_i171;

assign local_bb4_or1237_i171 = ((local_bb4__30_i165 & 8'h1) | (local_bb4__29_i163 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i173_stall_local;
wire [7:0] local_bb4__33_i173;

assign local_bb4__33_i173 = (local_bb4_cmp116_i170 ? (local_bb4__29_i163 & 8'h1) : (local_bb4__31_i167 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and72_i_stall_local;
wire [31:0] local_bb4_and72_i;

assign local_bb4_and72_i = ((local_bb4__28_i43 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i_stall_local;
wire [31:0] local_bb4_and75_i;

assign local_bb4_and75_i = ((local_bb4__28_i43 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and78_i_stall_local;
wire [31:0] local_bb4_and78_i;

assign local_bb4_and78_i = ((local_bb4__28_i43 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr94_i_stall_local;
wire [31:0] local_bb4_shr94_i;

assign local_bb4_shr94_i = ((local_bb4__28_i43 & 32'h7FFFFF8) >> (local_bb4_and93_i & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i_stall_local;
wire [31:0] local_bb4_and90_i;

assign local_bb4_and90_i = ((local_bb4__28_i43 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and87_i_stall_local;
wire [31:0] local_bb4_and87_i;

assign local_bb4_and87_i = ((local_bb4__28_i43 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and84_i_stall_local;
wire [31:0] local_bb4_and84_i;

assign local_bb4_and84_i = ((local_bb4__28_i43 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u41_stall_local;
wire [31:0] local_bb4_var__u41;

assign local_bb4_var__u41 = ((local_bb4__28_i43 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i33_stall_local;
wire local_bb4_or_cond_not_i33;

assign local_bb4_or_cond_not_i33 = (local_bb4_cmp25_i23 & local_bb4_lnot30_not_i32);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i42_stall_local;
wire [31:0] local_bb4__27_i42;

assign local_bb4__27_i42 = (local_bb4_lnot_i21 ? 32'h0 : ((local_bb4_shl_i41 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i37_stall_local;
wire local_bb4_reduction_8_i37;

assign local_bb4_reduction_8_i37 = (rnode_180to182_bb4_cmp27_i24_1_NO_SHIFT_REG & local_bb4_or_cond_i29);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i_stall_local;
wire [31:0] local_bb4_reduction_3_i;

assign local_bb4_reduction_3_i = ((local_bb4__32_i & 32'h1) | (local_bb4_or125_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or137_i_stall_local;
wire [31:0] local_bb4_or137_i;

assign local_bb4_or137_i = (local_bb4_cmp132_not_i ? (local_bb4_conv136_i & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i187_stall_local;
wire [31:0] local_bb4__37_v_i187;

assign local_bb4__37_v_i187 = (local_bb4_Pivot20_i182 ? 32'h0 : (local_bb4_or162_i186 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or123_i172_stall_local;
wire [31:0] local_bb4_or123_i172;

assign local_bb4_or123_i172[31:8] = 24'h0;
assign local_bb4_or123_i172[7:0] = (local_bb4_or1237_i171 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u42_stall_local;
wire [7:0] local_bb4_var__u42;

assign local_bb4_var__u42 = ((local_bb4__33_i173 & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and72_tr_i_stall_local;
wire [7:0] local_bb4_and72_tr_i;
wire [31:0] local_bb4_and72_tr_i$ps;

assign local_bb4_and72_tr_i$ps = (local_bb4_and72_i & 32'hFFFFFF);
assign local_bb4_and72_tr_i = local_bb4_and72_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp76_i_stall_local;
wire local_bb4_cmp76_i;

assign local_bb4_cmp76_i = ((local_bb4_and75_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp79_i_stall_local;
wire local_bb4_cmp79_i;

assign local_bb4_cmp79_i = ((local_bb4_and78_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and142_i_stall_local;
wire [31:0] local_bb4_and142_i;

assign local_bb4_and142_i = (local_bb4_shr94_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr150_i_stall_local;
wire [31:0] local_bb4_shr150_i;

assign local_bb4_shr150_i = (local_bb4_shr94_i >> (local_bb4_and149_i & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u43_stall_local;
wire [31:0] local_bb4_var__u43;

assign local_bb4_var__u43 = (local_bb4_shr94_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and146_i_stall_local;
wire [31:0] local_bb4_and146_i;

assign local_bb4_and146_i = (local_bb4_shr94_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i_stall_local;
wire local_bb4_cmp91_i;

assign local_bb4_cmp91_i = ((local_bb4_and90_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp88_i_stall_local;
wire local_bb4_cmp88_i;

assign local_bb4_cmp88_i = ((local_bb4_and87_i & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp85_i_stall_local;
wire local_bb4_cmp85_i;

assign local_bb4_cmp85_i = ((local_bb4_and84_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u44_stall_local;
wire local_bb4_var__u44;

assign local_bb4_var__u44 = ((local_bb4_var__u41 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i_stall_local;
wire [31:0] local_bb4_reduction_5_i;

assign local_bb4_reduction_5_i = (local_bb4_shr151_i | (local_bb4_reduction_3_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i_stall_local;
wire [31:0] local_bb4_reduction_4_i;

assign local_bb4_reduction_4_i = ((local_bb4_or137_i & 32'h1) | (local_bb4__39_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i188_stall_local;
wire [31:0] local_bb4__39_v_i188;

assign local_bb4__39_v_i188 = (local_bb4_SwitchLeaf_i183 ? (local_bb4_var__u36 & 32'h1) : (local_bb4__37_v_i187 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i174_stall_local;
wire [31:0] local_bb4_or124_i174;

assign local_bb4_or124_i174 = (local_bb4_cmp116_i170 ? 32'h0 : (local_bb4_or123_i172 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv135_i176_stall_local;
wire [31:0] local_bb4_conv135_i176;

assign local_bb4_conv135_i176[31:8] = 24'h0;
assign local_bb4_conv135_i176[7:0] = (local_bb4_var__u42 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool74_i_stall_local;
wire [7:0] local_bb4_frombool74_i;

assign local_bb4_frombool74_i = (local_bb4_and72_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u45_stall_local;
wire [31:0] local_bb4_var__u45;

assign local_bb4_var__u45 = ((local_bb4_and146_i & 32'h3FFFFFFF) | local_bb4_shr94_i);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i49_stall_local;
wire local_bb4__31_v_i49;

assign local_bb4__31_v_i49 = (local_bb4_cmp96_i ? local_bb4_cmp79_i : local_bb4_cmp91_i);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i47_stall_local;
wire local_bb4__30_v_i47;

assign local_bb4__30_v_i47 = (local_bb4_cmp96_i ? local_bb4_cmp76_i : local_bb4_cmp88_i);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool109_i_stall_local;
wire [7:0] local_bb4_frombool109_i;

assign local_bb4_frombool109_i[7:1] = 7'h0;
assign local_bb4_frombool109_i[0] = local_bb4_cmp85_i;

// This section implements an unregistered operation.
// 
wire local_bb4_or107_i_stall_local;
wire [31:0] local_bb4_or107_i;

assign local_bb4_or107_i[31:1] = 31'h0;
assign local_bb4_or107_i[0] = local_bb4_var__u44;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i_stall_local;
wire [31:0] local_bb4_reduction_6_i;

assign local_bb4_reduction_6_i = ((local_bb4_reduction_4_i & 32'h1) | local_bb4_reduction_5_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i189_stall_local;
wire [31:0] local_bb4_reduction_3_i189;

assign local_bb4_reduction_3_i189 = ((local_bb4__32_i168 & 32'h1) | (local_bb4_or124_i174 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or136_i178_stall_local;
wire [31:0] local_bb4_or136_i178;

assign local_bb4_or136_i178 = (local_bb4_cmp131_not_i177 ? (local_bb4_conv135_i176 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or1596_i_stall_local;
wire [31:0] local_bb4_or1596_i;

assign local_bb4_or1596_i = (local_bb4_var__u45 | (local_bb4_and142_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i50_stall_local;
wire [7:0] local_bb4__31_i50;

assign local_bb4__31_i50[7:1] = 7'h0;
assign local_bb4__31_i50[0] = local_bb4__31_v_i49;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i48_stall_local;
wire [7:0] local_bb4__30_i48;

assign local_bb4__30_i48[7:1] = 7'h0;
assign local_bb4__30_i48[0] = local_bb4__30_v_i47;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i46_stall_local;
wire [7:0] local_bb4__29_i46;

assign local_bb4__29_i46 = (local_bb4_cmp96_i ? (local_bb4_frombool74_i & 8'h1) : (local_bb4_frombool109_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i51_stall_local;
wire [31:0] local_bb4__32_i51;

assign local_bb4__32_i51 = (local_bb4_cmp96_i ? 32'h0 : (local_bb4_or107_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i_valid_out;
wire local_bb4_lnot33_not_i_stall_in;
wire local_bb4_cmp38_i_valid_out;
wire local_bb4_cmp38_i_stall_in;
wire local_bb4_and37_lobit_i_valid_out;
wire local_bb4_and37_lobit_i_stall_in;
wire local_bb4_xor189_i_valid_out;
wire local_bb4_xor189_i_stall_in;
wire local_bb4_xor189_i_inputs_ready;
wire local_bb4_xor189_i_stall_local;
wire [31:0] local_bb4_xor189_i;

assign local_bb4_xor189_i_inputs_ready = (rnode_178to179_bb4__22_i_0_valid_out_0_NO_SHIFT_REG & rnode_178to179_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i_0_valid_out_0_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i_0_valid_out_4_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i_0_valid_out_1_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i_0_valid_out_2_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i_0_valid_out_3_NO_SHIFT_REG & rnode_178to179_bb4__23_i_0_valid_out_2_NO_SHIFT_REG & rnode_178to179_bb4__22_i_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor189_i = (local_bb4_reduction_6_i ^ local_bb4_xor36_lobit_i);
assign local_bb4_lnot33_not_i_valid_out = 1'b1;
assign local_bb4_cmp38_i_valid_out = 1'b1;
assign local_bb4_and37_lobit_i_valid_out = 1'b1;
assign local_bb4_xor189_i_valid_out = 1'b1;
assign rnode_178to179_bb4__22_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_lnot23_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__23_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__22_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i191_stall_local;
wire [31:0] local_bb4_reduction_5_i191;

assign local_bb4_reduction_5_i191 = (local_bb4_shr150_i181 | (local_bb4_reduction_3_i189 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i190_stall_local;
wire [31:0] local_bb4_reduction_4_i190;

assign local_bb4_reduction_4_i190 = ((local_bb4_or136_i178 & 32'h1) | (local_bb4__39_v_i188 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or162_i_stall_local;
wire [31:0] local_bb4_or162_i;

assign local_bb4_or162_i = (local_bb4_or1596_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1237_i_stall_local;
wire [7:0] local_bb4_or1237_i;

assign local_bb4_or1237_i = ((local_bb4__30_i48 & 8'h1) | (local_bb4__29_i46 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i52_stall_local;
wire [7:0] local_bb4__33_i52;

assign local_bb4__33_i52 = (local_bb4_cmp116_i ? (local_bb4__29_i46 & 8'h1) : (local_bb4__31_i50 & 8'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_lnot33_not_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_lnot33_not_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_lnot33_not_i_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_lnot33_not_i_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_lnot33_not_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i),
	.data_out(rnode_179to180_bb4_lnot33_not_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_lnot33_not_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_lnot33_not_i_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb4_lnot33_not_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_lnot33_not_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_lnot33_not_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i_stall_in = 1'b0;
assign rnode_179to180_bb4_lnot33_not_i_0_NO_SHIFT_REG = rnode_179to180_bb4_lnot33_not_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_lnot33_not_i_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_cmp38_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_cmp38_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_cmp38_i_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_cmp38_i_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_cmp38_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_cmp38_i),
	.data_out(rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_cmp38_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp38_i_stall_in = 1'b0;
assign rnode_179to180_bb4_cmp38_i_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp38_i_0_NO_SHIFT_REG = rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp38_i_1_NO_SHIFT_REG = rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and37_lobit_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and37_lobit_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_and37_lobit_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_and37_lobit_i_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_and37_lobit_i_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_and37_lobit_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_and37_lobit_i & 32'h1)),
	.data_out(rnode_179to180_bb4_and37_lobit_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_and37_lobit_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and37_lobit_i_stall_in = 1'b0;
assign rnode_179to180_bb4_and37_lobit_i_0_NO_SHIFT_REG = rnode_179to180_bb4_and37_lobit_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_and37_lobit_i_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_xor189_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_xor189_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_xor189_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_xor189_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_xor189_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_xor189_i_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_xor189_i_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_xor189_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_xor189_i),
	.data_out(rnode_179to180_bb4_xor189_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_xor189_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor189_i_stall_in = 1'b0;
assign rnode_179to180_bb4_xor189_i_0_NO_SHIFT_REG = rnode_179to180_bb4_xor189_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_xor189_i_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_xor189_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i192_stall_local;
wire [31:0] local_bb4_reduction_6_i192;

assign local_bb4_reduction_6_i192 = ((local_bb4_reduction_4_i190 & 32'h1) | local_bb4_reduction_5_i191);

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i56_stall_local;
wire [31:0] local_bb4__37_v_i56;

assign local_bb4__37_v_i56 = (local_bb4_Pivot20_i54 ? 32'h0 : (local_bb4_or162_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or123_i_stall_local;
wire [31:0] local_bb4_or123_i;

assign local_bb4_or123_i[31:8] = 24'h0;
assign local_bb4_or123_i[7:0] = (local_bb4_or1237_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u46_stall_local;
wire [7:0] local_bb4_var__u46;

assign local_bb4_var__u46 = ((local_bb4__33_i52 & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i_stall_local;
wire local_bb4_brmerge_not_i;

assign local_bb4_brmerge_not_i = (rnode_178to180_bb4_cmp27_i_0_NO_SHIFT_REG & rnode_179to180_bb4_lnot33_not_i_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_cmp38_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_cmp38_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_cmp38_i_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_cmp38_i_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_cmp38_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_179to180_bb4_cmp38_i_1_NO_SHIFT_REG),
	.data_out(rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_cmp38_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp38_i_0_NO_SHIFT_REG = rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp38_i_1_NO_SHIFT_REG = rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp38_i_2_NO_SHIFT_REG = rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i_stall_local;
wire [31:0] local_bb4_add_i;

assign local_bb4_add_i = ((local_bb4__27_i & 32'h7FFFFF8) | (rnode_179to180_bb4_and37_lobit_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i124_valid_out;
wire local_bb4_lnot33_not_i124_stall_in;
wire local_bb4_cmp37_i120_valid_out;
wire local_bb4_cmp37_i120_stall_in;
wire local_bb4_and36_lobit_i195_valid_out;
wire local_bb4_and36_lobit_i195_stall_in;
wire local_bb4_xor188_i194_valid_out;
wire local_bb4_xor188_i194_stall_in;
wire local_bb4_xor188_i194_inputs_ready;
wire local_bb4_xor188_i194_stall_local;
wire [31:0] local_bb4_xor188_i194;

assign local_bb4_xor188_i194_inputs_ready = (rnode_180to181_bb4__22_i106_0_valid_out_0_NO_SHIFT_REG & rnode_180to181_bb4_lnot23_i115_0_valid_out_NO_SHIFT_REG & rnode_180to181_bb4_and93_i151_0_valid_out_NO_SHIFT_REG & rnode_180to181_bb4_and149_i180_0_valid_out_0_NO_SHIFT_REG & rnode_180to181_bb4_and95_i153_0_valid_out_NO_SHIFT_REG & rnode_180to181_bb4_and149_i180_0_valid_out_2_NO_SHIFT_REG & rnode_180to181_bb4_and115_i169_0_valid_out_NO_SHIFT_REG & rnode_180to181_bb4_and130_i175_0_valid_out_NO_SHIFT_REG & rnode_180to181_bb4_and149_i180_0_valid_out_1_NO_SHIFT_REG & rnode_180to181_bb4__23_i107_0_valid_out_2_NO_SHIFT_REG & rnode_180to181_bb4__22_i106_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor188_i194 = (local_bb4_reduction_6_i192 ^ local_bb4_xor_lobit_i193);
assign local_bb4_lnot33_not_i124_valid_out = 1'b1;
assign local_bb4_cmp37_i120_valid_out = 1'b1;
assign local_bb4_and36_lobit_i195_valid_out = 1'b1;
assign local_bb4_xor188_i194_valid_out = 1'b1;
assign rnode_180to181_bb4__22_i106_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_lnot23_i115_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and93_i151_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and149_i180_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and95_i153_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and149_i180_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and115_i169_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and130_i175_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_and149_i180_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__23_i107_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__22_i106_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i57_stall_local;
wire [31:0] local_bb4__39_v_i57;

assign local_bb4__39_v_i57 = (local_bb4_SwitchLeaf_i55 ? (local_bb4_var__u43 & 32'h1) : (local_bb4__37_v_i56 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i53_stall_local;
wire [31:0] local_bb4_or124_i53;

assign local_bb4_or124_i53 = (local_bb4_cmp116_i ? 32'h0 : (local_bb4_or123_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv135_i_stall_local;
wire [31:0] local_bb4_conv135_i;

assign local_bb4_conv135_i[31:8] = 24'h0;
assign local_bb4_conv135_i[7:0] = (local_bb4_var__u46 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i_stall_local;
wire local_bb4__24_i;

assign local_bb4__24_i = (local_bb4_or_cond_not_i | local_bb4_brmerge_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i_stall_local;
wire local_bb4_brmerge_not_not_i;

assign local_bb4_brmerge_not_not_i = (local_bb4_brmerge_not_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp38_i_stall_local;
wire local_bb4_not_cmp38_i;

assign local_bb4_not_cmp38_i = (rnode_180to182_bb4_cmp38_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add193_i_stall_local;
wire [31:0] local_bb4_add193_i;

assign local_bb4_add193_i = ((local_bb4_add_i & 32'h7FFFFF9) + rnode_179to180_bb4_xor189_i_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_lnot33_not_i124_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i124_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i124_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i124_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i124_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i124_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i124_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i124_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_lnot33_not_i124_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_lnot33_not_i124_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_lnot33_not_i124_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_lnot33_not_i124_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_lnot33_not_i124_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i124),
	.data_out(rnode_181to182_bb4_lnot33_not_i124_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_lnot33_not_i124_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_lnot33_not_i124_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb4_lnot33_not_i124_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_lnot33_not_i124_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_lnot33_not_i124_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i124_stall_in = 1'b0;
assign rnode_181to182_bb4_lnot33_not_i124_0_NO_SHIFT_REG = rnode_181to182_bb4_lnot33_not_i124_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_lnot33_not_i124_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_lnot33_not_i124_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_cmp37_i120_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i120_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_cmp37_i120_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_cmp37_i120_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_cmp37_i120_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_cmp37_i120_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_cmp37_i120_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_cmp37_i120),
	.data_out(rnode_181to182_bb4_cmp37_i120_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_cmp37_i120_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_cmp37_i120_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb4_cmp37_i120_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_cmp37_i120_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_cmp37_i120_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp37_i120_stall_in = 1'b0;
assign rnode_181to182_bb4_cmp37_i120_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_cmp37_i120_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_cmp37_i120_0_NO_SHIFT_REG = rnode_181to182_bb4_cmp37_i120_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_cmp37_i120_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_cmp37_i120_1_NO_SHIFT_REG = rnode_181to182_bb4_cmp37_i120_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and36_lobit_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and36_lobit_i195_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i195_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and36_lobit_i195_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i195_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i195_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i195_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and36_lobit_i195_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and36_lobit_i195_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and36_lobit_i195_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and36_lobit_i195_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and36_lobit_i195_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and36_lobit_i195 & 32'h1)),
	.data_out(rnode_181to182_bb4_and36_lobit_i195_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and36_lobit_i195_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and36_lobit_i195_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and36_lobit_i195_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and36_lobit_i195_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and36_lobit_i195_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and36_lobit_i195_stall_in = 1'b0;
assign rnode_181to182_bb4_and36_lobit_i195_0_NO_SHIFT_REG = rnode_181to182_bb4_and36_lobit_i195_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and36_lobit_i195_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and36_lobit_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_xor188_i194_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i194_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_xor188_i194_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i194_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_xor188_i194_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i194_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i194_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i194_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_xor188_i194_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_xor188_i194_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_xor188_i194_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_xor188_i194_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_xor188_i194_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_xor188_i194),
	.data_out(rnode_181to182_bb4_xor188_i194_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_xor188_i194_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_xor188_i194_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_xor188_i194_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_xor188_i194_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_xor188_i194_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor188_i194_stall_in = 1'b0;
assign rnode_181to182_bb4_xor188_i194_0_NO_SHIFT_REG = rnode_181to182_bb4_xor188_i194_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_xor188_i194_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_xor188_i194_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i58_stall_local;
wire [31:0] local_bb4_reduction_3_i58;

assign local_bb4_reduction_3_i58 = ((local_bb4__32_i51 & 32'h1) | (local_bb4_or124_i53 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or136_i_stall_local;
wire [31:0] local_bb4_or136_i;

assign local_bb4_or136_i = (local_bb4_cmp131_not_i ? (local_bb4_conv135_i & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i_stall_local;
wire local_bb4_reduction_7_i;

assign local_bb4_reduction_7_i = (local_bb4_cmp25_i & local_bb4_brmerge_not_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i125_stall_local;
wire local_bb4_brmerge_not_i125;

assign local_bb4_brmerge_not_i125 = (rnode_180to182_bb4_cmp27_i117_0_NO_SHIFT_REG & rnode_181to182_bb4_lnot33_not_i124_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_cmp37_i120_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_1_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_2_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i120_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_cmp37_i120_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_cmp37_i120_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_cmp37_i120_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_cmp37_i120_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_cmp37_i120_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb4_cmp37_i120_1_NO_SHIFT_REG),
	.data_out(rnode_182to184_bb4_cmp37_i120_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_cmp37_i120_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_cmp37_i120_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_182to184_bb4_cmp37_i120_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_cmp37_i120_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_cmp37_i120_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_cmp37_i120_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i120_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i120_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_cmp37_i120_0_NO_SHIFT_REG = rnode_182to184_bb4_cmp37_i120_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_cmp37_i120_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_cmp37_i120_1_NO_SHIFT_REG = rnode_182to184_bb4_cmp37_i120_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_cmp37_i120_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_cmp37_i120_2_NO_SHIFT_REG = rnode_182to184_bb4_cmp37_i120_0_reg_184_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i196_stall_local;
wire [31:0] local_bb4_add_i196;

assign local_bb4_add_i196 = ((local_bb4__27_i136 & 32'h7FFFFF8) | (rnode_181to182_bb4_and36_lobit_i195_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i60_stall_local;
wire [31:0] local_bb4_reduction_5_i60;

assign local_bb4_reduction_5_i60 = (local_bb4_shr150_i | (local_bb4_reduction_3_i58 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i59_stall_local;
wire [31:0] local_bb4_reduction_4_i59;

assign local_bb4_reduction_4_i59 = ((local_bb4_or136_i & 32'h1) | (local_bb4__39_v_i57 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i_stall_local;
wire local_bb4_reduction_9_i;

assign local_bb4_reduction_9_i = (local_bb4_reduction_7_i & local_bb4_reduction_8_i);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i128_stall_local;
wire local_bb4__24_i128;

assign local_bb4__24_i128 = (local_bb4_or_cond_not_i127 | local_bb4_brmerge_not_i125);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i129_stall_local;
wire local_bb4_brmerge_not_not_i129;

assign local_bb4_brmerge_not_not_i129 = (local_bb4_brmerge_not_i125 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp37_i226_stall_local;
wire local_bb4_not_cmp37_i226;

assign local_bb4_not_cmp37_i226 = (rnode_182to184_bb4_cmp37_i120_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add192_i197_stall_local;
wire [31:0] local_bb4_add192_i197;

assign local_bb4_add192_i197 = ((local_bb4_add_i196 & 32'h7FFFFF9) + rnode_181to182_bb4_xor188_i194_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i61_stall_local;
wire [31:0] local_bb4_reduction_6_i61;

assign local_bb4_reduction_6_i61 = ((local_bb4_reduction_4_i59 & 32'h1) | local_bb4_reduction_5_i60);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i_valid_out_2;
wire local_bb4_and17_i_stall_in_2;
wire local_bb4_var__u29_valid_out;
wire local_bb4_var__u29_stall_in;
wire local_bb4_add193_i_valid_out;
wire local_bb4_add193_i_stall_in;
wire local_bb4__26_i_valid_out;
wire local_bb4__26_i_stall_in;
wire local_bb4__26_i_inputs_ready;
wire local_bb4__26_i_stall_local;
wire local_bb4__26_i;

assign local_bb4__26_i_inputs_ready = (rnode_178to180_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG & rnode_178to180_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_179to180_bb4_xor189_i_0_valid_out_NO_SHIFT_REG & rnode_179to180_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG & rnode_178to180_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG & rnode_178to180_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i = (local_bb4_reduction_9_i ? rnode_179to180_bb4_cmp38_i_0_NO_SHIFT_REG : local_bb4__24_i);
assign local_bb4_and17_i_valid_out_2 = 1'b1;
assign local_bb4_var__u29_valid_out = 1'b1;
assign local_bb4_add193_i_valid_out = 1'b1;
assign local_bb4__26_i_valid_out = 1'b1;
assign rnode_178to180_bb4_shr16_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and37_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_xor189_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and20_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_lnot33_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and20_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i130_stall_local;
wire local_bb4_reduction_7_i130;

assign local_bb4_reduction_7_i130 = (local_bb4_cmp25_i116 & local_bb4_brmerge_not_not_i129);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i30_valid_out;
wire local_bb4_lnot33_not_i30_stall_in;
wire local_bb4_cmp37_i_valid_out;
wire local_bb4_cmp37_i_stall_in;
wire local_bb4_and36_lobit_i_valid_out;
wire local_bb4_and36_lobit_i_stall_in;
wire local_bb4_xor188_i_valid_out;
wire local_bb4_xor188_i_stall_in;
wire local_bb4_xor188_i_inputs_ready;
wire local_bb4_xor188_i_stall_local;
wire [31:0] local_bb4_xor188_i;

assign local_bb4_xor188_i_inputs_ready = (rnode_180to181_bb4__22_i13_0_valid_out_0_NO_SHIFT_REG & rnode_180to181_bb4_lnot23_i22_0_valid_out_NO_SHIFT_REG & rnode_180to181_bb4_align_0_i45_0_valid_out_0_NO_SHIFT_REG & rnode_180to181_bb4_align_0_i45_0_valid_out_4_NO_SHIFT_REG & rnode_180to181_bb4_align_0_i45_0_valid_out_1_NO_SHIFT_REG & rnode_180to181_bb4_align_0_i45_0_valid_out_2_NO_SHIFT_REG & rnode_180to181_bb4_align_0_i45_0_valid_out_3_NO_SHIFT_REG & rnode_180to181_bb4__23_i14_0_valid_out_2_NO_SHIFT_REG & rnode_180to181_bb4__22_i13_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor188_i = (local_bb4_reduction_6_i61 ^ local_bb4_xor_lobit_i);
assign local_bb4_lnot33_not_i30_valid_out = 1'b1;
assign local_bb4_cmp37_i_valid_out = 1'b1;
assign local_bb4_and36_lobit_i_valid_out = 1'b1;
assign local_bb4_xor188_i_valid_out = 1'b1;
assign rnode_180to181_bb4__22_i13_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_lnot23_i22_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_align_0_i45_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_align_0_i45_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_align_0_i45_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_align_0_i45_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_align_0_i45_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__23_i14_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__22_i13_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_and17_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and17_i_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and17_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_and17_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_and17_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_and17_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_and17_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_and17_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i & 32'hFF)),
	.data_out(rnode_180to182_bb4_and17_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_and17_i_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_and17_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_and17_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_and17_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_and17_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i_stall_in_2 = 1'b0;
assign rnode_180to182_bb4_and17_i_0_NO_SHIFT_REG = rnode_180to182_bb4_and17_i_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_and17_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and17_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_var__u29_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u29_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u29_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u29_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u29_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u29_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u29_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u29_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_var__u29_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_var__u29_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_var__u29_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_var__u29_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_var__u29_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4_var__u29),
	.data_out(rnode_180to181_bb4_var__u29_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_var__u29_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_var__u29_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb4_var__u29_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_var__u29_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_var__u29_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u29_stall_in = 1'b0;
assign rnode_180to181_bb4_var__u29_0_NO_SHIFT_REG = rnode_180to181_bb4_var__u29_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_var__u29_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_var__u29_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_3_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_add193_i_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_add193_i_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_add193_i_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_add193_i_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_add193_i_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4_add193_i),
	.data_out(rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_add193_i_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add193_i_stall_in = 1'b0;
assign rnode_180to181_bb4_add193_i_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_0_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_1_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_2_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_3_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4__26_i_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4__26_i_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4__26_i_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4__26_i_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4__26_i_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4__26_i),
	.data_out(rnode_180to181_bb4__26_i_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4__26_i_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4__26_i_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb4__26_i_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4__26_i_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4__26_i_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i_stall_in = 1'b0;
assign rnode_180to181_bb4__26_i_0_NO_SHIFT_REG = rnode_180to181_bb4__26_i_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__26_i_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i132_stall_local;
wire local_bb4_reduction_9_i132;

assign local_bb4_reduction_9_i132 = (local_bb4_reduction_7_i130 & local_bb4_reduction_8_i131);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_lnot33_not_i30_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i30_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i30_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i30_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i30_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i30_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i30_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_lnot33_not_i30_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_lnot33_not_i30_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_lnot33_not_i30_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_lnot33_not_i30_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_lnot33_not_i30_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_lnot33_not_i30_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i30),
	.data_out(rnode_181to182_bb4_lnot33_not_i30_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_lnot33_not_i30_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_lnot33_not_i30_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb4_lnot33_not_i30_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_lnot33_not_i30_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_lnot33_not_i30_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i30_stall_in = 1'b0;
assign rnode_181to182_bb4_lnot33_not_i30_0_NO_SHIFT_REG = rnode_181to182_bb4_lnot33_not_i30_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_lnot33_not_i30_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_lnot33_not_i30_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_cmp37_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_cmp37_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_cmp37_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_cmp37_i_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_cmp37_i_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_cmp37_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_cmp37_i),
	.data_out(rnode_181to182_bb4_cmp37_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_cmp37_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_cmp37_i_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb4_cmp37_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_cmp37_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_cmp37_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp37_i_stall_in = 1'b0;
assign rnode_181to182_bb4_cmp37_i_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_cmp37_i_0_NO_SHIFT_REG = rnode_181to182_bb4_cmp37_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_cmp37_i_1_NO_SHIFT_REG = rnode_181to182_bb4_cmp37_i_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and36_lobit_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and36_lobit_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and36_lobit_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and36_lobit_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and36_lobit_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and36_lobit_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and36_lobit_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and36_lobit_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and36_lobit_i & 32'h1)),
	.data_out(rnode_181to182_bb4_and36_lobit_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and36_lobit_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and36_lobit_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and36_lobit_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and36_lobit_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and36_lobit_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and36_lobit_i_stall_in = 1'b0;
assign rnode_181to182_bb4_and36_lobit_i_0_NO_SHIFT_REG = rnode_181to182_bb4_and36_lobit_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and36_lobit_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_xor188_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_xor188_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_xor188_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_xor188_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_xor188_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_xor188_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_xor188_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_xor188_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_xor188_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb4_xor188_i),
	.data_out(rnode_181to182_bb4_xor188_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_xor188_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_xor188_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_xor188_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_xor188_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_xor188_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor188_i_stall_in = 1'b0;
assign rnode_181to182_bb4_xor188_i_0_NO_SHIFT_REG = rnode_181to182_bb4_xor188_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_xor188_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_xor188_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_var__u29_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u29_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u29_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u29_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u29_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u29_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u29_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u29_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_var__u29_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_var__u29_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_var__u29_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_var__u29_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_var__u29_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb4_var__u29_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb4_var__u29_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_var__u29_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_var__u29_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb4_var__u29_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_var__u29_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_var__u29_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_var__u29_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_var__u29_0_NO_SHIFT_REG = rnode_181to182_bb4_var__u29_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_var__u29_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_var__u29_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and194_i_valid_out;
wire local_bb4_and194_i_stall_in;
wire local_bb4_and194_i_inputs_ready;
wire local_bb4_and194_i_stall_local;
wire [31:0] local_bb4_and194_i;

assign local_bb4_and194_i_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and194_i = (rnode_180to181_bb4_add193_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and194_i_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and196_i_valid_out;
wire local_bb4_and196_i_stall_in;
wire local_bb4_and196_i_inputs_ready;
wire local_bb4_and196_i_stall_local;
wire [31:0] local_bb4_and196_i;

assign local_bb4_and196_i_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and196_i = (rnode_180to181_bb4_add193_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and196_i_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and199_i_valid_out;
wire local_bb4_and199_i_stall_in;
wire local_bb4_and199_i_inputs_ready;
wire local_bb4_and199_i_stall_local;
wire [31:0] local_bb4_and199_i;

assign local_bb4_and199_i_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and199_i = (rnode_180to181_bb4_add193_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and199_i_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and202_i_stall_local;
wire [31:0] local_bb4_and202_i;

assign local_bb4_and202_i = (rnode_180to181_bb4_add193_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_181to183_bb4__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_181to183_bb4__26_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to183_bb4__26_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to183_bb4__26_i_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_181to183_bb4__26_i_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_181to183_bb4__26_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb4__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_181to183_bb4__26_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_181to183_bb4__26_i_0_reg_183_fifo.DEPTH = 2;
defparam rnode_181to183_bb4__26_i_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_181to183_bb4__26_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to183_bb4__26_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_181to183_bb4__26_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to183_bb4__26_i_0_NO_SHIFT_REG = rnode_181to183_bb4__26_i_0_reg_183_NO_SHIFT_REG;
assign rnode_181to183_bb4__26_i_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_181to183_bb4__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i109_valid_out_2;
wire local_bb4_and17_i109_stall_in_2;
wire local_bb4_var__u31_valid_out;
wire local_bb4_var__u31_stall_in;
wire local_bb4_add192_i197_valid_out;
wire local_bb4_add192_i197_stall_in;
wire local_bb4__26_i133_valid_out;
wire local_bb4__26_i133_stall_in;
wire local_bb4__26_i133_inputs_ready;
wire local_bb4__26_i133_stall_local;
wire local_bb4__26_i133;

assign local_bb4__26_i133_inputs_ready = (rnode_180to182_bb4_shr16_i108_0_valid_out_0_NO_SHIFT_REG & rnode_180to182_bb4_cmp27_i117_0_valid_out_2_NO_SHIFT_REG & rnode_181to182_bb4_and36_lobit_i195_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_xor188_i194_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_and20_i112_0_valid_out_0_NO_SHIFT_REG & rnode_180to182_bb4_cmp27_i117_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb4_lnot33_not_i124_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb4_cmp27_i117_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_and20_i112_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_cmp37_i120_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i133 = (local_bb4_reduction_9_i132 ? rnode_181to182_bb4_cmp37_i120_0_NO_SHIFT_REG : local_bb4__24_i128);
assign local_bb4_and17_i109_valid_out_2 = 1'b1;
assign local_bb4_var__u31_valid_out = 1'b1;
assign local_bb4_add192_i197_valid_out = 1'b1;
assign local_bb4__26_i133_valid_out = 1'b1;
assign rnode_180to182_bb4_shr16_i108_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i117_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and36_lobit_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_xor188_i194_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and20_i112_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i117_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_lnot33_not_i124_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i117_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and20_i112_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_cmp37_i120_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i31_stall_local;
wire local_bb4_brmerge_not_i31;

assign local_bb4_brmerge_not_i31 = (rnode_180to182_bb4_cmp27_i24_0_NO_SHIFT_REG & rnode_181to182_bb4_lnot33_not_i30_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_2_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_cmp37_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_cmp37_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_cmp37_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_cmp37_i_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_cmp37_i_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_cmp37_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb4_cmp37_i_1_NO_SHIFT_REG),
	.data_out(rnode_182to184_bb4_cmp37_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_cmp37_i_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_cmp37_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_182to184_bb4_cmp37_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_cmp37_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_cmp37_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_cmp37_i_0_NO_SHIFT_REG = rnode_182to184_bb4_cmp37_i_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_cmp37_i_1_NO_SHIFT_REG = rnode_182to184_bb4_cmp37_i_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to184_bb4_cmp37_i_2_NO_SHIFT_REG = rnode_182to184_bb4_cmp37_i_0_reg_184_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i62_stall_local;
wire [31:0] local_bb4_add_i62;

assign local_bb4_add_i62 = ((local_bb4__27_i42 & 32'h7FFFFF8) | (rnode_181to182_bb4_and36_lobit_i_0_NO_SHIFT_REG & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_var__u29_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u29_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u29_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u29_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u29_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u29_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u29_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u29_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_var__u29_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_var__u29_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_var__u29_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_var__u29_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_var__u29_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb4_var__u29_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb4_var__u29_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_var__u29_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_var__u29_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4_var__u29_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_var__u29_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_var__u29_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_var__u29_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u29_0_NO_SHIFT_REG = rnode_182to183_bb4_var__u29_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_var__u29_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u29_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and194_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and194_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and194_i_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and194_i_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and194_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and194_i & 32'hFFFFFFF)),
	.data_out(rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and194_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and194_i_stall_in = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and194_i_0_NO_SHIFT_REG = rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and194_i_1_NO_SHIFT_REG = rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and194_i_2_NO_SHIFT_REG = rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and196_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and196_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and196_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and196_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and196_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and196_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and196_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and196_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and196_i & 32'h1F)),
	.data_out(rnode_181to182_bb4_and196_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and196_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and196_i_stall_in = 1'b0;
assign rnode_181to182_bb4_and196_i_0_NO_SHIFT_REG = rnode_181to182_bb4_and196_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and196_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and196_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and199_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and199_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and199_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and199_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and199_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and199_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and199_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and199_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and199_i & 32'h1)),
	.data_out(rnode_181to182_bb4_and199_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and199_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and199_i_stall_in = 1'b0;
assign rnode_181to182_bb4_and199_i_0_NO_SHIFT_REG = rnode_181to182_bb4_and199_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and199_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and199_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i_stall_local;
wire [31:0] local_bb4_shr_i_i;

assign local_bb4_shr_i_i = ((local_bb4_and202_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4__26_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4__26_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4__26_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4__26_i_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4__26_i_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4__26_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_181to183_bb4__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_183to184_bb4__26_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4__26_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4__26_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4__26_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4__26_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4__26_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to183_bb4__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__26_i_0_NO_SHIFT_REG = rnode_183to184_bb4__26_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__26_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__26_i_1_NO_SHIFT_REG = rnode_183to184_bb4__26_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__26_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__26_i_2_NO_SHIFT_REG = rnode_183to184_bb4__26_i_0_reg_184_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_and17_i109_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i109_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and17_i109_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i109_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and17_i109_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i109_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i109_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i109_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_and17_i109_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_and17_i109_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_and17_i109_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_and17_i109_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_and17_i109_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i109 & 32'hFF)),
	.data_out(rnode_182to184_bb4_and17_i109_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_and17_i109_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_and17_i109_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_and17_i109_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_and17_i109_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_and17_i109_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i109_stall_in_2 = 1'b0;
assign rnode_182to184_bb4_and17_i109_0_NO_SHIFT_REG = rnode_182to184_bb4_and17_i109_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_and17_i109_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and17_i109_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_var__u31_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u31_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u31_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u31_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u31_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u31_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u31_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u31_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_var__u31_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_var__u31_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_var__u31_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_var__u31_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_var__u31_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_var__u31),
	.data_out(rnode_182to183_bb4_var__u31_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_var__u31_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_var__u31_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4_var__u31_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_var__u31_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_var__u31_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u31_stall_in = 1'b0;
assign rnode_182to183_bb4_var__u31_0_NO_SHIFT_REG = rnode_182to183_bb4_var__u31_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_var__u31_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u31_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_add192_i197_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i197_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i197_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i197_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i197_3_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i197_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i197_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_add192_i197_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_add192_i197_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_add192_i197_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_add192_i197_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_add192_i197_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_add192_i197),
	.data_out(rnode_182to183_bb4_add192_i197_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_add192_i197_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_add192_i197_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_add192_i197_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_add192_i197_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_add192_i197_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add192_i197_stall_in = 1'b0;
assign rnode_182to183_bb4_add192_i197_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add192_i197_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i197_0_NO_SHIFT_REG = rnode_182to183_bb4_add192_i197_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add192_i197_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i197_1_NO_SHIFT_REG = rnode_182to183_bb4_add192_i197_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add192_i197_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i197_2_NO_SHIFT_REG = rnode_182to183_bb4_add192_i197_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add192_i197_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i197_3_NO_SHIFT_REG = rnode_182to183_bb4_add192_i197_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4__26_i133_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i133_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i133_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i133_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i133_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i133_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i133_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i133_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4__26_i133_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4__26_i133_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4__26_i133_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4__26_i133_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4__26_i133_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4__26_i133),
	.data_out(rnode_182to183_bb4__26_i133_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4__26_i133_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4__26_i133_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4__26_i133_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4__26_i133_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4__26_i133_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i133_stall_in = 1'b0;
assign rnode_182to183_bb4__26_i133_0_NO_SHIFT_REG = rnode_182to183_bb4__26_i133_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4__26_i133_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4__26_i133_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__24_i34_stall_local;
wire local_bb4__24_i34;

assign local_bb4__24_i34 = (local_bb4_or_cond_not_i33 | local_bb4_brmerge_not_i31);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i35_stall_local;
wire local_bb4_brmerge_not_not_i35;

assign local_bb4_brmerge_not_not_i35 = (local_bb4_brmerge_not_i31 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp37_i_stall_local;
wire local_bb4_not_cmp37_i;

assign local_bb4_not_cmp37_i = (rnode_182to184_bb4_cmp37_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add192_i_stall_local;
wire [31:0] local_bb4_add192_i;

assign local_bb4_add192_i = ((local_bb4_add_i62 & 32'h7FFFFF9) + rnode_181to182_bb4_xor188_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_shr217_i_stall_local;
wire [31:0] local_bb4_shr217_i;

assign local_bb4_shr217_i = ((rnode_181to182_bb4_and194_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i_stall_local;
wire [31:0] local_bb4__pre_i;

assign local_bb4__pre_i = ((rnode_181to182_bb4_and196_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i_stall_local;
wire [31:0] local_bb4_or_i_i;

assign local_bb4_or_i_i = ((local_bb4_shr_i_i & 32'h3FFFFFF) | (local_bb4_and202_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond293_i_stall_local;
wire [31:0] local_bb4_cond293_i;

assign local_bb4_cond293_i = (rnode_183to184_bb4__26_i_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u47_stall_local;
wire [31:0] local_bb4_var__u47;

assign local_bb4_var__u47[31:1] = 31'h0;
assign local_bb4_var__u47[0] = rnode_183to184_bb4__26_i_2_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_var__u31_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u31_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u31_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u31_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u31_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u31_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u31_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u31_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_var__u31_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_var__u31_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_var__u31_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_var__u31_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_var__u31_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_182to183_bb4_var__u31_0_NO_SHIFT_REG),
	.data_out(rnode_183to184_bb4_var__u31_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_var__u31_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_var__u31_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_var__u31_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_var__u31_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_var__u31_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_var__u31_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_var__u31_0_NO_SHIFT_REG = rnode_183to184_bb4_var__u31_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_var__u31_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_var__u31_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and193_i198_valid_out;
wire local_bb4_and193_i198_stall_in;
wire local_bb4_and193_i198_inputs_ready;
wire local_bb4_and193_i198_stall_local;
wire [31:0] local_bb4_and193_i198;

assign local_bb4_and193_i198_inputs_ready = rnode_182to183_bb4_add192_i197_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and193_i198 = (rnode_182to183_bb4_add192_i197_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and193_i198_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i197_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and195_i199_valid_out;
wire local_bb4_and195_i199_stall_in;
wire local_bb4_and195_i199_inputs_ready;
wire local_bb4_and195_i199_stall_local;
wire [31:0] local_bb4_and195_i199;

assign local_bb4_and195_i199_inputs_ready = rnode_182to183_bb4_add192_i197_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and195_i199 = (rnode_182to183_bb4_add192_i197_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and195_i199_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i197_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and198_i200_valid_out;
wire local_bb4_and198_i200_stall_in;
wire local_bb4_and198_i200_inputs_ready;
wire local_bb4_and198_i200_stall_local;
wire [31:0] local_bb4_and198_i200;

assign local_bb4_and198_i200_inputs_ready = rnode_182to183_bb4_add192_i197_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and198_i200 = (rnode_182to183_bb4_add192_i197_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and198_i200_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i197_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and201_i201_stall_local;
wire [31:0] local_bb4_and201_i201;

assign local_bb4_and201_i201 = (rnode_182to183_bb4_add192_i197_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_183to185_bb4__26_i133_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i133_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i133_0_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i133_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i133_0_reg_185_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i133_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i133_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i133_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_183to185_bb4__26_i133_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to185_bb4__26_i133_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to185_bb4__26_i133_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_183to185_bb4__26_i133_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_183to185_bb4__26_i133_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(rnode_182to183_bb4__26_i133_0_NO_SHIFT_REG),
	.data_out(rnode_183to185_bb4__26_i133_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_183to185_bb4__26_i133_0_reg_185_fifo.DEPTH = 2;
defparam rnode_183to185_bb4__26_i133_0_reg_185_fifo.DATA_WIDTH = 1;
defparam rnode_183to185_bb4__26_i133_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to185_bb4__26_i133_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_183to185_bb4__26_i133_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__26_i133_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to185_bb4__26_i133_0_NO_SHIFT_REG = rnode_183to185_bb4__26_i133_0_reg_185_NO_SHIFT_REG;
assign rnode_183to185_bb4__26_i133_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_183to185_bb4__26_i133_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i36_stall_local;
wire local_bb4_reduction_7_i36;

assign local_bb4_reduction_7_i36 = (local_bb4_cmp25_i23 & local_bb4_brmerge_not_not_i35);

// This section implements an unregistered operation.
// 
wire local_bb4_or220_i_stall_local;
wire [31:0] local_bb4_or220_i;

assign local_bb4_or220_i = ((local_bb4_shr217_i & 32'h7FFFFFF) | (rnode_181to182_bb4_and199_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool214_i_stall_local;
wire local_bb4_tobool214_i;

assign local_bb4_tobool214_i = ((local_bb4__pre_i & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i_stall_local;
wire [31:0] local_bb4_shr1_i_i;

assign local_bb4_shr1_i_i = ((local_bb4_or_i_i & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i_stall_local;
wire [31:0] local_bb4_lnot_ext_i;

assign local_bb4_lnot_ext_i = ((local_bb4_var__u47 & 32'h1) ^ 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_var__u31_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u31_0_stall_in_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u31_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u31_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u31_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u31_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u31_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u31_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_var__u31_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_var__u31_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_var__u31_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_var__u31_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_var__u31_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(rnode_183to184_bb4_var__u31_0_NO_SHIFT_REG),
	.data_out(rnode_184to185_bb4_var__u31_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_var__u31_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_var__u31_0_reg_185_fifo.DATA_WIDTH = 1;
defparam rnode_184to185_bb4_var__u31_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_var__u31_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_var__u31_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_var__u31_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_var__u31_0_NO_SHIFT_REG = rnode_184to185_bb4_var__u31_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_var__u31_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_var__u31_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_and193_i198_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i198_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i198_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i198_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i198_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i198_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_and193_i198_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_and193_i198_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_and193_i198_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_and193_i198_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_and193_i198_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and193_i198 & 32'hFFFFFFF)),
	.data_out(rnode_183to184_bb4_and193_i198_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_and193_i198_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_and193_i198_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_and193_i198_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_and193_i198_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_and193_i198_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and193_i198_stall_in = 1'b0;
assign rnode_183to184_bb4_and193_i198_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i198_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_and193_i198_0_NO_SHIFT_REG = rnode_183to184_bb4_and193_i198_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and193_i198_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_and193_i198_1_NO_SHIFT_REG = rnode_183to184_bb4_and193_i198_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and193_i198_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_and193_i198_2_NO_SHIFT_REG = rnode_183to184_bb4_and193_i198_0_reg_184_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_and195_i199_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i199_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and195_i199_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i199_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and195_i199_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i199_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i199_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i199_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_and195_i199_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_and195_i199_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_and195_i199_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_and195_i199_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_and195_i199_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and195_i199 & 32'h1F)),
	.data_out(rnode_183to184_bb4_and195_i199_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_and195_i199_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_and195_i199_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_and195_i199_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_and195_i199_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_and195_i199_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and195_i199_stall_in = 1'b0;
assign rnode_183to184_bb4_and195_i199_0_NO_SHIFT_REG = rnode_183to184_bb4_and195_i199_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and195_i199_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and195_i199_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_and198_i200_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i200_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and198_i200_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i200_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and198_i200_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i200_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i200_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i200_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_and198_i200_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_and198_i200_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_and198_i200_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_and198_i200_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_and198_i200_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and198_i200 & 32'h1)),
	.data_out(rnode_183to184_bb4_and198_i200_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_and198_i200_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_and198_i200_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_and198_i200_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_and198_i200_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_and198_i200_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and198_i200_stall_in = 1'b0;
assign rnode_183to184_bb4_and198_i200_0_NO_SHIFT_REG = rnode_183to184_bb4_and198_i200_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and198_i200_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and198_i200_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i202_stall_local;
wire [31:0] local_bb4_shr_i_i202;

assign local_bb4_shr_i_i202 = ((local_bb4_and201_i201 & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4__26_i133_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i133_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4__26_i133_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4__26_i133_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4__26_i133_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4__26_i133_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4__26_i133_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_183to185_bb4__26_i133_0_NO_SHIFT_REG),
	.data_out(rnode_185to186_bb4__26_i133_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4__26_i133_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4__26_i133_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4__26_i133_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4__26_i133_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4__26_i133_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_183to185_bb4__26_i133_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i133_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i133_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__26_i133_0_NO_SHIFT_REG = rnode_185to186_bb4__26_i133_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4__26_i133_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__26_i133_1_NO_SHIFT_REG = rnode_185to186_bb4__26_i133_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4__26_i133_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__26_i133_2_NO_SHIFT_REG = rnode_185to186_bb4__26_i133_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i38_stall_local;
wire local_bb4_reduction_9_i38;

assign local_bb4_reduction_9_i38 = (local_bb4_reduction_7_i36 & local_bb4_reduction_8_i37);

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i_stall_local;
wire local_bb4__40_demorgan_i;

assign local_bb4__40_demorgan_i = (rnode_180to182_bb4_cmp38_i_0_NO_SHIFT_REG | local_bb4_tobool214_i);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i_stall_local;
wire local_bb4__42_i;

assign local_bb4__42_i = (local_bb4_tobool214_i & local_bb4_not_cmp38_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i_stall_local;
wire [31:0] local_bb4_or2_i_i;

assign local_bb4_or2_i_i = ((local_bb4_shr1_i_i & 32'h1FFFFFF) | (local_bb4_or_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_shr216_i223_stall_local;
wire [31:0] local_bb4_shr216_i223;

assign local_bb4_shr216_i223 = ((rnode_183to184_bb4_and193_i198_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i221_stall_local;
wire [31:0] local_bb4__pre_i221;

assign local_bb4__pre_i221 = ((rnode_183to184_bb4_and195_i199_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i203_stall_local;
wire [31:0] local_bb4_or_i_i203;

assign local_bb4_or_i_i203 = ((local_bb4_shr_i_i202 & 32'h3FFFFFF) | (local_bb4_and201_i201 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond292_i260_stall_local;
wire [31:0] local_bb4_cond292_i260;

assign local_bb4_cond292_i260 = (rnode_185to186_bb4__26_i133_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u48_stall_local;
wire [31:0] local_bb4_var__u48;

assign local_bb4_var__u48[31:1] = 31'h0;
assign local_bb4_var__u48[0] = rnode_185to186_bb4__26_i133_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i16_valid_out_2;
wire local_bb4_and17_i16_stall_in_2;
wire local_bb4_var__u39_valid_out;
wire local_bb4_var__u39_stall_in;
wire local_bb4_add192_i_valid_out;
wire local_bb4_add192_i_stall_in;
wire local_bb4__26_i39_valid_out;
wire local_bb4__26_i39_stall_in;
wire local_bb4__26_i39_inputs_ready;
wire local_bb4__26_i39_stall_local;
wire local_bb4__26_i39;

assign local_bb4__26_i39_inputs_ready = (rnode_180to182_bb4_shr16_i15_0_valid_out_0_NO_SHIFT_REG & rnode_180to182_bb4_cmp27_i24_0_valid_out_2_NO_SHIFT_REG & rnode_181to182_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_xor188_i_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_and20_i19_0_valid_out_0_NO_SHIFT_REG & rnode_180to182_bb4_cmp27_i24_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb4_lnot33_not_i30_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb4_cmp27_i24_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_and20_i19_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i39 = (local_bb4_reduction_9_i38 ? rnode_181to182_bb4_cmp37_i_0_NO_SHIFT_REG : local_bb4__24_i34);
assign local_bb4_and17_i16_valid_out_2 = 1'b1;
assign local_bb4_var__u39_valid_out = 1'b1;
assign local_bb4_add192_i_valid_out = 1'b1;
assign local_bb4__26_i39_valid_out = 1'b1;
assign rnode_180to182_bb4_shr16_i15_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i24_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and36_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_xor188_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and20_i19_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i24_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_lnot33_not_i30_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp27_i24_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and20_i19_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__43_i_stall_local;
wire [31:0] local_bb4__43_i;

assign local_bb4__43_i = (local_bb4__42_i ? 32'h0 : (local_bb4__pre_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i_stall_local;
wire [31:0] local_bb4_shr3_i_i;

assign local_bb4_shr3_i_i = ((local_bb4_or2_i_i & 32'h7FFFFFF) >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_or219_i224_stall_local;
wire [31:0] local_bb4_or219_i224;

assign local_bb4_or219_i224 = ((local_bb4_shr216_i223 & 32'h7FFFFFF) | (rnode_183to184_bb4_and198_i200_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool213_i222_stall_local;
wire local_bb4_tobool213_i222;

assign local_bb4_tobool213_i222 = ((local_bb4__pre_i221 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i204_stall_local;
wire [31:0] local_bb4_shr1_i_i204;

assign local_bb4_shr1_i_i204 = ((local_bb4_or_i_i203 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i270_stall_local;
wire [31:0] local_bb4_lnot_ext_i270;

assign local_bb4_lnot_ext_i270 = ((local_bb4_var__u48 & 32'h1) ^ 32'h1);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_and17_i16_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i16_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and17_i16_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i16_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and17_i16_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i16_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i16_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and17_i16_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_and17_i16_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_and17_i16_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_and17_i16_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_and17_i16_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_and17_i16_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i16 & 32'hFF)),
	.data_out(rnode_182to184_bb4_and17_i16_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_and17_i16_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_and17_i16_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_and17_i16_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_and17_i16_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_and17_i16_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i16_stall_in_2 = 1'b0;
assign rnode_182to184_bb4_and17_i16_0_NO_SHIFT_REG = rnode_182to184_bb4_and17_i16_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_and17_i16_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and17_i16_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_var__u39_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u39_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u39_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u39_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u39_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u39_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u39_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u39_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_var__u39_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_var__u39_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_var__u39_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_var__u39_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_var__u39_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_var__u39),
	.data_out(rnode_182to183_bb4_var__u39_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_var__u39_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_var__u39_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4_var__u39_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_var__u39_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_var__u39_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u39_stall_in = 1'b0;
assign rnode_182to183_bb4_var__u39_0_NO_SHIFT_REG = rnode_182to183_bb4_var__u39_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_var__u39_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u39_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i_3_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add192_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add192_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_add192_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_add192_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_add192_i_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_add192_i_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_add192_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_add192_i),
	.data_out(rnode_182to183_bb4_add192_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_add192_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_add192_i_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_add192_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_add192_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_add192_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add192_i_stall_in = 1'b0;
assign rnode_182to183_bb4_add192_i_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i_0_NO_SHIFT_REG = rnode_182to183_bb4_add192_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i_1_NO_SHIFT_REG = rnode_182to183_bb4_add192_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i_2_NO_SHIFT_REG = rnode_182to183_bb4_add192_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add192_i_3_NO_SHIFT_REG = rnode_182to183_bb4_add192_i_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4__26_i39_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i39_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i39_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i39_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i39_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i39_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i39_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__26_i39_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4__26_i39_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4__26_i39_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4__26_i39_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4__26_i39_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4__26_i39_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4__26_i39),
	.data_out(rnode_182to183_bb4__26_i39_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4__26_i39_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4__26_i39_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4__26_i39_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4__26_i39_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4__26_i39_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i39_stall_in = 1'b0;
assign rnode_182to183_bb4__26_i39_0_NO_SHIFT_REG = rnode_182to183_bb4__26_i39_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4__26_i39_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4__26_i39_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i_stall_local;
wire [31:0] local_bb4_or4_i_i;

assign local_bb4_or4_i_i = ((local_bb4_shr3_i_i & 32'h7FFFFF) | (local_bb4_or2_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i225_stall_local;
wire local_bb4__40_demorgan_i225;

assign local_bb4__40_demorgan_i225 = (rnode_182to184_bb4_cmp37_i120_0_NO_SHIFT_REG | local_bb4_tobool213_i222);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i227_stall_local;
wire local_bb4__42_i227;

assign local_bb4__42_i227 = (local_bb4_tobool213_i222 & local_bb4_not_cmp37_i226);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i205_stall_local;
wire [31:0] local_bb4_or2_i_i205;

assign local_bb4_or2_i_i205 = ((local_bb4_shr1_i_i204 & 32'h1FFFFFF) | (local_bb4_or_i_i203 & 32'h7FFFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_var__u39_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u39_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u39_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u39_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u39_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u39_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u39_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_var__u39_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_var__u39_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_var__u39_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_var__u39_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_var__u39_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_var__u39_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_182to183_bb4_var__u39_0_NO_SHIFT_REG),
	.data_out(rnode_183to184_bb4_var__u39_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_var__u39_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_var__u39_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_var__u39_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_var__u39_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_var__u39_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_var__u39_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_var__u39_0_NO_SHIFT_REG = rnode_183to184_bb4_var__u39_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_var__u39_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_var__u39_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and193_i_valid_out;
wire local_bb4_and193_i_stall_in;
wire local_bb4_and193_i_inputs_ready;
wire local_bb4_and193_i_stall_local;
wire [31:0] local_bb4_and193_i;

assign local_bb4_and193_i_inputs_ready = rnode_182to183_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and193_i = (rnode_182to183_bb4_add192_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and193_i_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and195_i_valid_out;
wire local_bb4_and195_i_stall_in;
wire local_bb4_and195_i_inputs_ready;
wire local_bb4_and195_i_stall_local;
wire [31:0] local_bb4_and195_i;

assign local_bb4_and195_i_inputs_ready = rnode_182to183_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and195_i = (rnode_182to183_bb4_add192_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and195_i_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and198_i_valid_out;
wire local_bb4_and198_i_stall_in;
wire local_bb4_and198_i_inputs_ready;
wire local_bb4_and198_i_stall_local;
wire [31:0] local_bb4_and198_i;

assign local_bb4_and198_i_inputs_ready = rnode_182to183_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and198_i = (rnode_182to183_bb4_add192_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and198_i_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and201_i_stall_local;
wire [31:0] local_bb4_and201_i;

assign local_bb4_and201_i = (rnode_182to183_bb4_add192_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_183to185_bb4__26_i39_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i39_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i39_0_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i39_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i39_0_reg_185_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i39_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i39_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_183to185_bb4__26_i39_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_183to185_bb4__26_i39_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to185_bb4__26_i39_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to185_bb4__26_i39_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_183to185_bb4__26_i39_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_183to185_bb4__26_i39_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(rnode_182to183_bb4__26_i39_0_NO_SHIFT_REG),
	.data_out(rnode_183to185_bb4__26_i39_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_183to185_bb4__26_i39_0_reg_185_fifo.DEPTH = 2;
defparam rnode_183to185_bb4__26_i39_0_reg_185_fifo.DATA_WIDTH = 1;
defparam rnode_183to185_bb4__26_i39_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to185_bb4__26_i39_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_183to185_bb4__26_i39_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__26_i39_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to185_bb4__26_i39_0_NO_SHIFT_REG = rnode_183to185_bb4__26_i39_0_reg_185_NO_SHIFT_REG;
assign rnode_183to185_bb4__26_i39_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_183to185_bb4__26_i39_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i_stall_local;
wire [31:0] local_bb4_shr5_i_i;

assign local_bb4_shr5_i_i = ((local_bb4_or4_i_i & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4__43_i228_stall_local;
wire [31:0] local_bb4__43_i228;

assign local_bb4__43_i228 = (local_bb4__42_i227 ? 32'h0 : (local_bb4__pre_i221 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i206_stall_local;
wire [31:0] local_bb4_shr3_i_i206;

assign local_bb4_shr3_i_i206 = ((local_bb4_or2_i_i205 & 32'h7FFFFFF) >> 32'h4);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_var__u39_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u39_0_stall_in_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u39_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u39_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u39_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u39_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u39_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_var__u39_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_var__u39_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_var__u39_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_var__u39_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_var__u39_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_var__u39_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(rnode_183to184_bb4_var__u39_0_NO_SHIFT_REG),
	.data_out(rnode_184to185_bb4_var__u39_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_var__u39_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_var__u39_0_reg_185_fifo.DATA_WIDTH = 1;
defparam rnode_184to185_bb4_var__u39_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_var__u39_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_var__u39_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_var__u39_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_var__u39_0_NO_SHIFT_REG = rnode_184to185_bb4_var__u39_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_var__u39_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_var__u39_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and193_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and193_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_and193_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_and193_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_and193_i_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_and193_i_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_and193_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and193_i & 32'hFFFFFFF)),
	.data_out(rnode_183to184_bb4_and193_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_and193_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_and193_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_and193_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_and193_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_and193_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and193_i_stall_in = 1'b0;
assign rnode_183to184_bb4_and193_i_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_and193_i_0_NO_SHIFT_REG = rnode_183to184_bb4_and193_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_and193_i_1_NO_SHIFT_REG = rnode_183to184_bb4_and193_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_and193_i_2_NO_SHIFT_REG = rnode_183to184_bb4_and193_i_0_reg_184_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_and195_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and195_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and195_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and195_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_and195_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_and195_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_and195_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_and195_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_and195_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and195_i & 32'h1F)),
	.data_out(rnode_183to184_bb4_and195_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_and195_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_and195_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_and195_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_and195_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_and195_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and195_i_stall_in = 1'b0;
assign rnode_183to184_bb4_and195_i_0_NO_SHIFT_REG = rnode_183to184_bb4_and195_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and195_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and195_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_and198_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and198_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_and198_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_and198_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_and198_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_and198_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_and198_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_and198_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_and198_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and198_i & 32'h1)),
	.data_out(rnode_183to184_bb4_and198_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_and198_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_and198_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_and198_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_and198_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_and198_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and198_i_stall_in = 1'b0;
assign rnode_183to184_bb4_and198_i_0_NO_SHIFT_REG = rnode_183to184_bb4_and198_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_and198_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and198_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i63_stall_local;
wire [31:0] local_bb4_shr_i_i63;

assign local_bb4_shr_i_i63 = ((local_bb4_and201_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4__26_i39_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__26_i39_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4__26_i39_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4__26_i39_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4__26_i39_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4__26_i39_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4__26_i39_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_183to185_bb4__26_i39_0_NO_SHIFT_REG),
	.data_out(rnode_185to186_bb4__26_i39_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4__26_i39_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4__26_i39_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4__26_i39_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4__26_i39_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4__26_i39_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_183to185_bb4__26_i39_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i39_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i39_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__26_i39_0_NO_SHIFT_REG = rnode_185to186_bb4__26_i39_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4__26_i39_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__26_i39_1_NO_SHIFT_REG = rnode_185to186_bb4__26_i39_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4__26_i39_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__26_i39_2_NO_SHIFT_REG = rnode_185to186_bb4__26_i39_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i_stall_local;
wire [31:0] local_bb4_or6_i_i;

assign local_bb4_or6_i_i = ((local_bb4_shr5_i_i & 32'h7FFFF) | (local_bb4_or4_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i207_stall_local;
wire [31:0] local_bb4_or4_i_i207;

assign local_bb4_or4_i_i207 = ((local_bb4_shr3_i_i206 & 32'h7FFFFF) | (local_bb4_or2_i_i205 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_shr216_i_stall_local;
wire [31:0] local_bb4_shr216_i;

assign local_bb4_shr216_i = ((rnode_183to184_bb4_and193_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i77_stall_local;
wire [31:0] local_bb4__pre_i77;

assign local_bb4__pre_i77 = ((rnode_183to184_bb4_and195_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i64_stall_local;
wire [31:0] local_bb4_or_i_i64;

assign local_bb4_or_i_i64 = ((local_bb4_shr_i_i63 & 32'h3FFFFFF) | (local_bb4_and201_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond292_i_stall_local;
wire [31:0] local_bb4_cond292_i;

assign local_bb4_cond292_i = (rnode_185to186_bb4__26_i39_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u49_stall_local;
wire [31:0] local_bb4_var__u49;

assign local_bb4_var__u49[31:1] = 31'h0;
assign local_bb4_var__u49[0] = rnode_185to186_bb4__26_i39_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i_stall_local;
wire [31:0] local_bb4_shr7_i_i;

assign local_bb4_shr7_i_i = ((local_bb4_or6_i_i & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i_stall_local;
wire [31:0] local_bb4_or6_masked_i_i;

assign local_bb4_or6_masked_i_i = ((local_bb4_or6_i_i & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i208_stall_local;
wire [31:0] local_bb4_shr5_i_i208;

assign local_bb4_shr5_i_i208 = ((local_bb4_or4_i_i207 & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_or219_i_stall_local;
wire [31:0] local_bb4_or219_i;

assign local_bb4_or219_i = ((local_bb4_shr216_i & 32'h7FFFFFF) | (rnode_183to184_bb4_and198_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool213_i_stall_local;
wire local_bb4_tobool213_i;

assign local_bb4_tobool213_i = ((local_bb4__pre_i77 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i65_stall_local;
wire [31:0] local_bb4_shr1_i_i65;

assign local_bb4_shr1_i_i65 = ((local_bb4_or_i_i64 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i94_stall_local;
wire [31:0] local_bb4_lnot_ext_i94;

assign local_bb4_lnot_ext_i94 = ((local_bb4_var__u49 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i_stall_local;
wire [31:0] local_bb4_neg_i_i;

assign local_bb4_neg_i_i = ((local_bb4_or6_masked_i_i & 32'h7FFFFFF) | (local_bb4_shr7_i_i & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i209_stall_local;
wire [31:0] local_bb4_or6_i_i209;

assign local_bb4_or6_i_i209 = ((local_bb4_shr5_i_i208 & 32'h7FFFF) | (local_bb4_or4_i_i207 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i78_stall_local;
wire local_bb4__40_demorgan_i78;

assign local_bb4__40_demorgan_i78 = (rnode_182to184_bb4_cmp37_i_0_NO_SHIFT_REG | local_bb4_tobool213_i);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i79_stall_local;
wire local_bb4__42_i79;

assign local_bb4__42_i79 = (local_bb4_tobool213_i & local_bb4_not_cmp37_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i66_stall_local;
wire [31:0] local_bb4_or2_i_i66;

assign local_bb4_or2_i_i66 = ((local_bb4_shr1_i_i65 & 32'h1FFFFFF) | (local_bb4_or_i_i64 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i1_stall_local;
wire [31:0] local_bb4_and_i_i1;

assign local_bb4_and_i_i1 = ((local_bb4_neg_i_i & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i210_stall_local;
wire [31:0] local_bb4_shr7_i_i210;

assign local_bb4_shr7_i_i210 = ((local_bb4_or6_i_i209 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i211_stall_local;
wire [31:0] local_bb4_or6_masked_i_i211;

assign local_bb4_or6_masked_i_i211 = ((local_bb4_or6_i_i209 & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__43_i80_stall_local;
wire [31:0] local_bb4__43_i80;

assign local_bb4__43_i80 = (local_bb4__42_i79 ? 32'h0 : (local_bb4__pre_i77 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i67_stall_local;
wire [31:0] local_bb4_shr3_i_i67;

assign local_bb4_shr3_i_i67 = ((local_bb4_or2_i_i66 & 32'h7FFFFFF) >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i1_valid_out;
wire local_bb4__and_i_i1_stall_in;
wire local_bb4__and_i_i1_inputs_ready;
wire local_bb4__and_i_i1_stall_local;
wire [31:0] local_bb4__and_i_i1;

thirtysix_six_comp local_bb4__and_i_i1_popcnt_instance (
	.data((local_bb4_and_i_i1 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i1)
);


assign local_bb4__and_i_i1_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i1_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i212_stall_local;
wire [31:0] local_bb4_neg_i_i212;

assign local_bb4_neg_i_i212 = ((local_bb4_or6_masked_i_i211 & 32'h7FFFFFF) | (local_bb4_shr7_i_i210 & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i68_stall_local;
wire [31:0] local_bb4_or4_i_i68;

assign local_bb4_or4_i_i68 = ((local_bb4_shr3_i_i67 & 32'h7FFFFF) | (local_bb4_or2_i_i66 & 32'h7FFFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4__and_i_i1_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i1_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i1_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i1_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i1_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i1_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4__and_i_i1_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4__and_i_i1_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4__and_i_i1_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4__and_i_i1_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4__and_i_i1_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i1 & 32'h3F)),
	.data_out(rnode_181to182_bb4__and_i_i1_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4__and_i_i1_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4__and_i_i1_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4__and_i_i1_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4__and_i_i1_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4__and_i_i1_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i1_stall_in = 1'b0;
assign rnode_181to182_bb4__and_i_i1_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i1_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4__and_i_i1_0_NO_SHIFT_REG = rnode_181to182_bb4__and_i_i1_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4__and_i_i1_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4__and_i_i1_1_NO_SHIFT_REG = rnode_181to182_bb4__and_i_i1_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4__and_i_i1_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4__and_i_i1_2_NO_SHIFT_REG = rnode_181to182_bb4__and_i_i1_0_reg_182_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i213_stall_local;
wire [31:0] local_bb4_and_i_i213;

assign local_bb4_and_i_i213 = ((local_bb4_neg_i_i212 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i69_stall_local;
wire [31:0] local_bb4_shr5_i_i69;

assign local_bb4_shr5_i_i69 = ((local_bb4_or4_i_i68 & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i_stall_local;
wire [31:0] local_bb4_and9_i_i;

assign local_bb4_and9_i_i = ((rnode_181to182_bb4__and_i_i1_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and204_i_stall_local;
wire [31:0] local_bb4_and204_i;

assign local_bb4_and204_i = ((rnode_181to182_bb4__and_i_i1_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and207_i_stall_local;
wire [31:0] local_bb4_and207_i;

assign local_bb4_and207_i = ((rnode_181to182_bb4__and_i_i1_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i213_valid_out;
wire local_bb4__and_i_i213_stall_in;
wire local_bb4__and_i_i213_inputs_ready;
wire local_bb4__and_i_i213_stall_local;
wire [31:0] local_bb4__and_i_i213;

thirtysix_six_comp local_bb4__and_i_i213_popcnt_instance (
	.data((local_bb4_and_i_i213 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i213)
);


assign local_bb4__and_i_i213_inputs_ready = rnode_182to183_bb4_add192_i197_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i213_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i197_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i70_stall_local;
wire [31:0] local_bb4_or6_i_i70;

assign local_bb4_or6_i_i70 = ((local_bb4_shr5_i_i69 & 32'h7FFFF) | (local_bb4_or4_i_i68 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_sub240_i_stall_local;
wire [31:0] local_bb4_sub240_i;

assign local_bb4_sub240_i = (32'h0 - (local_bb4_and9_i_i & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl205_i_stall_local;
wire [31:0] local_bb4_shl205_i;

assign local_bb4_shl205_i = ((rnode_181to182_bb4_and194_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and204_i & 32'h18));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4__and_i_i213_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i213_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i213_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i213_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i213_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i213_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4__and_i_i213_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4__and_i_i213_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4__and_i_i213_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4__and_i_i213_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4__and_i_i213_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i213 & 32'h3F)),
	.data_out(rnode_183to184_bb4__and_i_i213_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4__and_i_i213_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4__and_i_i213_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4__and_i_i213_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4__and_i_i213_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4__and_i_i213_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i213_stall_in = 1'b0;
assign rnode_183to184_bb4__and_i_i213_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i213_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__and_i_i213_0_NO_SHIFT_REG = rnode_183to184_bb4__and_i_i213_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__and_i_i213_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__and_i_i213_1_NO_SHIFT_REG = rnode_183to184_bb4__and_i_i213_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__and_i_i213_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__and_i_i213_2_NO_SHIFT_REG = rnode_183to184_bb4__and_i_i213_0_reg_184_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i71_stall_local;
wire [31:0] local_bb4_shr7_i_i71;

assign local_bb4_shr7_i_i71 = ((local_bb4_or6_i_i70 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i72_stall_local;
wire [31:0] local_bb4_or6_masked_i_i72;

assign local_bb4_or6_masked_i_i72 = ((local_bb4_or6_i_i70 & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond245_i_stall_local;
wire [31:0] local_bb4_cond245_i;

assign local_bb4_cond245_i = (rnode_180to182_bb4_cmp38_i_2_NO_SHIFT_REG ? local_bb4_sub240_i : (local_bb4__43_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i_stall_local;
wire [31:0] local_bb4_and206_i;

assign local_bb4_and206_i = (local_bb4_shl205_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i214_stall_local;
wire [31:0] local_bb4_and9_i_i214;

assign local_bb4_and9_i_i214 = ((rnode_183to184_bb4__and_i_i213_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and203_i215_stall_local;
wire [31:0] local_bb4_and203_i215;

assign local_bb4_and203_i215 = ((rnode_183to184_bb4__and_i_i213_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i217_stall_local;
wire [31:0] local_bb4_and206_i217;

assign local_bb4_and206_i217 = ((rnode_183to184_bb4__and_i_i213_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i73_stall_local;
wire [31:0] local_bb4_neg_i_i73;

assign local_bb4_neg_i_i73 = ((local_bb4_or6_masked_i_i72 & 32'h7FFFFFF) | (local_bb4_shr7_i_i71 & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb4_add246_i_stall_local;
wire [31:0] local_bb4_add246_i;

assign local_bb4_add246_i = (local_bb4_cond245_i + (rnode_180to182_bb4_and17_i_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i_stall_local;
wire [31:0] local_bb4_fold_i;

assign local_bb4_fold_i = (local_bb4_cond245_i + (rnode_180to182_bb4_shr16_i_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl208_i_stall_local;
wire [31:0] local_bb4_shl208_i;

assign local_bb4_shl208_i = ((local_bb4_and206_i & 32'h7FFFFFF) << (local_bb4_and207_i & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb4_sub239_i236_stall_local;
wire [31:0] local_bb4_sub239_i236;

assign local_bb4_sub239_i236 = (32'h0 - (local_bb4_and9_i_i214 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl204_i216_stall_local;
wire [31:0] local_bb4_shl204_i216;

assign local_bb4_shl204_i216 = ((rnode_183to184_bb4_and193_i198_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and203_i215 & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i74_stall_local;
wire [31:0] local_bb4_and_i_i74;

assign local_bb4_and_i_i74 = ((local_bb4_neg_i_i73 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and251_i_stall_local;
wire [31:0] local_bb4_and251_i;

assign local_bb4_and251_i = (local_bb4_fold_i & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i_stall_local;
wire [31:0] local_bb4_and270_i;

assign local_bb4_and270_i = (local_bb4_fold_i << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and209_i_stall_local;
wire [31:0] local_bb4_and209_i;

assign local_bb4_and209_i = (local_bb4_shl208_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond244_i237_stall_local;
wire [31:0] local_bb4_cond244_i237;

assign local_bb4_cond244_i237 = (rnode_182to184_bb4_cmp37_i120_2_NO_SHIFT_REG ? local_bb4_sub239_i236 : (local_bb4__43_i228 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and205_i218_stall_local;
wire [31:0] local_bb4_and205_i218;

assign local_bb4_and205_i218 = (local_bb4_shl204_i216 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i74_valid_out;
wire local_bb4__and_i_i74_stall_in;
wire local_bb4__and_i_i74_inputs_ready;
wire local_bb4__and_i_i74_stall_local;
wire [31:0] local_bb4__and_i_i74;

thirtysix_six_comp local_bb4__and_i_i74_popcnt_instance (
	.data((local_bb4_and_i_i74 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i74)
);


assign local_bb4__and_i_i74_inputs_ready = rnode_182to183_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i74_valid_out = 1'b1;
assign rnode_182to183_bb4_add192_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__44_i_stall_local;
wire [31:0] local_bb4__44_i;

assign local_bb4__44_i = (local_bb4__40_demorgan_i ? (local_bb4_and209_i & 32'h7FFFFFF) : (local_bb4_or220_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add245_i238_stall_local;
wire [31:0] local_bb4_add245_i238;

assign local_bb4_add245_i238 = (local_bb4_cond244_i237 + (rnode_182to184_bb4_and17_i109_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i240_stall_local;
wire [31:0] local_bb4_fold_i240;

assign local_bb4_fold_i240 = (local_bb4_cond244_i237 + (rnode_182to184_bb4_shr16_i108_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl207_i219_stall_local;
wire [31:0] local_bb4_shl207_i219;

assign local_bb4_shl207_i219 = ((local_bb4_and205_i218 & 32'h7FFFFFF) << (local_bb4_and206_i217 & 32'h7));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4__and_i_i74_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i74_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i74_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i74_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4__and_i_i74_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__and_i_i74_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4__and_i_i74_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4__and_i_i74_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4__and_i_i74_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4__and_i_i74_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4__and_i_i74_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i74 & 32'h3F)),
	.data_out(rnode_183to184_bb4__and_i_i74_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4__and_i_i74_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4__and_i_i74_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4__and_i_i74_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4__and_i_i74_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4__and_i_i74_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i74_stall_in = 1'b0;
assign rnode_183to184_bb4__and_i_i74_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i74_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__and_i_i74_0_NO_SHIFT_REG = rnode_183to184_bb4__and_i_i74_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__and_i_i74_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__and_i_i74_1_NO_SHIFT_REG = rnode_183to184_bb4__and_i_i74_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__and_i_i74_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__and_i_i74_2_NO_SHIFT_REG = rnode_183to184_bb4__and_i_i74_0_reg_184_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and251_i_valid_out;
wire local_bb4_and251_i_stall_in;
wire local_bb4_and270_i_valid_out;
wire local_bb4_and270_i_stall_in;
wire local_bb4_add246_i_valid_out;
wire local_bb4_add246_i_stall_in;
wire local_bb4__45_i_valid_out;
wire local_bb4__45_i_stall_in;
wire local_bb4_not_cmp38_i_valid_out_1;
wire local_bb4_not_cmp38_i_stall_in_1;
wire local_bb4__45_i_inputs_ready;
wire local_bb4__45_i_stall_local;
wire [31:0] local_bb4__45_i;

assign local_bb4__45_i_inputs_ready = (rnode_180to182_bb4_shr16_i_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb4_and17_i_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_and196_i_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_and199_i_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb4__and_i_i1_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4__and_i_i1_0_valid_out_2_NO_SHIFT_REG & rnode_181to182_bb4__and_i_i1_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i = (local_bb4__42_i ? (rnode_181to182_bb4_and194_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i & 32'h7FFFFFF));
assign local_bb4_and251_i_valid_out = 1'b1;
assign local_bb4_and270_i_valid_out = 1'b1;
assign local_bb4_add246_i_valid_out = 1'b1;
assign local_bb4__45_i_valid_out = 1'b1;
assign local_bb4_not_cmp38_i_valid_out_1 = 1'b1;
assign rnode_180to182_bb4_shr16_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and17_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and196_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and199_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i1_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i1_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i1_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i241_stall_local;
wire [31:0] local_bb4_and250_i241;

assign local_bb4_and250_i241 = (local_bb4_fold_i240 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and269_i252_stall_local;
wire [31:0] local_bb4_and269_i252;

assign local_bb4_and269_i252 = (local_bb4_fold_i240 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and208_i220_stall_local;
wire [31:0] local_bb4_and208_i220;

assign local_bb4_and208_i220 = (local_bb4_shl207_i219 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i75_stall_local;
wire [31:0] local_bb4_and9_i_i75;

assign local_bb4_and9_i_i75 = ((rnode_183to184_bb4__and_i_i74_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and203_i_stall_local;
wire [31:0] local_bb4_and203_i;

assign local_bb4_and203_i = ((rnode_183to184_bb4__and_i_i74_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i76_stall_local;
wire [31:0] local_bb4_and206_i76;

assign local_bb4_and206_i76 = ((rnode_183to184_bb4__and_i_i74_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_and251_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and251_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and251_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_and251_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_and251_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_and251_i_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_and251_i_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_and251_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in((local_bb4_and251_i & 32'hFF)),
	.data_out(rnode_182to183_bb4_and251_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_and251_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and251_i_stall_in = 1'b0;
assign rnode_182to183_bb4_and251_i_0_NO_SHIFT_REG = rnode_182to183_bb4_and251_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_and251_i_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and251_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_and270_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and270_i_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and270_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_and270_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_and270_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_and270_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_and270_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_and270_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and270_i & 32'hFF800000)),
	.data_out(rnode_182to184_bb4_and270_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_and270_i_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_and270_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_and270_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_and270_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_and270_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and270_i_stall_in = 1'b0;
assign rnode_182to184_bb4_and270_i_0_NO_SHIFT_REG = rnode_182to184_bb4_and270_i_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_and270_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and270_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add246_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add246_i_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_add246_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_add246_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_add246_i_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_add246_i_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_add246_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_add246_i),
	.data_out(rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_add246_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add246_i_stall_in = 1'b0;
assign rnode_182to183_bb4_add246_i_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add246_i_0_NO_SHIFT_REG = rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add246_i_1_NO_SHIFT_REG = rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4__45_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4__45_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4__45_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4__45_i_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4__45_i_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4__45_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in((local_bb4__45_i & 32'hFFFFFFF)),
	.data_out(rnode_182to183_bb4__45_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4__45_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4__45_i_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4__45_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4__45_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4__45_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i_stall_in = 1'b0;
assign rnode_182to183_bb4__45_i_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4__45_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__45_i_0_NO_SHIFT_REG = rnode_182to183_bb4__45_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4__45_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__45_i_1_NO_SHIFT_REG = rnode_182to183_bb4__45_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4__45_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__45_i_2_NO_SHIFT_REG = rnode_182to183_bb4__45_i_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_not_cmp38_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_not_cmp38_i_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_not_cmp38_i_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_not_cmp38_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp38_i),
	.data_out(rnode_182to183_bb4_not_cmp38_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_not_cmp38_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp38_i_stall_in_1 = 1'b0;
assign rnode_182to183_bb4_not_cmp38_i_0_NO_SHIFT_REG = rnode_182to183_bb4_not_cmp38_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_not_cmp38_i_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__44_i229_stall_local;
wire [31:0] local_bb4__44_i229;

assign local_bb4__44_i229 = (local_bb4__40_demorgan_i225 ? (local_bb4_and208_i220 & 32'h7FFFFFF) : (local_bb4_or219_i224 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_sub239_i_stall_local;
wire [31:0] local_bb4_sub239_i;

assign local_bb4_sub239_i = (32'h0 - (local_bb4_and9_i_i75 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl204_i_stall_local;
wire [31:0] local_bb4_shl204_i;

assign local_bb4_shl204_i = ((rnode_183to184_bb4_and193_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and203_i & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i_stall_local;
wire local_bb4_notrhs_i;

assign local_bb4_notrhs_i = ((rnode_182to183_bb4_and251_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl274_i_stall_local;
wire [31:0] local_bb4_shl274_i;

assign local_bb4_shl274_i = ((rnode_182to184_bb4_and270_i_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and248_i_stall_local;
wire [31:0] local_bb4_and248_i;

assign local_bb4_and248_i = (rnode_182to183_bb4_add246_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp259_i_stall_local;
wire local_bb4_cmp259_i;

assign local_bb4_cmp259_i = ($signed(rnode_182to183_bb4_add246_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and226_i_stall_local;
wire [31:0] local_bb4_and226_i;

assign local_bb4_and226_i = ((rnode_182to183_bb4__45_i_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and271_i_stall_local;
wire [31:0] local_bb4_and271_i;

assign local_bb4_and271_i = ((rnode_182to183_bb4__45_i_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr272_i_valid_out;
wire local_bb4_shr272_i_stall_in;
wire local_bb4_shr272_i_inputs_ready;
wire local_bb4_shr272_i_stall_local;
wire [31:0] local_bb4_shr272_i;

assign local_bb4_shr272_i_inputs_ready = rnode_182to183_bb4__45_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr272_i = ((rnode_182to183_bb4__45_i_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr272_i_valid_out = 1'b1;
assign rnode_182to183_bb4__45_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i241_valid_out;
wire local_bb4_and250_i241_stall_in;
wire local_bb4_and269_i252_valid_out;
wire local_bb4_and269_i252_stall_in;
wire local_bb4_add245_i238_valid_out;
wire local_bb4_add245_i238_stall_in;
wire local_bb4__45_i230_valid_out;
wire local_bb4__45_i230_stall_in;
wire local_bb4_not_cmp37_i226_valid_out_1;
wire local_bb4_not_cmp37_i226_stall_in_1;
wire local_bb4__45_i230_inputs_ready;
wire local_bb4__45_i230_stall_local;
wire [31:0] local_bb4__45_i230;

assign local_bb4__45_i230_inputs_ready = (rnode_182to184_bb4_shr16_i108_0_valid_out_NO_SHIFT_REG & rnode_182to184_bb4_and17_i109_0_valid_out_NO_SHIFT_REG & rnode_182to184_bb4_cmp37_i120_0_valid_out_2_NO_SHIFT_REG & rnode_182to184_bb4_cmp37_i120_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4_and193_i198_0_valid_out_2_NO_SHIFT_REG & rnode_182to184_bb4_cmp37_i120_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4_and195_i199_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_and193_i198_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4_and198_i200_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_and193_i198_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4__and_i_i213_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4__and_i_i213_0_valid_out_2_NO_SHIFT_REG & rnode_183to184_bb4__and_i_i213_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i230 = (local_bb4__42_i227 ? (rnode_183to184_bb4_and193_i198_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i229 & 32'h7FFFFFF));
assign local_bb4_and250_i241_valid_out = 1'b1;
assign local_bb4_and269_i252_valid_out = 1'b1;
assign local_bb4_add245_i238_valid_out = 1'b1;
assign local_bb4__45_i230_valid_out = 1'b1;
assign local_bb4_not_cmp37_i226_valid_out_1 = 1'b1;
assign rnode_182to184_bb4_shr16_i108_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and17_i109_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i120_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i120_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i198_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i120_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and195_i199_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i198_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and198_i200_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i198_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i213_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i213_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i213_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cond244_i_stall_local;
wire [31:0] local_bb4_cond244_i;

assign local_bb4_cond244_i = (rnode_182to184_bb4_cmp37_i_2_NO_SHIFT_REG ? local_bb4_sub239_i : (local_bb4__43_i80 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and205_i_stall_local;
wire [31:0] local_bb4_and205_i;

assign local_bb4_and205_i = (local_bb4_shl204_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i_stall_local;
wire local_bb4_notlhs_i;

assign local_bb4_notlhs_i = ((local_bb4_and248_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp227_i_stall_local;
wire local_bb4_cmp227_i;

assign local_bb4_cmp227_i = ((local_bb4_and226_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp297_i_stall_local;
wire local_bb4_cmp297_i;

assign local_bb4_cmp297_i = ((local_bb4_and271_i & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp297_i_valid_out;
wire local_bb4_cmp297_i_stall_in;
wire local_bb4_cmp300_i_valid_out;
wire local_bb4_cmp300_i_stall_in;
wire local_bb4_cmp300_i_inputs_ready;
wire local_bb4_cmp300_i_stall_local;
wire local_bb4_cmp300_i;

assign local_bb4_cmp300_i_inputs_ready = rnode_182to183_bb4__45_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp300_i = ((local_bb4_and271_i & 32'h7) == 32'h4);
assign local_bb4_cmp297_i_valid_out = 1'b1;
assign local_bb4_cmp300_i_valid_out = 1'b1;
assign rnode_182to183_bb4__45_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_shr272_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_shr272_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_shr272_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_shr272_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_shr272_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_shr272_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_shr272_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_shr272_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_shr272_i & 32'h1FFFFFF)),
	.data_out(rnode_183to184_bb4_shr272_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_shr272_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr272_i_stall_in = 1'b0;
assign rnode_183to184_bb4_shr272_i_0_NO_SHIFT_REG = rnode_183to184_bb4_shr272_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_shr272_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_shr272_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_and250_i241_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i241_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and250_i241_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i241_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and250_i241_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i241_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i241_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i241_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_and250_i241_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_and250_i241_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_and250_i241_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_and250_i241_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_and250_i241_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in((local_bb4_and250_i241 & 32'hFF)),
	.data_out(rnode_184to185_bb4_and250_i241_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_and250_i241_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_and250_i241_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4_and250_i241_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_and250_i241_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_and250_i241_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and250_i241_stall_in = 1'b0;
assign rnode_184to185_bb4_and250_i241_0_NO_SHIFT_REG = rnode_184to185_bb4_and250_i241_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_and250_i241_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and250_i241_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_184to186_bb4_and269_i252_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i252_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_184to186_bb4_and269_i252_0_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i252_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to186_bb4_and269_i252_0_reg_186_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i252_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i252_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i252_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_184to186_bb4_and269_i252_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to186_bb4_and269_i252_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to186_bb4_and269_i252_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_184to186_bb4_and269_i252_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_184to186_bb4_and269_i252_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in((local_bb4_and269_i252 & 32'hFF800000)),
	.data_out(rnode_184to186_bb4_and269_i252_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_184to186_bb4_and269_i252_0_reg_186_fifo.DEPTH = 2;
defparam rnode_184to186_bb4_and269_i252_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_184to186_bb4_and269_i252_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to186_bb4_and269_i252_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_184to186_bb4_and269_i252_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and269_i252_stall_in = 1'b0;
assign rnode_184to186_bb4_and269_i252_0_NO_SHIFT_REG = rnode_184to186_bb4_and269_i252_0_reg_186_NO_SHIFT_REG;
assign rnode_184to186_bb4_and269_i252_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_184to186_bb4_and269_i252_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_add245_i238_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i238_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_add245_i238_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i238_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i238_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_add245_i238_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i238_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_add245_i238_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i238_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i238_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i238_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_add245_i238_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_add245_i238_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_add245_i238_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_add245_i238_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_add245_i238_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(local_bb4_add245_i238),
	.data_out(rnode_184to185_bb4_add245_i238_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_add245_i238_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_add245_i238_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4_add245_i238_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_add245_i238_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_add245_i238_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add245_i238_stall_in = 1'b0;
assign rnode_184to185_bb4_add245_i238_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_add245_i238_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4_add245_i238_0_NO_SHIFT_REG = rnode_184to185_bb4_add245_i238_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_add245_i238_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4_add245_i238_1_NO_SHIFT_REG = rnode_184to185_bb4_add245_i238_0_reg_185_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4__45_i230_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i230_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i230_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i230_2_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i230_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i230_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4__45_i230_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4__45_i230_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4__45_i230_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4__45_i230_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4__45_i230_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in((local_bb4__45_i230 & 32'hFFFFFFF)),
	.data_out(rnode_184to185_bb4__45_i230_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4__45_i230_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4__45_i230_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4__45_i230_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4__45_i230_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4__45_i230_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i230_stall_in = 1'b0;
assign rnode_184to185_bb4__45_i230_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4__45_i230_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4__45_i230_0_NO_SHIFT_REG = rnode_184to185_bb4__45_i230_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4__45_i230_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4__45_i230_1_NO_SHIFT_REG = rnode_184to185_bb4__45_i230_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4__45_i230_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4__45_i230_2_NO_SHIFT_REG = rnode_184to185_bb4__45_i230_0_reg_185_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_not_cmp37_i226_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i226_0_stall_in_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i226_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i226_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i226_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i226_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i226_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i226_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_not_cmp37_i226_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_not_cmp37_i226_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_not_cmp37_i226_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_not_cmp37_i226_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_not_cmp37_i226_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp37_i226),
	.data_out(rnode_184to185_bb4_not_cmp37_i226_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_not_cmp37_i226_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_not_cmp37_i226_0_reg_185_fifo.DATA_WIDTH = 1;
defparam rnode_184to185_bb4_not_cmp37_i226_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_not_cmp37_i226_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_not_cmp37_i226_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp37_i226_stall_in_1 = 1'b0;
assign rnode_184to185_bb4_not_cmp37_i226_0_NO_SHIFT_REG = rnode_184to185_bb4_not_cmp37_i226_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_not_cmp37_i226_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_not_cmp37_i226_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_add245_i_stall_local;
wire [31:0] local_bb4_add245_i;

assign local_bb4_add245_i = (local_bb4_cond244_i + (rnode_182to184_bb4_and17_i16_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i85_stall_local;
wire [31:0] local_bb4_fold_i85;

assign local_bb4_fold_i85 = (local_bb4_cond244_i + (rnode_182to184_bb4_shr16_i15_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl207_i_stall_local;
wire [31:0] local_bb4_shl207_i;

assign local_bb4_shl207_i = ((local_bb4_and205_i & 32'h7FFFFFF) << (local_bb4_and206_i76 & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i_stall_local;
wire local_bb4_not__46_i;

assign local_bb4_not__46_i = (local_bb4_notrhs_i | local_bb4_notlhs_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp227_not_i_stall_local;
wire local_bb4_cmp227_not_i;

assign local_bb4_cmp227_not_i = (local_bb4_cmp227_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_cmp297_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_cmp297_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_cmp297_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_cmp297_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_cmp297_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4_cmp297_i),
	.data_out(rnode_183to184_bb4_cmp297_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_cmp297_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp297_i_stall_in = 1'b0;
assign rnode_183to184_bb4_cmp297_i_0_NO_SHIFT_REG = rnode_183to184_bb4_cmp297_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_cmp297_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_cmp300_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_cmp300_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_cmp300_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_cmp300_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_cmp300_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4_cmp300_i),
	.data_out(rnode_183to184_bb4_cmp300_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_cmp300_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp300_i_stall_in = 1'b0;
assign rnode_183to184_bb4_cmp300_i_0_NO_SHIFT_REG = rnode_183to184_bb4_cmp300_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_cmp300_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and273_i_stall_local;
wire [31:0] local_bb4_and273_i;

assign local_bb4_and273_i = ((rnode_183to184_bb4_shr272_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i243_stall_local;
wire local_bb4_notrhs_i243;

assign local_bb4_notrhs_i243 = ((rnode_184to185_bb4_and250_i241_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl273_i253_stall_local;
wire [31:0] local_bb4_shl273_i253;

assign local_bb4_shl273_i253 = ((rnode_184to186_bb4_and269_i252_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and247_i239_stall_local;
wire [31:0] local_bb4_and247_i239;

assign local_bb4_and247_i239 = (rnode_184to185_bb4_add245_i238_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp258_i246_stall_local;
wire local_bb4_cmp258_i246;

assign local_bb4_cmp258_i246 = ($signed(rnode_184to185_bb4_add245_i238_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and225_i231_stall_local;
wire [31:0] local_bb4_and225_i231;

assign local_bb4_and225_i231 = ((rnode_184to185_bb4__45_i230_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i249_stall_local;
wire [31:0] local_bb4_and270_i249;

assign local_bb4_and270_i249 = ((rnode_184to185_bb4__45_i230_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr271_i250_valid_out;
wire local_bb4_shr271_i250_stall_in;
wire local_bb4_shr271_i250_inputs_ready;
wire local_bb4_shr271_i250_stall_local;
wire [31:0] local_bb4_shr271_i250;

assign local_bb4_shr271_i250_inputs_ready = rnode_184to185_bb4__45_i230_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr271_i250 = ((rnode_184to185_bb4__45_i230_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr271_i250_valid_out = 1'b1;
assign rnode_184to185_bb4__45_i230_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i_stall_local;
wire [31:0] local_bb4_and250_i;

assign local_bb4_and250_i = (local_bb4_fold_i85 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and269_i_stall_local;
wire [31:0] local_bb4_and269_i;

assign local_bb4_and269_i = (local_bb4_fold_i85 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and208_i_stall_local;
wire [31:0] local_bb4_and208_i;

assign local_bb4_and208_i = (local_bb4_shl207_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__47_i_stall_local;
wire local_bb4__47_i;

assign local_bb4__47_i = (local_bb4_cmp227_i | local_bb4_not__46_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i_stall_local;
wire local_bb4_brmerge12_i;

assign local_bb4_brmerge12_i = (local_bb4_cmp227_not_i | rnode_182to183_bb4_not_cmp38_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot263__i_stall_local;
wire local_bb4_lnot263__i;

assign local_bb4_lnot263__i = (local_bb4_cmp259_i & local_bb4_cmp227_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29749_i_stall_local;
wire [31:0] local_bb4_cmp29749_i;

assign local_bb4_cmp29749_i[31:1] = 31'h0;
assign local_bb4_cmp29749_i[0] = rnode_183to184_bb4_cmp297_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv301_i_stall_local;
wire [31:0] local_bb4_conv301_i;

assign local_bb4_conv301_i[31:1] = 31'h0;
assign local_bb4_conv301_i[0] = rnode_183to184_bb4_cmp300_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i_stall_local;
wire [31:0] local_bb4_or275_i;

assign local_bb4_or275_i = ((local_bb4_and273_i & 32'h7FFFFF) | (local_bb4_shl274_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i242_stall_local;
wire local_bb4_notlhs_i242;

assign local_bb4_notlhs_i242 = ((local_bb4_and247_i239 & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_i232_stall_local;
wire local_bb4_cmp226_i232;

assign local_bb4_cmp226_i232 = ((local_bb4_and225_i231 & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i264_stall_local;
wire local_bb4_cmp296_i264;

assign local_bb4_cmp296_i264 = ((local_bb4_and270_i249 & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i264_valid_out;
wire local_bb4_cmp296_i264_stall_in;
wire local_bb4_cmp299_i265_valid_out;
wire local_bb4_cmp299_i265_stall_in;
wire local_bb4_cmp299_i265_inputs_ready;
wire local_bb4_cmp299_i265_stall_local;
wire local_bb4_cmp299_i265;

assign local_bb4_cmp299_i265_inputs_ready = rnode_184to185_bb4__45_i230_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp299_i265 = ((local_bb4_and270_i249 & 32'h7) == 32'h4);
assign local_bb4_cmp296_i264_valid_out = 1'b1;
assign local_bb4_cmp299_i265_valid_out = 1'b1;
assign rnode_184to185_bb4__45_i230_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_shr271_i250_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i250_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_shr271_i250_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i250_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_shr271_i250_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i250_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i250_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i250_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_shr271_i250_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_shr271_i250_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_shr271_i250_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_shr271_i250_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_shr271_i250_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in((local_bb4_shr271_i250 & 32'h1FFFFFF)),
	.data_out(rnode_185to186_bb4_shr271_i250_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_shr271_i250_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_shr271_i250_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb4_shr271_i250_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_shr271_i250_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_shr271_i250_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr271_i250_stall_in = 1'b0;
assign rnode_185to186_bb4_shr271_i250_0_NO_SHIFT_REG = rnode_185to186_bb4_shr271_i250_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_shr271_i250_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_shr271_i250_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__44_i81_stall_local;
wire [31:0] local_bb4__44_i81;

assign local_bb4__44_i81 = (local_bb4__40_demorgan_i78 ? (local_bb4_and208_i & 32'h7FFFFFF) : (local_bb4_or219_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i_stall_local;
wire [31:0] local_bb4_resultSign_0_i;

assign local_bb4_resultSign_0_i = (local_bb4_brmerge12_i ? (rnode_182to183_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i_valid_out;
wire local_bb4_resultSign_0_i_stall_in;
wire local_bb4__47_i_valid_out;
wire local_bb4__47_i_stall_in;
wire local_bb4_or2672_i_valid_out;
wire local_bb4_or2672_i_stall_in;
wire local_bb4_or2672_i_inputs_ready;
wire local_bb4_or2672_i_stall_local;
wire local_bb4_or2672_i;

assign local_bb4_or2672_i_inputs_ready = (rnode_182to183_bb4_and35_i_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb4_and251_i_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb4__45_i_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG & rnode_182to183_bb4_var__u29_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2672_i = (rnode_182to183_bb4_var__u29_0_NO_SHIFT_REG | local_bb4_lnot263__i);
assign local_bb4_resultSign_0_i_valid_out = 1'b1;
assign local_bb4__47_i_valid_out = 1'b1;
assign local_bb4_or2672_i_valid_out = 1'b1;
assign rnode_182to183_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_not_cmp38_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add246_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and251_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4__45_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add246_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u29_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i244_stall_local;
wire local_bb4_not__46_i244;

assign local_bb4_not__46_i244 = (local_bb4_notrhs_i243 | local_bb4_notlhs_i242);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_not_i233_stall_local;
wire local_bb4_cmp226_not_i233;

assign local_bb4_cmp226_not_i233 = (local_bb4_cmp226_i232 ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_cmp296_i264_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i264_0_stall_in_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i264_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i264_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i264_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i264_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i264_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i264_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_cmp296_i264_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_cmp296_i264_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_cmp296_i264_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_cmp296_i264_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_cmp296_i264_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4_cmp296_i264),
	.data_out(rnode_185to186_bb4_cmp296_i264_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_cmp296_i264_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_cmp296_i264_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4_cmp296_i264_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_cmp296_i264_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_cmp296_i264_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp296_i264_stall_in = 1'b0;
assign rnode_185to186_bb4_cmp296_i264_0_NO_SHIFT_REG = rnode_185to186_bb4_cmp296_i264_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_cmp296_i264_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp296_i264_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_cmp299_i265_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i265_0_stall_in_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i265_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i265_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i265_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i265_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i265_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i265_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_cmp299_i265_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_cmp299_i265_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_cmp299_i265_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_cmp299_i265_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_cmp299_i265_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4_cmp299_i265),
	.data_out(rnode_185to186_bb4_cmp299_i265_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_cmp299_i265_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_cmp299_i265_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4_cmp299_i265_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_cmp299_i265_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_cmp299_i265_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp299_i265_stall_in = 1'b0;
assign rnode_185to186_bb4_cmp299_i265_0_NO_SHIFT_REG = rnode_185to186_bb4_cmp299_i265_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_cmp299_i265_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp299_i265_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and272_i251_stall_local;
wire [31:0] local_bb4_and272_i251;

assign local_bb4_and272_i251 = ((rnode_185to186_bb4_shr271_i250_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i_valid_out;
wire local_bb4_and250_i_stall_in;
wire local_bb4_and269_i_valid_out;
wire local_bb4_and269_i_stall_in;
wire local_bb4_add245_i_valid_out;
wire local_bb4_add245_i_stall_in;
wire local_bb4__45_i82_valid_out;
wire local_bb4__45_i82_stall_in;
wire local_bb4_not_cmp37_i_valid_out_1;
wire local_bb4_not_cmp37_i_stall_in_1;
wire local_bb4__45_i82_inputs_ready;
wire local_bb4__45_i82_stall_local;
wire [31:0] local_bb4__45_i82;

assign local_bb4__45_i82_inputs_ready = (rnode_182to184_bb4_shr16_i15_0_valid_out_NO_SHIFT_REG & rnode_182to184_bb4_and17_i16_0_valid_out_NO_SHIFT_REG & rnode_182to184_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG & rnode_182to184_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG & rnode_182to184_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4_and195_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4_and198_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4__and_i_i74_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4__and_i_i74_0_valid_out_2_NO_SHIFT_REG & rnode_183to184_bb4__and_i_i74_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i82 = (local_bb4__42_i79 ? (rnode_183to184_bb4_and193_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i81 & 32'h7FFFFFF));
assign local_bb4_and250_i_valid_out = 1'b1;
assign local_bb4_and269_i_valid_out = 1'b1;
assign local_bb4_add245_i_valid_out = 1'b1;
assign local_bb4__45_i82_valid_out = 1'b1;
assign local_bb4_not_cmp37_i_valid_out_1 = 1'b1;
assign rnode_182to184_bb4_shr16_i15_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and17_i16_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and195_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and198_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_and193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i74_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i74_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__and_i_i74_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_resultSign_0_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_resultSign_0_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_resultSign_0_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_resultSign_0_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_resultSign_0_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_resultSign_0_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_resultSign_0_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i & 32'h80000000)),
	.data_out(rnode_183to184_bb4_resultSign_0_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_resultSign_0_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_resultSign_0_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_resultSign_0_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_resultSign_0_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_resultSign_0_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i_stall_in = 1'b0;
assign rnode_183to184_bb4_resultSign_0_i_0_NO_SHIFT_REG = rnode_183to184_bb4_resultSign_0_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_resultSign_0_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4__47_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4__47_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4__47_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4__47_i_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4__47_i_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4__47_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4__47_i),
	.data_out(rnode_183to184_bb4__47_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4__47_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4__47_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4__47_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4__47_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4__47_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i_stall_in = 1'b0;
assign rnode_183to184_bb4__47_i_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__47_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__47_i_0_NO_SHIFT_REG = rnode_183to184_bb4__47_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__47_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__47_i_1_NO_SHIFT_REG = rnode_183to184_bb4__47_i_0_reg_184_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_or2672_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_or2672_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_or2672_i_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_or2672_i_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_or2672_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4_or2672_i),
	.data_out(rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_or2672_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2672_i_stall_in = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_or2672_i_0_NO_SHIFT_REG = rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_or2672_i_1_NO_SHIFT_REG = rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_or2672_i_2_NO_SHIFT_REG = rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__47_i245_stall_local;
wire local_bb4__47_i245;

assign local_bb4__47_i245 = (local_bb4_cmp226_i232 | local_bb4_not__46_i244);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i234_stall_local;
wire local_bb4_brmerge12_i234;

assign local_bb4_brmerge12_i234 = (local_bb4_cmp226_not_i233 | rnode_184to185_bb4_not_cmp37_i226_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot262__i247_stall_local;
wire local_bb4_lnot262__i247;

assign local_bb4_lnot262__i247 = (local_bb4_cmp258_i246 & local_bb4_cmp226_not_i233);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29649_i268_stall_local;
wire [31:0] local_bb4_cmp29649_i268;

assign local_bb4_cmp29649_i268[31:1] = 31'h0;
assign local_bb4_cmp29649_i268[0] = rnode_185to186_bb4_cmp296_i264_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv300_i266_stall_local;
wire [31:0] local_bb4_conv300_i266;

assign local_bb4_conv300_i266[31:1] = 31'h0;
assign local_bb4_conv300_i266[0] = rnode_185to186_bb4_cmp299_i265_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or274_i254_stall_local;
wire [31:0] local_bb4_or274_i254;

assign local_bb4_or274_i254 = ((local_bb4_and272_i251 & 32'h7FFFFF) | (local_bb4_shl273_i253 & 32'h7F800000));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_and250_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and250_i_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_and250_i_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_and250_i_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_and250_i_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_and250_i_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_and250_i_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_and250_i_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_and250_i_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in((local_bb4_and250_i & 32'hFF)),
	.data_out(rnode_184to185_bb4_and250_i_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_and250_i_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_and250_i_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4_and250_i_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_and250_i_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_and250_i_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and250_i_stall_in = 1'b0;
assign rnode_184to185_bb4_and250_i_0_NO_SHIFT_REG = rnode_184to185_bb4_and250_i_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_and250_i_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and250_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_184to186_bb4_and269_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_184to186_bb4_and269_i_0_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to186_bb4_and269_i_0_reg_186_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_184to186_bb4_and269_i_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_184to186_bb4_and269_i_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to186_bb4_and269_i_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to186_bb4_and269_i_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_184to186_bb4_and269_i_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_184to186_bb4_and269_i_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in((local_bb4_and269_i & 32'hFF800000)),
	.data_out(rnode_184to186_bb4_and269_i_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_184to186_bb4_and269_i_0_reg_186_fifo.DEPTH = 2;
defparam rnode_184to186_bb4_and269_i_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_184to186_bb4_and269_i_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to186_bb4_and269_i_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_184to186_bb4_and269_i_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and269_i_stall_in = 1'b0;
assign rnode_184to186_bb4_and269_i_0_NO_SHIFT_REG = rnode_184to186_bb4_and269_i_0_reg_186_NO_SHIFT_REG;
assign rnode_184to186_bb4_and269_i_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_184to186_bb4_and269_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_add245_i_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_add245_i_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4_add245_i_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_add245_i_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_add245_i_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_add245_i_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_add245_i_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_add245_i_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_add245_i_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(local_bb4_add245_i),
	.data_out(rnode_184to185_bb4_add245_i_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_add245_i_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_add245_i_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4_add245_i_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_add245_i_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_add245_i_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add245_i_stall_in = 1'b0;
assign rnode_184to185_bb4_add245_i_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4_add245_i_0_NO_SHIFT_REG = rnode_184to185_bb4_add245_i_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4_add245_i_1_NO_SHIFT_REG = rnode_184to185_bb4_add245_i_0_reg_185_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4__45_i82_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i82_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i82_1_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i82_2_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb4__45_i82_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4__45_i82_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4__45_i82_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4__45_i82_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4__45_i82_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4__45_i82_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4__45_i82_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in((local_bb4__45_i82 & 32'hFFFFFFF)),
	.data_out(rnode_184to185_bb4__45_i82_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4__45_i82_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4__45_i82_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb4__45_i82_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4__45_i82_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4__45_i82_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i82_stall_in = 1'b0;
assign rnode_184to185_bb4__45_i82_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4__45_i82_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4__45_i82_0_NO_SHIFT_REG = rnode_184to185_bb4__45_i82_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4__45_i82_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4__45_i82_1_NO_SHIFT_REG = rnode_184to185_bb4__45_i82_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4__45_i82_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb4__45_i82_2_NO_SHIFT_REG = rnode_184to185_bb4__45_i82_0_reg_185_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i_0_valid_out_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i_0_stall_in_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb4_not_cmp37_i_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb4_not_cmp37_i_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb4_not_cmp37_i_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb4_not_cmp37_i_0_stall_in_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb4_not_cmp37_i_0_valid_out_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb4_not_cmp37_i_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp37_i),
	.data_out(rnode_184to185_bb4_not_cmp37_i_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb4_not_cmp37_i_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb4_not_cmp37_i_0_reg_185_fifo.DATA_WIDTH = 1;
defparam rnode_184to185_bb4_not_cmp37_i_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb4_not_cmp37_i_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb4_not_cmp37_i_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp37_i_stall_in_1 = 1'b0;
assign rnode_184to185_bb4_not_cmp37_i_0_NO_SHIFT_REG = rnode_184to185_bb4_not_cmp37_i_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb4_not_cmp37_i_0_stall_in_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or276_i_stall_local;
wire [31:0] local_bb4_or276_i;

assign local_bb4_or276_i = ((local_bb4_or275_i & 32'h7FFFFFFF) | (rnode_183to184_bb4_resultSign_0_i_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u50_stall_local;
wire [31:0] local_bb4_var__u50;

assign local_bb4_var__u50[31:1] = 31'h0;
assign local_bb4_var__u50[0] = rnode_183to184_bb4__47_i_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2814_i_stall_local;
wire local_bb4_or2814_i;

assign local_bb4_or2814_i = (rnode_183to184_bb4__47_i_0_NO_SHIFT_REG | rnode_183to184_bb4_or2672_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2885_i_stall_local;
wire local_bb4_or2885_i;

assign local_bb4_or2885_i = (rnode_183to184_bb4_or2672_i_1_NO_SHIFT_REG | rnode_183to184_bb4__26_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u51_stall_local;
wire [31:0] local_bb4_var__u51;

assign local_bb4_var__u51[31:1] = 31'h0;
assign local_bb4_var__u51[0] = rnode_183to184_bb4_or2672_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i235_stall_local;
wire [31:0] local_bb4_resultSign_0_i235;

assign local_bb4_resultSign_0_i235 = (local_bb4_brmerge12_i234 ? (rnode_184to185_bb4_and35_i118_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i235_valid_out;
wire local_bb4_resultSign_0_i235_stall_in;
wire local_bb4__47_i245_valid_out;
wire local_bb4__47_i245_stall_in;
wire local_bb4_or2662_i248_valid_out;
wire local_bb4_or2662_i248_stall_in;
wire local_bb4_or2662_i248_inputs_ready;
wire local_bb4_or2662_i248_stall_local;
wire local_bb4_or2662_i248;

assign local_bb4_or2662_i248_inputs_ready = (rnode_184to185_bb4_and35_i118_0_valid_out_NO_SHIFT_REG & rnode_184to185_bb4_not_cmp37_i226_0_valid_out_NO_SHIFT_REG & rnode_184to185_bb4_add245_i238_0_valid_out_0_NO_SHIFT_REG & rnode_184to185_bb4_and250_i241_0_valid_out_NO_SHIFT_REG & rnode_184to185_bb4__45_i230_0_valid_out_0_NO_SHIFT_REG & rnode_184to185_bb4_add245_i238_0_valid_out_1_NO_SHIFT_REG & rnode_184to185_bb4_var__u31_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2662_i248 = (rnode_184to185_bb4_var__u31_0_NO_SHIFT_REG | local_bb4_lnot262__i247);
assign local_bb4_resultSign_0_i235_valid_out = 1'b1;
assign local_bb4__47_i245_valid_out = 1'b1;
assign local_bb4_or2662_i248_valid_out = 1'b1;
assign rnode_184to185_bb4_and35_i118_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_not_cmp37_i226_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_add245_i238_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and250_i241_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4__45_i230_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_add245_i238_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_var__u31_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i87_stall_local;
wire local_bb4_notrhs_i87;

assign local_bb4_notrhs_i87 = ((rnode_184to185_bb4_and250_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl273_i_stall_local;
wire [31:0] local_bb4_shl273_i;

assign local_bb4_shl273_i = ((rnode_184to186_bb4_and269_i_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and247_i_stall_local;
wire [31:0] local_bb4_and247_i;

assign local_bb4_and247_i = (rnode_184to185_bb4_add245_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp258_i_stall_local;
wire local_bb4_cmp258_i;

assign local_bb4_cmp258_i = ($signed(rnode_184to185_bb4_add245_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and225_i_stall_local;
wire [31:0] local_bb4_and225_i;

assign local_bb4_and225_i = ((rnode_184to185_bb4__45_i82_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i90_stall_local;
wire [31:0] local_bb4_and270_i90;

assign local_bb4_and270_i90 = ((rnode_184to185_bb4__45_i82_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr271_i_valid_out;
wire local_bb4_shr271_i_stall_in;
wire local_bb4_shr271_i_inputs_ready;
wire local_bb4_shr271_i_stall_local;
wire [31:0] local_bb4_shr271_i;

assign local_bb4_shr271_i_inputs_ready = rnode_184to185_bb4__45_i82_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr271_i = ((rnode_184to185_bb4__45_i82_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr271_i_valid_out = 1'b1;
assign rnode_184to185_bb4__45_i82_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext315_i_stall_local;
wire [31:0] local_bb4_lnot_ext315_i;

assign local_bb4_lnot_ext315_i = ((local_bb4_var__u50 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond283_i_stall_local;
wire [31:0] local_bb4_cond283_i;

assign local_bb4_cond283_i = (local_bb4_or2814_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond290_i_stall_local;
wire [31:0] local_bb4_cond290_i;

assign local_bb4_cond290_i = (local_bb4_or2885_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext311_i_stall_local;
wire [31:0] local_bb4_lnot_ext311_i;

assign local_bb4_lnot_ext311_i = ((local_bb4_var__u51 & 32'h1) ^ 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_resultSign_0_i235_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i235_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_resultSign_0_i235_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i235_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_resultSign_0_i235_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i235_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i235_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i235_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_resultSign_0_i235_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_resultSign_0_i235_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_resultSign_0_i235_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_resultSign_0_i235_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_resultSign_0_i235_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i235 & 32'h80000000)),
	.data_out(rnode_185to186_bb4_resultSign_0_i235_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_resultSign_0_i235_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_resultSign_0_i235_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb4_resultSign_0_i235_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_resultSign_0_i235_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_resultSign_0_i235_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i235_stall_in = 1'b0;
assign rnode_185to186_bb4_resultSign_0_i235_0_NO_SHIFT_REG = rnode_185to186_bb4_resultSign_0_i235_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_resultSign_0_i235_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_resultSign_0_i235_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4__47_i245_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i245_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4__47_i245_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4__47_i245_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4__47_i245_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4__47_i245_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4__47_i245_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4__47_i245),
	.data_out(rnode_185to186_bb4__47_i245_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4__47_i245_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4__47_i245_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4__47_i245_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4__47_i245_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4__47_i245_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i245_stall_in = 1'b0;
assign rnode_185to186_bb4__47_i245_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__47_i245_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__47_i245_0_NO_SHIFT_REG = rnode_185to186_bb4__47_i245_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4__47_i245_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__47_i245_1_NO_SHIFT_REG = rnode_185to186_bb4__47_i245_0_reg_186_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_or2662_i248_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i248_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_or2662_i248_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_or2662_i248_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_or2662_i248_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_or2662_i248_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_or2662_i248_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4_or2662_i248),
	.data_out(rnode_185to186_bb4_or2662_i248_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_or2662_i248_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_or2662_i248_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4_or2662_i248_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_or2662_i248_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_or2662_i248_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2662_i248_stall_in = 1'b0;
assign rnode_185to186_bb4_or2662_i248_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i248_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4_or2662_i248_0_NO_SHIFT_REG = rnode_185to186_bb4_or2662_i248_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_or2662_i248_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4_or2662_i248_1_NO_SHIFT_REG = rnode_185to186_bb4_or2662_i248_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_or2662_i248_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4_or2662_i248_2_NO_SHIFT_REG = rnode_185to186_bb4_or2662_i248_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i86_stall_local;
wire local_bb4_notlhs_i86;

assign local_bb4_notlhs_i86 = ((local_bb4_and247_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_i_stall_local;
wire local_bb4_cmp226_i;

assign local_bb4_cmp226_i = ((local_bb4_and225_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i_stall_local;
wire local_bb4_cmp296_i;

assign local_bb4_cmp296_i = ((local_bb4_and270_i90 & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i_valid_out;
wire local_bb4_cmp296_i_stall_in;
wire local_bb4_cmp299_i_valid_out;
wire local_bb4_cmp299_i_stall_in;
wire local_bb4_cmp299_i_inputs_ready;
wire local_bb4_cmp299_i_stall_local;
wire local_bb4_cmp299_i;

assign local_bb4_cmp299_i_inputs_ready = rnode_184to185_bb4__45_i82_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp299_i = ((local_bb4_and270_i90 & 32'h7) == 32'h4);
assign local_bb4_cmp296_i_valid_out = 1'b1;
assign local_bb4_cmp299_i_valid_out = 1'b1;
assign rnode_184to185_bb4__45_i82_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_shr271_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_shr271_i_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_shr271_i_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_shr271_i_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_shr271_i_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_shr271_i_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_shr271_i_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_shr271_i_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_shr271_i_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in((local_bb4_shr271_i & 32'h1FFFFFF)),
	.data_out(rnode_185to186_bb4_shr271_i_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_shr271_i_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_shr271_i_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb4_shr271_i_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_shr271_i_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_shr271_i_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr271_i_stall_in = 1'b0;
assign rnode_185to186_bb4_shr271_i_0_NO_SHIFT_REG = rnode_185to186_bb4_shr271_i_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_shr271_i_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_shr271_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and294_i_stall_local;
wire [31:0] local_bb4_and294_i;

assign local_bb4_and294_i = ((local_bb4_cond283_i | 32'h80000000) & local_bb4_or276_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i_stall_local;
wire [31:0] local_bb4_or295_i;

assign local_bb4_or295_i = ((local_bb4_cond290_i & 32'h7F800000) | (local_bb4_cond293_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i_stall_local;
wire [31:0] local_bb4_reduction_0_i;

assign local_bb4_reduction_0_i = ((local_bb4_lnot_ext311_i & 32'h1) & (local_bb4_lnot_ext_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i255_stall_local;
wire [31:0] local_bb4_or275_i255;

assign local_bb4_or275_i255 = ((local_bb4_or274_i254 & 32'h7FFFFFFF) | (rnode_185to186_bb4_resultSign_0_i235_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u52_stall_local;
wire [31:0] local_bb4_var__u52;

assign local_bb4_var__u52[31:1] = 31'h0;
assign local_bb4_var__u52[0] = rnode_185to186_bb4__47_i245_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2804_i256_stall_local;
wire local_bb4_or2804_i256;

assign local_bb4_or2804_i256 = (rnode_185to186_bb4__47_i245_0_NO_SHIFT_REG | rnode_185to186_bb4_or2662_i248_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2875_i258_stall_local;
wire local_bb4_or2875_i258;

assign local_bb4_or2875_i258 = (rnode_185to186_bb4_or2662_i248_1_NO_SHIFT_REG | rnode_185to186_bb4__26_i133_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u53_stall_local;
wire [31:0] local_bb4_var__u53;

assign local_bb4_var__u53[31:1] = 31'h0;
assign local_bb4_var__u53[0] = rnode_185to186_bb4_or2662_i248_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i88_stall_local;
wire local_bb4_not__46_i88;

assign local_bb4_not__46_i88 = (local_bb4_notrhs_i87 | local_bb4_notlhs_i86);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_not_i_stall_local;
wire local_bb4_cmp226_not_i;

assign local_bb4_cmp226_not_i = (local_bb4_cmp226_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp296_i_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_cmp296_i_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_cmp296_i_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_cmp296_i_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_cmp296_i_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_cmp296_i_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4_cmp296_i),
	.data_out(rnode_185to186_bb4_cmp296_i_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_cmp296_i_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_cmp296_i_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4_cmp296_i_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_cmp296_i_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_cmp296_i_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp296_i_stall_in = 1'b0;
assign rnode_185to186_bb4_cmp296_i_0_NO_SHIFT_REG = rnode_185to186_bb4_cmp296_i_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_cmp296_i_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_cmp299_i_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_cmp299_i_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_cmp299_i_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_cmp299_i_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_cmp299_i_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_cmp299_i_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4_cmp299_i),
	.data_out(rnode_185to186_bb4_cmp299_i_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_cmp299_i_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_cmp299_i_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4_cmp299_i_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_cmp299_i_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_cmp299_i_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp299_i_stall_in = 1'b0;
assign rnode_185to186_bb4_cmp299_i_0_NO_SHIFT_REG = rnode_185to186_bb4_cmp299_i_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_cmp299_i_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and272_i_stall_local;
wire [31:0] local_bb4_and272_i;

assign local_bb4_and272_i = ((rnode_185to186_bb4_shr271_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and303_i_stall_local;
wire [31:0] local_bb4_and303_i;

assign local_bb4_and303_i = ((local_bb4_conv301_i & 32'h1) & local_bb4_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or296_i_stall_local;
wire [31:0] local_bb4_or296_i;

assign local_bb4_or296_i = ((local_bb4_or295_i & 32'h7FC00000) | local_bb4_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext314_i272_stall_local;
wire [31:0] local_bb4_lnot_ext314_i272;

assign local_bb4_lnot_ext314_i272 = ((local_bb4_var__u52 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond282_i257_stall_local;
wire [31:0] local_bb4_cond282_i257;

assign local_bb4_cond282_i257 = (local_bb4_or2804_i256 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond289_i259_stall_local;
wire [31:0] local_bb4_cond289_i259;

assign local_bb4_cond289_i259 = (local_bb4_or2875_i258 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext310_i271_stall_local;
wire [31:0] local_bb4_lnot_ext310_i271;

assign local_bb4_lnot_ext310_i271 = ((local_bb4_var__u53 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__47_i89_stall_local;
wire local_bb4__47_i89;

assign local_bb4__47_i89 = (local_bb4_cmp226_i | local_bb4_not__46_i88);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i83_stall_local;
wire local_bb4_brmerge12_i83;

assign local_bb4_brmerge12_i83 = (local_bb4_cmp226_not_i | rnode_184to185_bb4_not_cmp37_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot262__i_stall_local;
wire local_bb4_lnot262__i;

assign local_bb4_lnot262__i = (local_bb4_cmp258_i & local_bb4_cmp226_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29649_i_stall_local;
wire [31:0] local_bb4_cmp29649_i;

assign local_bb4_cmp29649_i[31:1] = 31'h0;
assign local_bb4_cmp29649_i[0] = rnode_185to186_bb4_cmp296_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv300_i_stall_local;
wire [31:0] local_bb4_conv300_i;

assign local_bb4_conv300_i[31:1] = 31'h0;
assign local_bb4_conv300_i[0] = rnode_185to186_bb4_cmp299_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or274_i_stall_local;
wire [31:0] local_bb4_or274_i;

assign local_bb4_or274_i = ((local_bb4_and272_i & 32'h7FFFFF) | (local_bb4_shl273_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i_stall_local;
wire [31:0] local_bb4_lor_ext_i;

assign local_bb4_lor_ext_i = ((local_bb4_cmp29749_i & 32'h1) | (local_bb4_and303_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and293_i261_stall_local;
wire [31:0] local_bb4_and293_i261;

assign local_bb4_and293_i261 = ((local_bb4_cond282_i257 | 32'h80000000) & local_bb4_or275_i255);

// This section implements an unregistered operation.
// 
wire local_bb4_or294_i262_stall_local;
wire [31:0] local_bb4_or294_i262;

assign local_bb4_or294_i262 = ((local_bb4_cond289_i259 & 32'h7F800000) | (local_bb4_cond292_i260 & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i273_stall_local;
wire [31:0] local_bb4_reduction_0_i273;

assign local_bb4_reduction_0_i273 = ((local_bb4_lnot_ext310_i271 & 32'h1) & (local_bb4_lnot_ext_i270 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i84_stall_local;
wire [31:0] local_bb4_resultSign_0_i84;

assign local_bb4_resultSign_0_i84 = (local_bb4_brmerge12_i83 ? (rnode_184to185_bb4_and35_i25_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i84_valid_out;
wire local_bb4_resultSign_0_i84_stall_in;
wire local_bb4__47_i89_valid_out;
wire local_bb4__47_i89_stall_in;
wire local_bb4_or2662_i_valid_out;
wire local_bb4_or2662_i_stall_in;
wire local_bb4_or2662_i_inputs_ready;
wire local_bb4_or2662_i_stall_local;
wire local_bb4_or2662_i;

assign local_bb4_or2662_i_inputs_ready = (rnode_184to185_bb4_and35_i25_0_valid_out_NO_SHIFT_REG & rnode_184to185_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG & rnode_184to185_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG & rnode_184to185_bb4_and250_i_0_valid_out_NO_SHIFT_REG & rnode_184to185_bb4__45_i82_0_valid_out_0_NO_SHIFT_REG & rnode_184to185_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG & rnode_184to185_bb4_var__u39_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2662_i = (rnode_184to185_bb4_var__u39_0_NO_SHIFT_REG | local_bb4_lnot262__i);
assign local_bb4_resultSign_0_i84_valid_out = 1'b1;
assign local_bb4__47_i89_valid_out = 1'b1;
assign local_bb4_or2662_i_valid_out = 1'b1;
assign rnode_184to185_bb4_and35_i25_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_not_cmp37_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_add245_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_and250_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4__45_i82_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_add245_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb4_var__u39_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i_stall_local;
wire [31:0] local_bb4_reduction_1_i;

assign local_bb4_reduction_1_i = ((local_bb4_lnot_ext315_i & 32'h1) & (local_bb4_lor_ext_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and302_i267_stall_local;
wire [31:0] local_bb4_and302_i267;

assign local_bb4_and302_i267 = ((local_bb4_conv300_i266 & 32'h1) & local_bb4_and293_i261);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i263_stall_local;
wire [31:0] local_bb4_or295_i263;

assign local_bb4_or295_i263 = ((local_bb4_or294_i262 & 32'h7FC00000) | local_bb4_and293_i261);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_resultSign_0_i84_0_valid_out_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i84_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_resultSign_0_i84_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i84_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb4_resultSign_0_i84_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i84_0_valid_out_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i84_0_stall_in_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_resultSign_0_i84_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_resultSign_0_i84_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_resultSign_0_i84_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_resultSign_0_i84_0_stall_in_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_resultSign_0_i84_0_valid_out_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_resultSign_0_i84_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i84 & 32'h80000000)),
	.data_out(rnode_185to186_bb4_resultSign_0_i84_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_resultSign_0_i84_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_resultSign_0_i84_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb4_resultSign_0_i84_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_resultSign_0_i84_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_resultSign_0_i84_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i84_stall_in = 1'b0;
assign rnode_185to186_bb4_resultSign_0_i84_0_NO_SHIFT_REG = rnode_185to186_bb4_resultSign_0_i84_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_resultSign_0_i84_0_stall_in_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_resultSign_0_i84_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4__47_i89_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4__47_i89_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4__47_i89_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4__47_i89_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4__47_i89_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4__47_i89_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4__47_i89_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4__47_i89),
	.data_out(rnode_185to186_bb4__47_i89_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4__47_i89_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4__47_i89_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4__47_i89_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4__47_i89_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4__47_i89_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i89_stall_in = 1'b0;
assign rnode_185to186_bb4__47_i89_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__47_i89_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__47_i89_0_NO_SHIFT_REG = rnode_185to186_bb4__47_i89_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4__47_i89_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4__47_i89_1_NO_SHIFT_REG = rnode_185to186_bb4__47_i89_0_reg_186_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_1_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_2_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb4_or2662_i_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb4_or2662_i_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb4_or2662_i_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb4_or2662_i_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb4_or2662_i_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb4_or2662_i_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb4_or2662_i),
	.data_out(rnode_185to186_bb4_or2662_i_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb4_or2662_i_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb4_or2662_i_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb4_or2662_i_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb4_or2662_i_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb4_or2662_i_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2662_i_stall_in = 1'b0;
assign rnode_185to186_bb4_or2662_i_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4_or2662_i_0_NO_SHIFT_REG = rnode_185to186_bb4_or2662_i_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4_or2662_i_1_NO_SHIFT_REG = rnode_185to186_bb4_or2662_i_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb4_or2662_i_2_NO_SHIFT_REG = rnode_185to186_bb4_or2662_i_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i_stall_local;
wire [31:0] local_bb4_reduction_2_i;

assign local_bb4_reduction_2_i = ((local_bb4_reduction_0_i & 32'h1) & (local_bb4_reduction_1_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i269_stall_local;
wire [31:0] local_bb4_lor_ext_i269;

assign local_bb4_lor_ext_i269 = ((local_bb4_cmp29649_i268 & 32'h1) | (local_bb4_and302_i267 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i91_stall_local;
wire [31:0] local_bb4_or275_i91;

assign local_bb4_or275_i91 = ((local_bb4_or274_i & 32'h7FFFFFFF) | (rnode_185to186_bb4_resultSign_0_i84_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u54_stall_local;
wire [31:0] local_bb4_var__u54;

assign local_bb4_var__u54[31:1] = 31'h0;
assign local_bb4_var__u54[0] = rnode_185to186_bb4__47_i89_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2804_i_stall_local;
wire local_bb4_or2804_i;

assign local_bb4_or2804_i = (rnode_185to186_bb4__47_i89_0_NO_SHIFT_REG | rnode_185to186_bb4_or2662_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2875_i_stall_local;
wire local_bb4_or2875_i;

assign local_bb4_or2875_i = (rnode_185to186_bb4_or2662_i_1_NO_SHIFT_REG | rnode_185to186_bb4__26_i39_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u55_stall_local;
wire [31:0] local_bb4_var__u55;

assign local_bb4_var__u55[31:1] = 31'h0;
assign local_bb4_var__u55[0] = rnode_185to186_bb4_or2662_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add321_i_stall_local;
wire [31:0] local_bb4_add321_i;

assign local_bb4_add321_i = ((local_bb4_reduction_2_i & 32'h1) + local_bb4_or296_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i274_stall_local;
wire [31:0] local_bb4_reduction_1_i274;

assign local_bb4_reduction_1_i274 = ((local_bb4_lnot_ext314_i272 & 32'h1) & (local_bb4_lor_ext_i269 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext314_i_stall_local;
wire [31:0] local_bb4_lnot_ext314_i;

assign local_bb4_lnot_ext314_i = ((local_bb4_var__u54 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond282_i_stall_local;
wire [31:0] local_bb4_cond282_i;

assign local_bb4_cond282_i = (local_bb4_or2804_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond289_i_stall_local;
wire [31:0] local_bb4_cond289_i;

assign local_bb4_cond289_i = (local_bb4_or2875_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext310_i_stall_local;
wire [31:0] local_bb4_lnot_ext310_i;

assign local_bb4_lnot_ext310_i = ((local_bb4_var__u55 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i_stall_local;
wire [31:0] local_bb4_and_i_i;

assign local_bb4_and_i_i = (local_bb4_add321_i & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i275_stall_local;
wire [31:0] local_bb4_reduction_2_i275;

assign local_bb4_reduction_2_i275 = ((local_bb4_reduction_0_i273 & 32'h1) & (local_bb4_reduction_1_i274 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and293_i_stall_local;
wire [31:0] local_bb4_and293_i;

assign local_bb4_and293_i = ((local_bb4_cond282_i | 32'h80000000) & local_bb4_or275_i91);

// This section implements an unregistered operation.
// 
wire local_bb4_or294_i_stall_local;
wire [31:0] local_bb4_or294_i;

assign local_bb4_or294_i = ((local_bb4_cond289_i & 32'h7F800000) | (local_bb4_cond292_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i95_stall_local;
wire [31:0] local_bb4_reduction_0_i95;

assign local_bb4_reduction_0_i95 = ((local_bb4_lnot_ext310_i & 32'h1) & (local_bb4_lnot_ext_i94 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_astype1_i_i_valid_out;
wire local_bb4_astype1_i_i_stall_in;
wire local_bb4_astype1_i_i_inputs_ready;
wire local_bb4_astype1_i_i_stall_local;
wire [31:0] local_bb4_astype1_i_i;

assign local_bb4_astype1_i_i_inputs_ready = (rnode_182to184_bb4_and270_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4__26_i_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4__26_i_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4__47_i_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4__26_i_0_valid_out_2_NO_SHIFT_REG & rnode_183to184_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG & rnode_183to184_bb4_shr272_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4__47_i_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_astype1_i_i = (local_bb4_and_i_i & 32'h7FFFFFFF);
assign local_bb4_astype1_i_i_valid_out = 1'b1;
assign rnode_182to184_bb4_and270_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_resultSign_0_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__47_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_shr272_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__47_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp297_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp300_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_add320_i276_valid_out;
wire local_bb4_add320_i276_stall_in;
wire local_bb4_add320_i276_inputs_ready;
wire local_bb4_add320_i276_stall_local;
wire [31:0] local_bb4_add320_i276;

assign local_bb4_add320_i276_inputs_ready = (rnode_184to186_bb4_and269_i252_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4_resultSign_0_i235_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4_or2662_i248_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb4__26_i133_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb4__26_i133_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb4__47_i245_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb4_or2662_i248_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb4__26_i133_0_valid_out_2_NO_SHIFT_REG & rnode_185to186_bb4_or2662_i248_0_valid_out_2_NO_SHIFT_REG & rnode_185to186_bb4_shr271_i250_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4__47_i245_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb4_cmp296_i264_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4_cmp299_i265_0_valid_out_NO_SHIFT_REG);
assign local_bb4_add320_i276 = ((local_bb4_reduction_2_i275 & 32'h1) + local_bb4_or295_i263);
assign local_bb4_add320_i276_valid_out = 1'b1;
assign rnode_184to186_bb4_and269_i252_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_resultSign_0_i235_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i248_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i133_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i133_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__47_i245_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i248_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i133_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i248_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_shr271_i250_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__47_i245_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp296_i264_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp299_i265_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and302_i_stall_local;
wire [31:0] local_bb4_and302_i;

assign local_bb4_and302_i = ((local_bb4_conv300_i & 32'h1) & local_bb4_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i92_stall_local;
wire [31:0] local_bb4_or295_i92;

assign local_bb4_or295_i92 = ((local_bb4_or294_i & 32'h7FC00000) | local_bb4_and293_i);

// This section implements a registered operation.
// 
wire local_bb4_cmp30_inputs_ready;
 reg local_bb4_cmp30_valid_out_0_NO_SHIFT_REG;
wire local_bb4_cmp30_stall_in_0;
 reg local_bb4_cmp30_valid_out_1_NO_SHIFT_REG;
wire local_bb4_cmp30_stall_in_1;
wire local_bb4_cmp30_output_regs_ready;
wire local_bb4_cmp30;
 reg local_bb4_cmp30_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_cmp30_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_cmp30_causedstall;

acl_fp_cmp fp_module_local_bb4_cmp30 (
	.clock(clock),
	.dataa(local_bb4_astype1_i_i),
	.datab(input_e_d),
	.enable(local_bb4_cmp30_output_regs_ready),
	.result(local_bb4_cmp30)
);

defparam fp_module_local_bb4_cmp30.COMPARISON_MODE = 5;

assign local_bb4_cmp30_inputs_ready = 1'b1;
assign local_bb4_cmp30_output_regs_ready = 1'b1;
assign local_bb4_astype1_i_i_stall_in = 1'b0;
assign local_bb4_cmp30_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_cmp30_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_cmp30_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_cmp30_output_regs_ready)
		begin
			local_bb4_cmp30_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_cmp30_valid_pipe_1_NO_SHIFT_REG <= local_bb4_cmp30_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_cmp30_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_cmp30_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_cmp30_output_regs_ready)
		begin
			local_bb4_cmp30_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_cmp30_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_cmp30_stall_in_0))
			begin
				local_bb4_cmp30_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_cmp30_stall_in_1))
			begin
				local_bb4_cmp30_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb4_add320_i276_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i276_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_add320_i276_0_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i276_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_add320_i276_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i276_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i276_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i276_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb4_add320_i276_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb4_add320_i276_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb4_add320_i276_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb4_add320_i276_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb4_add320_i276_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb4_add320_i276),
	.data_out(rnode_186to187_bb4_add320_i276_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb4_add320_i276_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb4_add320_i276_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb4_add320_i276_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb4_add320_i276_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb4_add320_i276_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add320_i276_stall_in = 1'b0;
assign rnode_186to187_bb4_add320_i276_0_NO_SHIFT_REG = rnode_186to187_bb4_add320_i276_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb4_add320_i276_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_add320_i276_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i93_stall_local;
wire [31:0] local_bb4_lor_ext_i93;

assign local_bb4_lor_ext_i93 = ((local_bb4_cmp29649_i & 32'h1) | (local_bb4_and302_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u56_stall_local;
wire [31:0] local_bb4_var__u56;

assign local_bb4_var__u56 = rnode_186to187_bb4_add320_i276_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i96_stall_local;
wire [31:0] local_bb4_reduction_1_i96;

assign local_bb4_reduction_1_i96 = ((local_bb4_lnot_ext314_i & 32'h1) & (local_bb4_lor_ext_i93 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__23_stall_local;
wire [31:0] local_bb4__23;

assign local_bb4__23 = (local_bb4_cmp30 ? local_bb4_var__u56 : rnode_186to187_bb4_sum_33_pop32__0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i97_stall_local;
wire [31:0] local_bb4_reduction_2_i97;

assign local_bb4_reduction_2_i97 = ((local_bb4_reduction_0_i95 & 32'h1) & (local_bb4_reduction_1_i96 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__23_valid_out_0;
wire local_bb4__23_stall_in_0;
wire local_bb4_select28_valid_out;
wire local_bb4_select28_stall_in;
wire local_bb4_select28_inputs_ready;
wire local_bb4_select28_stall_local;
wire [31:0] local_bb4_select28;

assign local_bb4_select28_inputs_ready = (local_bb4_cmp30_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb4_sum_33_pop32__0_valid_out_NO_SHIFT_REG & rnode_186to187_bb4_add320_i276_0_valid_out_NO_SHIFT_REG);
assign local_bb4_select28 = (input_wii_var__u17 ? 32'h0 : local_bb4__23);
assign local_bb4__23_valid_out_0 = 1'b1;
assign local_bb4_select28_valid_out = 1'b1;
assign local_bb4_cmp30_stall_in_0 = 1'b0;
assign rnode_186to187_bb4_sum_33_pop32__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_add320_i276_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_add320_i_valid_out;
wire local_bb4_add320_i_stall_in;
wire local_bb4_add320_i_inputs_ready;
wire local_bb4_add320_i_stall_local;
wire [31:0] local_bb4_add320_i;

assign local_bb4_add320_i_inputs_ready = (rnode_184to186_bb4_and269_i_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4_resultSign_0_i84_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb4__26_i39_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb4__26_i39_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb4__47_i89_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb4__26_i39_0_valid_out_2_NO_SHIFT_REG & rnode_185to186_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG & rnode_185to186_bb4_shr271_i_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4__47_i89_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG & rnode_185to186_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_add320_i = ((local_bb4_reduction_2_i97 & 32'h1) + local_bb4_or295_i92);
assign local_bb4_add320_i_valid_out = 1'b1;
assign rnode_184to186_bb4_and269_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_resultSign_0_i84_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i39_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i39_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__47_i89_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__26_i39_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_or2662_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_shr271_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4__47_i89_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp296_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb4_cmp299_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_sum_33_push32__23_inputs_ready;
 reg local_bb4_sum_33_push32__23_valid_out_NO_SHIFT_REG;
wire local_bb4_sum_33_push32__23_stall_in;
wire local_bb4_sum_33_push32__23_output_regs_ready;
wire [31:0] local_bb4_sum_33_push32__23_result;
wire local_bb4_sum_33_push32__23_fu_valid_out;
wire local_bb4_sum_33_push32__23_fu_stall_out;
 reg [31:0] local_bb4_sum_33_push32__23_NO_SHIFT_REG;
wire local_bb4_sum_33_push32__23_causedstall;

acl_push local_bb4_sum_33_push32__23_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_186to187_bb4_notexitcond_or_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4__23),
	.stall_out(local_bb4_sum_33_push32__23_fu_stall_out),
	.valid_in(SFC_3_VALID_186_187_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sum_33_push32__23_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_sum_33_push32__23_result),
	.feedback_out(feedback_data_out_32),
	.feedback_valid_out(feedback_valid_out_32),
	.feedback_stall_in(feedback_stall_in_32)
);

defparam local_bb4_sum_33_push32__23_feedback.STALLFREE = 1;
defparam local_bb4_sum_33_push32__23_feedback.DATA_WIDTH = 32;
defparam local_bb4_sum_33_push32__23_feedback.FIFO_DEPTH = 9;
defparam local_bb4_sum_33_push32__23_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb4_sum_33_push32__23_feedback.STYLE = "REGULAR";

assign local_bb4_sum_33_push32__23_inputs_ready = 1'b1;
assign local_bb4_sum_33_push32__23_output_regs_ready = 1'b1;
assign local_bb4__23_stall_in_0 = 1'b0;
assign SFC_3_VALID_186_187_0_stall_in_1 = 1'b0;
assign rnode_186to187_bb4_notexitcond_or_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb4_sum_33_push32__23_causedstall = (SFC_3_VALID_186_187_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_sum_33_push32__23_NO_SHIFT_REG <= 'x;
		local_bb4_sum_33_push32__23_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_sum_33_push32__23_output_regs_ready)
		begin
			local_bb4_sum_33_push32__23_NO_SHIFT_REG <= local_bb4_sum_33_push32__23_result;
			local_bb4_sum_33_push32__23_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_sum_33_push32__23_stall_in))
			begin
				local_bb4_sum_33_push32__23_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb4_select28_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select28_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb4_select28_0_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select28_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb4_select28_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select28_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select28_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select28_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb4_select28_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb4_select28_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb4_select28_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb4_select28_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb4_select28_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb4_select28),
	.data_out(rnode_187to188_bb4_select28_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb4_select28_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb4_select28_0_reg_188_fifo.DATA_WIDTH = 32;
defparam rnode_187to188_bb4_select28_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb4_select28_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb4_select28_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_select28_stall_in = 1'b0;
assign rnode_187to188_bb4_select28_0_NO_SHIFT_REG = rnode_187to188_bb4_select28_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb4_select28_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb4_select28_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb4_add320_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_add320_i_0_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb4_add320_i_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb4_add320_i_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb4_add320_i_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb4_add320_i_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb4_add320_i_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb4_add320_i_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb4_add320_i_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb4_add320_i),
	.data_out(rnode_186to187_bb4_add320_i_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb4_add320_i_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb4_add320_i_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb4_add320_i_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb4_add320_i_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb4_add320_i_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add320_i_stall_in = 1'b0;
assign rnode_186to187_bb4_add320_i_0_NO_SHIFT_REG = rnode_186to187_bb4_add320_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb4_add320_i_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_add320_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u57_stall_local;
wire [31:0] local_bb4_var__u57;

assign local_bb4_var__u57 = rnode_186to187_bb4_add320_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__24_stall_local;
wire [31:0] local_bb4__24;

assign local_bb4__24 = (local_bb4_cmp30 ? local_bb4_var__u57 : rnode_186to187_bb4_t_34_pop31__0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__24_valid_out_0;
wire local_bb4__24_stall_in_0;
wire local_bb4_select25_valid_out;
wire local_bb4_select25_stall_in;
wire local_bb4_select25_inputs_ready;
wire local_bb4_select25_stall_local;
wire [31:0] local_bb4_select25;

assign local_bb4_select25_inputs_ready = (local_bb4_cmp30_valid_out_1_NO_SHIFT_REG & rnode_186to187_bb4_t_34_pop31__0_valid_out_NO_SHIFT_REG & rnode_186to187_bb4_add320_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_select25 = (input_wii_var__u17 ? 32'h0 : local_bb4__24);
assign local_bb4__24_valid_out_0 = 1'b1;
assign local_bb4_select25_valid_out = 1'b1;
assign local_bb4_cmp30_stall_in_1 = 1'b0;
assign rnode_186to187_bb4_t_34_pop31__0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb4_add320_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_t_34_push31__24_inputs_ready;
 reg local_bb4_t_34_push31__24_valid_out_NO_SHIFT_REG;
wire local_bb4_t_34_push31__24_stall_in;
wire local_bb4_t_34_push31__24_output_regs_ready;
wire [31:0] local_bb4_t_34_push31__24_result;
wire local_bb4_t_34_push31__24_fu_valid_out;
wire local_bb4_t_34_push31__24_fu_stall_out;
 reg [31:0] local_bb4_t_34_push31__24_NO_SHIFT_REG;
wire local_bb4_t_34_push31__24_causedstall;

acl_push local_bb4_t_34_push31__24_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_186to187_bb4_notexitcond_or_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4__24),
	.stall_out(local_bb4_t_34_push31__24_fu_stall_out),
	.valid_in(SFC_3_VALID_186_187_0_NO_SHIFT_REG),
	.valid_out(local_bb4_t_34_push31__24_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_t_34_push31__24_result),
	.feedback_out(feedback_data_out_31),
	.feedback_valid_out(feedback_valid_out_31),
	.feedback_stall_in(feedback_stall_in_31)
);

defparam local_bb4_t_34_push31__24_feedback.STALLFREE = 1;
defparam local_bb4_t_34_push31__24_feedback.DATA_WIDTH = 32;
defparam local_bb4_t_34_push31__24_feedback.FIFO_DEPTH = 9;
defparam local_bb4_t_34_push31__24_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_t_34_push31__24_feedback.STYLE = "REGULAR";

assign local_bb4_t_34_push31__24_inputs_ready = 1'b1;
assign local_bb4_t_34_push31__24_output_regs_ready = 1'b1;
assign local_bb4__24_stall_in_0 = 1'b0;
assign SFC_3_VALID_186_187_0_stall_in_2 = 1'b0;
assign rnode_186to187_bb4_notexitcond_or_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign local_bb4_t_34_push31__24_causedstall = (SFC_3_VALID_186_187_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_t_34_push31__24_NO_SHIFT_REG <= 'x;
		local_bb4_t_34_push31__24_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_t_34_push31__24_output_regs_ready)
		begin
			local_bb4_t_34_push31__24_NO_SHIFT_REG <= local_bb4_t_34_push31__24_result;
			local_bb4_t_34_push31__24_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_t_34_push31__24_stall_in))
			begin
				local_bb4_t_34_push31__24_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb4_select25_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb4_select25_0_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select25_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb4_select25_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select25_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select25_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb4_select25_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb4_select25_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb4_select25_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb4_select25_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb4_select25_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb4_select25_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb4_select25),
	.data_out(rnode_187to188_bb4_select25_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb4_select25_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb4_select25_0_reg_188_fifo.DATA_WIDTH = 32;
defparam rnode_187to188_bb4_select25_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb4_select25_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb4_select25_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_select25_stall_in = 1'b0;
assign rnode_187to188_bb4_select25_0_NO_SHIFT_REG = rnode_187to188_bb4_select25_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb4_select25_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb4_select25_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_exi1_stall_local;
wire [95:0] local_bb4_c1_exi1;

assign local_bb4_c1_exi1[31:0] = 32'bx;
assign local_bb4_c1_exi1[63:32] = rnode_187to188_bb4_select25_0_NO_SHIFT_REG;
assign local_bb4_c1_exi1[95:64] = 32'bx;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_exi2_valid_out;
wire local_bb4_c1_exi2_stall_in;
wire local_bb4_c1_exi2_inputs_ready;
wire local_bb4_c1_exi2_stall_local;
wire [95:0] local_bb4_c1_exi2;

assign local_bb4_c1_exi2_inputs_ready = (rnode_187to188_bb4_select28_0_valid_out_NO_SHIFT_REG & rnode_187to188_bb4_select25_0_valid_out_NO_SHIFT_REG);
assign local_bb4_c1_exi2[63:0] = local_bb4_c1_exi1[63:0];
assign local_bb4_c1_exi2[95:64] = rnode_187to188_bb4_select28_0_NO_SHIFT_REG;
assign local_bb4_c1_exi2_valid_out = 1'b1;
assign rnode_187to188_bb4_select28_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb4_select25_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_c1_exit_c1_exi2_inputs_ready;
 reg local_bb4_c1_exit_c1_exi2_valid_out_0_NO_SHIFT_REG;
wire local_bb4_c1_exit_c1_exi2_stall_in_0;
 reg local_bb4_c1_exit_c1_exi2_valid_out_1_NO_SHIFT_REG;
wire local_bb4_c1_exit_c1_exi2_stall_in_1;
 reg [95:0] local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG;
wire [95:0] local_bb4_c1_exit_c1_exi2_in;
wire local_bb4_c1_exit_c1_exi2_valid;
wire local_bb4_c1_exit_c1_exi2_causedstall;

acl_stall_free_sink local_bb4_c1_exit_c1_exi2_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb4_c1_exi2),
	.data_out(local_bb4_c1_exit_c1_exi2_in),
	.input_accepted(local_bb4_c1_enter_c1_eni6_input_accepted),
	.valid_out(local_bb4_c1_exit_c1_exi2_valid),
	.stall_in(~(local_bb4_c1_exit_c1_exi2_output_regs_ready)),
	.stall_entry(local_bb4_c1_exit_c1_exi2_entry_stall),
	.valid_in(local_bb4_c1_exit_c1_exi2_valid_in),
	.IIphases(local_bb4_c1_exit_c1_exi2_phases),
	.inc_pipelined_thread(local_bb4_c1_enter_c1_eni6_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb4_c1_enter_c1_eni6_dec_pipelined_thread)
);

defparam local_bb4_c1_exit_c1_exi2_instance.DATA_WIDTH = 96;
defparam local_bb4_c1_exit_c1_exi2_instance.PIPELINE_DEPTH = 17;
defparam local_bb4_c1_exit_c1_exi2_instance.SHARINGII = 1;
defparam local_bb4_c1_exit_c1_exi2_instance.SCHEDULEII = 9;
defparam local_bb4_c1_exit_c1_exi2_instance.ALWAYS_THROTTLE = 1;

assign local_bb4_c1_exit_c1_exi2_inputs_ready = 1'b1;
assign local_bb4_c1_exit_c1_exi2_output_regs_ready = ((~(local_bb4_c1_exit_c1_exi2_valid_out_0_NO_SHIFT_REG) | ~(local_bb4_c1_exit_c1_exi2_stall_in_0)) & (~(local_bb4_c1_exit_c1_exi2_valid_out_1_NO_SHIFT_REG) | ~(local_bb4_c1_exit_c1_exi2_stall_in_1)));
assign local_bb4_c1_exit_c1_exi2_valid_in = SFC_3_VALID_187_188_0_NO_SHIFT_REG;
assign local_bb4_c1_exi2_stall_in = 1'b0;
assign local_bb4_sum_33_push32__23_stall_in = 1'b0;
assign local_bb4_t_34_push31__24_stall_in = 1'b0;
assign SFC_3_VALID_187_188_0_stall_in = 1'b0;
assign rnode_187to188_bb4_notexitcond546_push48_notexitcond546_pop48_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_c1_exit_c1_exi2_causedstall = (1'b1 && (1'b0 && !(~(local_bb4_c1_exit_c1_exi2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG <= 'x;
		local_bb4_c1_exit_c1_exi2_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_exit_c1_exi2_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c1_exit_c1_exi2_output_regs_ready)
		begin
			local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_in;
			local_bb4_c1_exit_c1_exi2_valid_out_0_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_valid;
			local_bb4_c1_exit_c1_exi2_valid_out_1_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_valid;
		end
		else
		begin
			if (~(local_bb4_c1_exit_c1_exi2_stall_in_0))
			begin
				local_bb4_c1_exit_c1_exi2_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_exit_c1_exi2_stall_in_1))
			begin
				local_bb4_c1_exit_c1_exi2_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_exe1_stall_local;
wire [31:0] local_bb4_c1_exe1;

assign local_bb4_c1_exe1 = local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_exe2_valid_out;
wire local_bb4_c1_exe2_stall_in;
wire local_bb4_c1_exe1_valid_out;
wire local_bb4_c1_exe1_stall_in;
wire local_bb4_c1_exe2_inputs_ready;
wire local_bb4_c1_exe2_stall_local;
wire [31:0] local_bb4_c1_exe2;

assign local_bb4_c1_exe2_inputs_ready = (local_bb4_c1_exit_c1_exi2_valid_out_1_NO_SHIFT_REG & local_bb4_c1_exit_c1_exi2_valid_out_0_NO_SHIFT_REG);
assign local_bb4_c1_exe2 = local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG[95:64];
assign local_bb4_c1_exe2_stall_local = (local_bb4_c1_exe2_stall_in | local_bb4_c1_exe1_stall_in);
assign local_bb4_c1_exe2_valid_out = local_bb4_c1_exe2_inputs_ready;
assign local_bb4_c1_exe1_valid_out = local_bb4_c1_exe2_inputs_ready;
assign local_bb4_c1_exit_c1_exi2_stall_in_1 = (local_bb4_c1_exe2_stall_local | ~(local_bb4_c1_exe2_inputs_ready));
assign local_bb4_c1_exit_c1_exi2_stall_in_0 = (local_bb4_c1_exe2_stall_local | ~(local_bb4_c1_exe2_inputs_ready));

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [447:0] lvb_bb4_c0_exit87_c0_exi1386_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb4_c0_exe794_0_reg_NO_SHIFT_REG;
 reg lvb_bb4_c0_exe895_0_reg_NO_SHIFT_REG;
 reg lvb_bb4_c0_exe996_0_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb4_c0_exe1097_0_reg_NO_SHIFT_REG;
 reg lvb_bb4_c0_exe1198_0_reg_NO_SHIFT_REG;
 reg lvb_bb4_c0_exe1299_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb4_c1_exe1_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb4_c1_exe2_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb4_c1_exe2_valid_out & local_bb4_c1_exe1_valid_out & local_bb4_c0_exe1299_valid_out & local_bb4_c0_exe1198_valid_out & local_bb4_c0_exe1097_valid_out & local_bb4_c0_exe996_valid_out & local_bb4_c0_exe895_valid_out & local_bb4_c0_exe794_valid_out & local_bb4_c0_exe592_valid_out & rnode_192to193_bb4_c0_exit87_c0_exi1386_0_valid_out_7_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb4_c1_exe2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c1_exe1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe1299_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe1198_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe1097_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe996_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe895_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe794_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe592_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_192to193_bb4_c0_exit87_c0_exi1386_0_stall_in_7_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb4_c0_exit87_c0_exi1386_0 = lvb_bb4_c0_exit87_c0_exi1386_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exit87_c0_exi1386_1 = lvb_bb4_c0_exit87_c0_exi1386_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe794_0 = lvb_bb4_c0_exe794_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe794_1 = lvb_bb4_c0_exe794_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe895_0 = lvb_bb4_c0_exe895_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe895_1 = lvb_bb4_c0_exe895_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe996_0 = lvb_bb4_c0_exe996_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe996_1 = lvb_bb4_c0_exe996_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe1097_0 = lvb_bb4_c0_exe1097_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe1097_1 = lvb_bb4_c0_exe1097_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe1198_0 = lvb_bb4_c0_exe1198_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe1198_1 = lvb_bb4_c0_exe1198_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe1299_0 = lvb_bb4_c0_exe1299_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe1299_1 = lvb_bb4_c0_exe1299_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exe1_0 = lvb_bb4_c1_exe1_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exe1_1 = lvb_bb4_c1_exe1_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exe2_0 = lvb_bb4_c1_exe2_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exe2_1 = lvb_bb4_c1_exe2_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_bb4_c0_exit87_c0_exi1386_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe794_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe895_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe996_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe1097_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe1198_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe1299_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c1_exe1_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c1_exe2_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb4_c0_exit87_c0_exi1386_0_reg_NO_SHIFT_REG <= rnode_192to193_bb4_c0_exit87_c0_exi1386_7_NO_SHIFT_REG;
			lvb_bb4_c0_exe794_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe794;
			lvb_bb4_c0_exe895_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe895;
			lvb_bb4_c0_exe996_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe996;
			lvb_bb4_c0_exe1097_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe1097;
			lvb_bb4_c0_exe1198_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe1198;
			lvb_bb4_c0_exe1299_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe1299;
			lvb_bb4_c1_exe1_0_reg_NO_SHIFT_REG <= local_bb4_c1_exe1;
			lvb_bb4_c1_exe2_0_reg_NO_SHIFT_REG <= local_bb4_c1_exe2;
			branch_compare_result_NO_SHIFT_REG <= local_bb4_c0_exe592;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_5
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_wii_div,
		input [31:0] 		input_wii_div1,
		input 		input_wii_cmp19,
		input [31:0] 		input_wii_add7,
		input [31:0] 		input_wii_sub20,
		input [31:0] 		input_wii_sub22,
		input 		input_wii_var_,
		input 		input_wii_var__u58,
		input 		input_wii_var__u59,
		input 		input_wii_var__u60,
		input 		valid_in,
		output 		stall_out,
		input [447:0] 		input_c0_exit87_c0_exi1386,
		input [31:0] 		input_c0_exe794,
		input 		input_c0_exe895,
		input 		input_c0_exe996,
		input [63:0] 		input_c0_exe1097,
		input 		input_c0_exe1198,
		input 		input_c0_exe1299,
		input [31:0] 		input_c1_exe1,
		input [31:0] 		input_c1_exe2,
		output 		valid_out_0,
		input 		stall_in_0,
		output [31:0] 		lvb_c0_exe794_0,
		output 		lvb_c0_exe895_0,
		output 		lvb_c0_exe996_0,
		output [63:0] 		lvb_c0_exe1097_0,
		output 		lvb_c0_exe1198_0,
		output 		lvb_c0_exe1299_0,
		output [31:0] 		lvb_c1_exe1_0,
		output [31:0] 		lvb_c1_exe2_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [31:0] 		lvb_c0_exe794_1,
		output 		lvb_c0_exe895_1,
		output 		lvb_c0_exe996_1,
		output [63:0] 		lvb_c0_exe1097_1,
		output 		lvb_c0_exe1198_1,
		output 		lvb_c0_exe1299_1,
		output [31:0] 		lvb_c1_exe1_1,
		output [31:0] 		lvb_c1_exe2_1,
		input [31:0] 		workgroup_size,
		input 		start
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [447:0] input_c0_exit87_c0_exi1386_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe794_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe895_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe996_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_c0_exe1097_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe1198_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe1299_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c1_exe1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c1_exe2_staging_reg_NO_SHIFT_REG;
 reg [447:0] local_lvm_c0_exit87_c0_exi1386_NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe794_NO_SHIFT_REG;
 reg local_lvm_c0_exe895_NO_SHIFT_REG;
 reg local_lvm_c0_exe996_NO_SHIFT_REG;
 reg [63:0] local_lvm_c0_exe1097_NO_SHIFT_REG;
 reg local_lvm_c0_exe1198_NO_SHIFT_REG;
 reg local_lvm_c0_exe1299_NO_SHIFT_REG;
 reg [31:0] local_lvm_c1_exe1_NO_SHIFT_REG;
 reg [31:0] local_lvm_c1_exe2_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_c0_exit87_c0_exi1386_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe794_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe895_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe996_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1097_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1198_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1299_staging_reg_NO_SHIFT_REG <= 'x;
		input_c1_exe1_staging_reg_NO_SHIFT_REG <= 'x;
		input_c1_exe2_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_c0_exit87_c0_exi1386_staging_reg_NO_SHIFT_REG <= input_c0_exit87_c0_exi1386;
				input_c0_exe794_staging_reg_NO_SHIFT_REG <= input_c0_exe794;
				input_c0_exe895_staging_reg_NO_SHIFT_REG <= input_c0_exe895;
				input_c0_exe996_staging_reg_NO_SHIFT_REG <= input_c0_exe996;
				input_c0_exe1097_staging_reg_NO_SHIFT_REG <= input_c0_exe1097;
				input_c0_exe1198_staging_reg_NO_SHIFT_REG <= input_c0_exe1198;
				input_c0_exe1299_staging_reg_NO_SHIFT_REG <= input_c0_exe1299;
				input_c1_exe1_staging_reg_NO_SHIFT_REG <= input_c1_exe1;
				input_c1_exe2_staging_reg_NO_SHIFT_REG <= input_c1_exe2;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_c0_exit87_c0_exi1386_NO_SHIFT_REG <= input_c0_exit87_c0_exi1386_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe794_NO_SHIFT_REG <= input_c0_exe794_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe895_NO_SHIFT_REG <= input_c0_exe895_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe996_NO_SHIFT_REG <= input_c0_exe996_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1097_NO_SHIFT_REG <= input_c0_exe1097_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1198_NO_SHIFT_REG <= input_c0_exe1198_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1299_NO_SHIFT_REG <= input_c0_exe1299_staging_reg_NO_SHIFT_REG;
					local_lvm_c1_exe1_NO_SHIFT_REG <= input_c1_exe1_staging_reg_NO_SHIFT_REG;
					local_lvm_c1_exe2_NO_SHIFT_REG <= input_c1_exe2_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_c0_exit87_c0_exi1386_NO_SHIFT_REG <= input_c0_exit87_c0_exi1386;
					local_lvm_c0_exe794_NO_SHIFT_REG <= input_c0_exe794;
					local_lvm_c0_exe895_NO_SHIFT_REG <= input_c0_exe895;
					local_lvm_c0_exe996_NO_SHIFT_REG <= input_c0_exe996;
					local_lvm_c0_exe1097_NO_SHIFT_REG <= input_c0_exe1097;
					local_lvm_c0_exe1198_NO_SHIFT_REG <= input_c0_exe1198;
					local_lvm_c0_exe1299_NO_SHIFT_REG <= input_c0_exe1299;
					local_lvm_c1_exe1_NO_SHIFT_REG <= input_c1_exe1;
					local_lvm_c1_exe2_NO_SHIFT_REG <= input_c1_exe2;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5_c0_exe13100_valid_out;
wire local_bb5_c0_exe13100_stall_in;
wire local_bb5_c0_exe13100_inputs_ready;
wire local_bb5_c0_exe13100_stall_local;
wire local_bb5_c0_exe13100;

assign local_bb5_c0_exe13100_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb5_c0_exe13100 = local_lvm_c0_exit87_c0_exi1386_NO_SHIFT_REG[400];
assign local_bb5_c0_exe13100_valid_out = local_bb5_c0_exe13100_inputs_ready;
assign local_bb5_c0_exe13100_stall_local = local_bb5_c0_exe13100_stall_in;
assign merge_node_stall_in_0 = (|local_bb5_c0_exe13100_stall_local);

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [31:0] lvb_c0_exe794_0_reg_NO_SHIFT_REG;
 reg lvb_c0_exe895_0_reg_NO_SHIFT_REG;
 reg lvb_c0_exe996_0_reg_NO_SHIFT_REG;
 reg [63:0] lvb_c0_exe1097_0_reg_NO_SHIFT_REG;
 reg lvb_c0_exe1198_0_reg_NO_SHIFT_REG;
 reg lvb_c0_exe1299_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_c1_exe1_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_c1_exe2_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb5_c0_exe13100_valid_out & merge_node_valid_out_1_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb5_c0_exe13100_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign merge_node_stall_in_1 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_c0_exe794_0 = lvb_c0_exe794_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe794_1 = lvb_c0_exe794_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe895_0 = lvb_c0_exe895_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe895_1 = lvb_c0_exe895_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe996_0 = lvb_c0_exe996_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe996_1 = lvb_c0_exe996_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1097_0 = lvb_c0_exe1097_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1097_1 = lvb_c0_exe1097_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1198_0 = lvb_c0_exe1198_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1198_1 = lvb_c0_exe1198_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1299_0 = lvb_c0_exe1299_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe1299_1 = lvb_c0_exe1299_0_reg_NO_SHIFT_REG;
assign lvb_c1_exe1_0 = lvb_c1_exe1_0_reg_NO_SHIFT_REG;
assign lvb_c1_exe1_1 = lvb_c1_exe1_0_reg_NO_SHIFT_REG;
assign lvb_c1_exe2_0 = lvb_c1_exe2_0_reg_NO_SHIFT_REG;
assign lvb_c1_exe2_1 = lvb_c1_exe2_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_c0_exe794_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe895_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe996_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe1097_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe1198_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe1299_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c1_exe1_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c1_exe2_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_c0_exe794_0_reg_NO_SHIFT_REG <= local_lvm_c0_exe794_NO_SHIFT_REG;
			lvb_c0_exe895_0_reg_NO_SHIFT_REG <= local_lvm_c0_exe895_NO_SHIFT_REG;
			lvb_c0_exe996_0_reg_NO_SHIFT_REG <= local_lvm_c0_exe996_NO_SHIFT_REG;
			lvb_c0_exe1097_0_reg_NO_SHIFT_REG <= local_lvm_c0_exe1097_NO_SHIFT_REG;
			lvb_c0_exe1198_0_reg_NO_SHIFT_REG <= local_lvm_c0_exe1198_NO_SHIFT_REG;
			lvb_c0_exe1299_0_reg_NO_SHIFT_REG <= local_lvm_c0_exe1299_NO_SHIFT_REG;
			lvb_c1_exe1_0_reg_NO_SHIFT_REG <= local_lvm_c1_exe1_NO_SHIFT_REG;
			lvb_c1_exe2_0_reg_NO_SHIFT_REG <= local_lvm_c1_exe2_NO_SHIFT_REG;
			branch_compare_result_NO_SHIFT_REG <= local_bb5_c0_exe13100;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_6
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_out,
		input [31:0] 		input_wii_div,
		input [31:0] 		input_wii_div1,
		input 		input_wii_cmp19,
		input [31:0] 		input_wii_add7,
		input [31:0] 		input_wii_sub20,
		input [31:0] 		input_wii_sub22,
		input 		input_wii_var_,
		input 		input_wii_var__u61,
		input 		input_wii_var__u62,
		input 		input_wii_var__u63,
		input 		valid_in,
		output 		stall_out,
		input [31:0] 		input_c0_exe794,
		input 		input_c0_exe895,
		input 		input_c0_exe996,
		input [63:0] 		input_c0_exe1097,
		input 		input_c0_exe1198,
		input 		input_c0_exe1299,
		input [31:0] 		input_c1_exe1,
		input [31:0] 		input_c1_exe2,
		output 		valid_out_0,
		input 		stall_in_0,
		output 		lvb_c0_exe895_0,
		output 		lvb_c0_exe996_0,
		output 		lvb_bb6_st_c0_exe1108_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output 		lvb_c0_exe895_1,
		output 		lvb_c0_exe996_1,
		output 		lvb_bb6_st_c0_exe1108_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input [511:0] 		avm_local_bb6_st_c0_exe1108_readdata,
		input 		avm_local_bb6_st_c0_exe1108_readdatavalid,
		input 		avm_local_bb6_st_c0_exe1108_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe1108_address,
		output 		avm_local_bb6_st_c0_exe1108_read,
		output 		avm_local_bb6_st_c0_exe1108_write,
		input 		avm_local_bb6_st_c0_exe1108_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe1108_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe1108_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe1108_burstcount,
		output 		local_bb6_st_c0_exe1108_active,
		input 		clock2x,
		output 		feedback_valid_out_11,
		input 		feedback_stall_in_11,
		output 		feedback_data_out_11
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe794_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe895_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe996_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_c0_exe1097_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe1198_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe1299_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c1_exe1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c1_exe2_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe794_NO_SHIFT_REG;
 reg local_lvm_c0_exe895_NO_SHIFT_REG;
 reg local_lvm_c0_exe996_NO_SHIFT_REG;
 reg [63:0] local_lvm_c0_exe1097_NO_SHIFT_REG;
 reg local_lvm_c0_exe1198_NO_SHIFT_REG;
 reg local_lvm_c0_exe1299_NO_SHIFT_REG;
 reg [31:0] local_lvm_c1_exe1_NO_SHIFT_REG;
 reg [31:0] local_lvm_c1_exe2_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_c0_exe794_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe895_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe996_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1097_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1198_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe1299_staging_reg_NO_SHIFT_REG <= 'x;
		input_c1_exe1_staging_reg_NO_SHIFT_REG <= 'x;
		input_c1_exe2_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_c0_exe794_staging_reg_NO_SHIFT_REG <= input_c0_exe794;
				input_c0_exe895_staging_reg_NO_SHIFT_REG <= input_c0_exe895;
				input_c0_exe996_staging_reg_NO_SHIFT_REG <= input_c0_exe996;
				input_c0_exe1097_staging_reg_NO_SHIFT_REG <= input_c0_exe1097;
				input_c0_exe1198_staging_reg_NO_SHIFT_REG <= input_c0_exe1198;
				input_c0_exe1299_staging_reg_NO_SHIFT_REG <= input_c0_exe1299;
				input_c1_exe1_staging_reg_NO_SHIFT_REG <= input_c1_exe1;
				input_c1_exe2_staging_reg_NO_SHIFT_REG <= input_c1_exe2;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_c0_exe794_NO_SHIFT_REG <= input_c0_exe794_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe895_NO_SHIFT_REG <= input_c0_exe895_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe996_NO_SHIFT_REG <= input_c0_exe996_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1097_NO_SHIFT_REG <= input_c0_exe1097_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1198_NO_SHIFT_REG <= input_c0_exe1198_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe1299_NO_SHIFT_REG <= input_c0_exe1299_staging_reg_NO_SHIFT_REG;
					local_lvm_c1_exe1_NO_SHIFT_REG <= input_c1_exe1_staging_reg_NO_SHIFT_REG;
					local_lvm_c1_exe2_NO_SHIFT_REG <= input_c1_exe2_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_c0_exe794_NO_SHIFT_REG <= input_c0_exe794;
					local_lvm_c0_exe895_NO_SHIFT_REG <= input_c0_exe895;
					local_lvm_c0_exe996_NO_SHIFT_REG <= input_c0_exe996;
					local_lvm_c0_exe1097_NO_SHIFT_REG <= input_c0_exe1097;
					local_lvm_c0_exe1198_NO_SHIFT_REG <= input_c0_exe1198;
					local_lvm_c0_exe1299_NO_SHIFT_REG <= input_c0_exe1299;
					local_lvm_c1_exe1_NO_SHIFT_REG <= input_c1_exe1;
					local_lvm_c1_exe2_NO_SHIFT_REG <= input_c1_exe2;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_c0_eni1101_stall_local;
wire [95:0] local_bb6_c0_eni1101;

assign local_bb6_c0_eni1101[31:0] = 32'bx;
assign local_bb6_c0_eni1101[63:32] = local_lvm_c1_exe1_NO_SHIFT_REG;
assign local_bb6_c0_eni1101[95:64] = 32'bx;

// This section implements an unregistered operation.
// 
wire local_bb6_var__stall_local;
wire [31:0] local_bb6_var_;

assign local_bb6_var_ = local_lvm_c0_exe1097_NO_SHIFT_REG[31:0];

// Register node:
//  * latency = 19
//  * capacity = 19
 logic rnode_1to20_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_1to20_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_1to20_var__0_reg_20_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to20_var__0_valid_out_reg_20_NO_SHIFT_REG;
 logic rnode_1to20_var__0_stall_in_reg_20_NO_SHIFT_REG;
 logic rnode_1to20_var__0_stall_out_reg_20_NO_SHIFT_REG;

acl_data_fifo rnode_1to20_var__0_reg_20_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to20_var__0_reg_20_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to20_var__0_stall_in_reg_20_NO_SHIFT_REG),
	.valid_out(rnode_1to20_var__0_valid_out_reg_20_NO_SHIFT_REG),
	.stall_out(rnode_1to20_var__0_stall_out_reg_20_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to20_var__0_reg_20_fifo.DEPTH = 20;
defparam rnode_1to20_var__0_reg_20_fifo.DATA_WIDTH = 0;
defparam rnode_1to20_var__0_reg_20_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to20_var__0_reg_20_fifo.IMPL = "ram";

assign rnode_1to20_var__0_reg_20_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_4_NO_SHIFT_REG;
assign merge_node_stall_in_4 = rnode_1to20_var__0_stall_out_reg_20_NO_SHIFT_REG;
assign rnode_1to20_var__0_stall_in_reg_20_NO_SHIFT_REG = rnode_1to20_var__0_stall_in_NO_SHIFT_REG;
assign rnode_1to20_var__0_valid_out_NO_SHIFT_REG = rnode_1to20_var__0_valid_out_reg_20_NO_SHIFT_REG;

// Register node:
//  * latency = 179
//  * capacity = 179
 logic rnode_1to180_c0_exe1299_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to180_c0_exe1299_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to180_c0_exe1299_0_NO_SHIFT_REG;
 logic rnode_1to180_c0_exe1299_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to180_c0_exe1299_0_reg_180_NO_SHIFT_REG;
 logic rnode_1to180_c0_exe1299_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_1to180_c0_exe1299_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_1to180_c0_exe1299_0_stall_out_reg_180_NO_SHIFT_REG;
wire [2:0] rci_rcnode_1to181_rc6_c0_exe895_0_reg_1;

acl_data_fifo rnode_1to180_c0_exe1299_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to180_c0_exe1299_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to180_c0_exe1299_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_1to180_c0_exe1299_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_1to180_c0_exe1299_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_lvm_c0_exe1299_NO_SHIFT_REG),
	.data_out(rnode_1to180_c0_exe1299_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_1to180_c0_exe1299_0_reg_180_fifo.DEPTH = 180;
defparam rnode_1to180_c0_exe1299_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_1to180_c0_exe1299_0_reg_180_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to180_c0_exe1299_0_reg_180_fifo.IMPL = "ram";

assign rnode_1to180_c0_exe1299_0_reg_180_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign merge_node_stall_in_5 = rnode_1to180_c0_exe1299_0_stall_out_reg_180_NO_SHIFT_REG;
assign rnode_1to180_c0_exe1299_0_NO_SHIFT_REG = rnode_1to180_c0_exe1299_0_reg_180_NO_SHIFT_REG;
assign rnode_1to180_c0_exe1299_0_stall_in_reg_180_NO_SHIFT_REG = rnode_1to180_c0_exe1299_0_stall_in_NO_SHIFT_REG;
assign rnode_1to180_c0_exe1299_0_valid_out_NO_SHIFT_REG = rnode_1to180_c0_exe1299_0_valid_out_reg_180_NO_SHIFT_REG;
assign rci_rcnode_1to181_rc6_c0_exe895_0_reg_1[0] = local_lvm_c0_exe895_NO_SHIFT_REG;
assign rci_rcnode_1to181_rc6_c0_exe895_0_reg_1[1] = local_lvm_c0_exe996_NO_SHIFT_REG;
assign rci_rcnode_1to181_rc6_c0_exe895_0_reg_1[2] = local_lvm_c0_exe1198_NO_SHIFT_REG;

// Register node:
//  * latency = 180
//  * capacity = 180
 logic rcnode_1to181_rc6_c0_exe895_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to181_rc6_c0_exe895_0_stall_in_NO_SHIFT_REG;
 logic [2:0] rcnode_1to181_rc6_c0_exe895_0_NO_SHIFT_REG;
 logic rcnode_1to181_rc6_c0_exe895_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [2:0] rcnode_1to181_rc6_c0_exe895_0_reg_181_NO_SHIFT_REG;
 logic rcnode_1to181_rc6_c0_exe895_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rcnode_1to181_rc6_c0_exe895_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rcnode_1to181_rc6_c0_exe895_0_stall_out_reg_181_IP_NO_SHIFT_REG;
 logic rcnode_1to181_rc6_c0_exe895_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rcnode_1to181_rc6_c0_exe895_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to181_rc6_c0_exe895_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to181_rc6_c0_exe895_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rcnode_1to181_rc6_c0_exe895_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rcnode_1to181_rc6_c0_exe895_0_stall_out_reg_181_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to181_rc6_c0_exe895_0_reg_1),
	.data_out(rcnode_1to181_rc6_c0_exe895_0_reg_181_NO_SHIFT_REG)
);

defparam rcnode_1to181_rc6_c0_exe895_0_reg_181_fifo.DEPTH = 181;
defparam rcnode_1to181_rc6_c0_exe895_0_reg_181_fifo.DATA_WIDTH = 3;
defparam rcnode_1to181_rc6_c0_exe895_0_reg_181_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to181_rc6_c0_exe895_0_reg_181_fifo.IMPL = "ram";

assign rcnode_1to181_rc6_c0_exe895_0_reg_181_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_6_NO_SHIFT_REG;
assign rcnode_1to181_rc6_c0_exe895_0_stall_out_reg_181_NO_SHIFT_REG = (~(rcnode_1to181_rc6_c0_exe895_0_reg_181_inputs_ready_NO_SHIFT_REG) | rcnode_1to181_rc6_c0_exe895_0_stall_out_reg_181_IP_NO_SHIFT_REG);
assign merge_node_stall_in_6 = rcnode_1to181_rc6_c0_exe895_0_stall_out_reg_181_NO_SHIFT_REG;
assign rcnode_1to181_rc6_c0_exe895_0_NO_SHIFT_REG = rcnode_1to181_rc6_c0_exe895_0_reg_181_NO_SHIFT_REG;
assign rcnode_1to181_rc6_c0_exe895_0_stall_in_reg_181_NO_SHIFT_REG = rcnode_1to181_rc6_c0_exe895_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to181_rc6_c0_exe895_0_valid_out_NO_SHIFT_REG = rcnode_1to181_rc6_c0_exe895_0_valid_out_reg_181_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb6_c0_eni2102_valid_out;
wire local_bb6_c0_eni2102_stall_in;
wire local_bb6_c0_eni2102_inputs_ready;
wire local_bb6_c0_eni2102_stall_local;
wire [95:0] local_bb6_c0_eni2102;

assign local_bb6_c0_eni2102_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign local_bb6_c0_eni2102[63:0] = local_bb6_c0_eni1101[63:0];
assign local_bb6_c0_eni2102[95:64] = local_lvm_c1_exe2_NO_SHIFT_REG;
assign local_bb6_c0_eni2102_valid_out = local_bb6_c0_eni2102_inputs_ready;
assign local_bb6_c0_eni2102_stall_local = local_bb6_c0_eni2102_stall_in;
assign merge_node_stall_in_0 = (local_bb6_c0_eni2102_stall_local | ~(local_bb6_c0_eni2102_inputs_ready));
assign merge_node_stall_in_1 = (local_bb6_c0_eni2102_stall_local | ~(local_bb6_c0_eni2102_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb6_add38_valid_out;
wire local_bb6_add38_stall_in;
wire local_bb6_add38_inputs_ready;
wire local_bb6_add38_stall_local;
wire [31:0] local_bb6_add38;

assign local_bb6_add38_inputs_ready = (merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_3_NO_SHIFT_REG);
assign local_bb6_add38 = (local_bb6_var_ + local_lvm_c0_exe794_NO_SHIFT_REG);
assign local_bb6_add38_valid_out = local_bb6_add38_inputs_ready;
assign local_bb6_add38_stall_local = local_bb6_add38_stall_in;
assign merge_node_stall_in_2 = (local_bb6_add38_stall_local | ~(local_bb6_add38_inputs_ready));
assign merge_node_stall_in_3 = (local_bb6_add38_stall_local | ~(local_bb6_add38_inputs_ready));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_20to21_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_20to21_var__0_stall_in_NO_SHIFT_REG;
 logic rnode_20to21_var__0_reg_21_inputs_ready_NO_SHIFT_REG;
 logic rnode_20to21_var__0_valid_out_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_var__0_stall_in_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_var__0_stall_out_reg_21_NO_SHIFT_REG;

acl_data_fifo rnode_20to21_var__0_reg_21_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_20to21_var__0_reg_21_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_20to21_var__0_stall_in_reg_21_NO_SHIFT_REG),
	.valid_out(rnode_20to21_var__0_valid_out_reg_21_NO_SHIFT_REG),
	.stall_out(rnode_20to21_var__0_stall_out_reg_21_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_20to21_var__0_reg_21_fifo.DEPTH = 2;
defparam rnode_20to21_var__0_reg_21_fifo.DATA_WIDTH = 0;
defparam rnode_20to21_var__0_reg_21_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_20to21_var__0_reg_21_fifo.IMPL = "ll_reg";

assign rnode_20to21_var__0_reg_21_inputs_ready_NO_SHIFT_REG = rnode_1to20_var__0_valid_out_NO_SHIFT_REG;
assign rnode_1to20_var__0_stall_in_NO_SHIFT_REG = rnode_20to21_var__0_stall_out_reg_21_NO_SHIFT_REG;
assign rnode_20to21_var__0_stall_in_reg_21_NO_SHIFT_REG = rnode_20to21_var__0_stall_in_NO_SHIFT_REG;
assign rnode_20to21_var__0_valid_out_NO_SHIFT_REG = rnode_20to21_var__0_valid_out_reg_21_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_c0_exe1299_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_c0_exe1299_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_c0_exe1299_0_NO_SHIFT_REG;
 logic rnode_180to181_c0_exe1299_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_c0_exe1299_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_c0_exe1299_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_c0_exe1299_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_c0_exe1299_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_c0_exe1299_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_c0_exe1299_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_c0_exe1299_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_c0_exe1299_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_c0_exe1299_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(rnode_1to180_c0_exe1299_0_NO_SHIFT_REG),
	.data_out(rnode_180to181_c0_exe1299_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_c0_exe1299_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_c0_exe1299_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_c0_exe1299_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_c0_exe1299_0_reg_181_fifo.IMPL = "ll_reg";

assign rnode_180to181_c0_exe1299_0_reg_181_inputs_ready_NO_SHIFT_REG = rnode_1to180_c0_exe1299_0_valid_out_NO_SHIFT_REG;
assign rnode_1to180_c0_exe1299_0_stall_in_NO_SHIFT_REG = rnode_180to181_c0_exe1299_0_stall_out_reg_181_NO_SHIFT_REG;
assign rnode_180to181_c0_exe1299_0_NO_SHIFT_REG = rnode_180to181_c0_exe1299_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_c0_exe1299_0_stall_in_reg_181_NO_SHIFT_REG = rnode_180to181_c0_exe1299_0_stall_in_NO_SHIFT_REG;
assign rnode_180to181_c0_exe1299_0_valid_out_NO_SHIFT_REG = rnode_180to181_c0_exe1299_0_valid_out_reg_181_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb6_c0_enter103_c0_eni2102_inputs_ready;
 reg local_bb6_c0_enter103_c0_eni2102_valid_out_0_NO_SHIFT_REG;
wire local_bb6_c0_enter103_c0_eni2102_stall_in_0;
 reg local_bb6_c0_enter103_c0_eni2102_valid_out_1_NO_SHIFT_REG;
wire local_bb6_c0_enter103_c0_eni2102_stall_in_1;
 reg local_bb6_c0_enter103_c0_eni2102_valid_out_2_NO_SHIFT_REG;
wire local_bb6_c0_enter103_c0_eni2102_stall_in_2;
wire local_bb6_c0_enter103_c0_eni2102_output_regs_ready;
 reg [95:0] local_bb6_c0_enter103_c0_eni2102_NO_SHIFT_REG;
wire local_bb6_c0_enter103_c0_eni2102_input_accepted;
 reg local_bb6_c0_enter103_c0_eni2102_valid_bit_NO_SHIFT_REG;
wire local_bb6_c0_exit107_c0_exi1106_entry_stall;
wire local_bb6_c0_exit107_c0_exi1106_output_regs_ready;
wire [15:0] local_bb6_c0_exit107_c0_exi1106_valid_bits;
wire local_bb6_c0_exit107_c0_exi1106_valid_in;
wire local_bb6_c0_exit107_c0_exi1106_phases;
wire local_bb6_c0_enter103_c0_eni2102_inc_pipelined_thread;
wire local_bb6_c0_enter103_c0_eni2102_dec_pipelined_thread;
wire local_bb6_c0_enter103_c0_eni2102_causedstall;

assign local_bb6_c0_enter103_c0_eni2102_inputs_ready = local_bb6_c0_eni2102_valid_out;
assign local_bb6_c0_enter103_c0_eni2102_output_regs_ready = 1'b1;
assign local_bb6_c0_enter103_c0_eni2102_input_accepted = (local_bb6_c0_enter103_c0_eni2102_inputs_ready && !(local_bb6_c0_exit107_c0_exi1106_entry_stall));
assign local_bb6_c0_enter103_c0_eni2102_inc_pipelined_thread = 1'b1;
assign local_bb6_c0_enter103_c0_eni2102_dec_pipelined_thread = ~(1'b0);
assign local_bb6_c0_eni2102_stall_in = ((~(local_bb6_c0_enter103_c0_eni2102_inputs_ready) | local_bb6_c0_exit107_c0_exi1106_entry_stall) | ~(1'b1));
assign local_bb6_c0_enter103_c0_eni2102_causedstall = (1'b1 && ((~(local_bb6_c0_enter103_c0_eni2102_inputs_ready) | local_bb6_c0_exit107_c0_exi1106_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_enter103_c0_eni2102_valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb6_c0_enter103_c0_eni2102_valid_bit_NO_SHIFT_REG <= local_bb6_c0_enter103_c0_eni2102_input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_enter103_c0_eni2102_NO_SHIFT_REG <= 'x;
		local_bb6_c0_enter103_c0_eni2102_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter103_c0_eni2102_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter103_c0_eni2102_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_c0_enter103_c0_eni2102_output_regs_ready)
		begin
			local_bb6_c0_enter103_c0_eni2102_NO_SHIFT_REG <= local_bb6_c0_eni2102;
			local_bb6_c0_enter103_c0_eni2102_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter103_c0_eni2102_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter103_c0_eni2102_valid_out_2_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb6_c0_enter103_c0_eni2102_stall_in_0))
			begin
				local_bb6_c0_enter103_c0_eni2102_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter103_c0_eni2102_stall_in_1))
			begin
				local_bb6_c0_enter103_c0_eni2102_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter103_c0_eni2102_stall_in_2))
			begin
				local_bb6_c0_enter103_c0_eni2102_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 18
//  * capacity = 18
 logic rnode_1to19_bb6_add38_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to19_bb6_add38_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to19_bb6_add38_0_NO_SHIFT_REG;
 logic rnode_1to19_bb6_add38_0_reg_19_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to19_bb6_add38_0_reg_19_NO_SHIFT_REG;
 logic rnode_1to19_bb6_add38_0_valid_out_reg_19_NO_SHIFT_REG;
 logic rnode_1to19_bb6_add38_0_stall_in_reg_19_NO_SHIFT_REG;
 logic rnode_1to19_bb6_add38_0_stall_out_reg_19_NO_SHIFT_REG;

acl_data_fifo rnode_1to19_bb6_add38_0_reg_19_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to19_bb6_add38_0_reg_19_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to19_bb6_add38_0_stall_in_reg_19_NO_SHIFT_REG),
	.valid_out(rnode_1to19_bb6_add38_0_valid_out_reg_19_NO_SHIFT_REG),
	.stall_out(rnode_1to19_bb6_add38_0_stall_out_reg_19_NO_SHIFT_REG),
	.data_in(local_bb6_add38),
	.data_out(rnode_1to19_bb6_add38_0_reg_19_NO_SHIFT_REG)
);

defparam rnode_1to19_bb6_add38_0_reg_19_fifo.DEPTH = 19;
defparam rnode_1to19_bb6_add38_0_reg_19_fifo.DATA_WIDTH = 32;
defparam rnode_1to19_bb6_add38_0_reg_19_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to19_bb6_add38_0_reg_19_fifo.IMPL = "ram";

assign rnode_1to19_bb6_add38_0_reg_19_inputs_ready_NO_SHIFT_REG = local_bb6_add38_valid_out;
assign local_bb6_add38_stall_in = rnode_1to19_bb6_add38_0_stall_out_reg_19_NO_SHIFT_REG;
assign rnode_1to19_bb6_add38_0_NO_SHIFT_REG = rnode_1to19_bb6_add38_0_reg_19_NO_SHIFT_REG;
assign rnode_1to19_bb6_add38_0_stall_in_reg_19_NO_SHIFT_REG = rnode_1to19_bb6_add38_0_stall_in_NO_SHIFT_REG;
assign rnode_1to19_bb6_add38_0_valid_out_NO_SHIFT_REG = rnode_1to19_bb6_add38_0_valid_out_reg_19_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb6_c0_ene1104_valid_out;
wire local_bb6_c0_ene1104_stall_in;
wire local_bb6_c0_ene1104_inputs_ready;
wire local_bb6_c0_ene1104_stall_local;
wire [31:0] local_bb6_c0_ene1104;

assign local_bb6_c0_ene1104_inputs_ready = local_bb6_c0_enter103_c0_eni2102_valid_out_0_NO_SHIFT_REG;
assign local_bb6_c0_ene1104 = local_bb6_c0_enter103_c0_eni2102_NO_SHIFT_REG[63:32];
assign local_bb6_c0_ene1104_valid_out = 1'b1;
assign local_bb6_c0_enter103_c0_eni2102_stall_in_0 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb6_c0_ene2105_valid_out;
wire local_bb6_c0_ene2105_stall_in;
wire local_bb6_c0_ene2105_inputs_ready;
wire local_bb6_c0_ene2105_stall_local;
wire [31:0] local_bb6_c0_ene2105;

assign local_bb6_c0_ene2105_inputs_ready = local_bb6_c0_enter103_c0_eni2102_valid_out_1_NO_SHIFT_REG;
assign local_bb6_c0_ene2105 = local_bb6_c0_enter103_c0_eni2102_NO_SHIFT_REG[95:64];
assign local_bb6_c0_ene2105_valid_out = 1'b1;
assign local_bb6_c0_enter103_c0_eni2102_stall_in_1 = 1'b0;

// This section implements an unregistered operation.
// 
wire SFC_4_VALID_2_2_0_valid_out;
wire SFC_4_VALID_2_2_0_stall_in;
wire SFC_4_VALID_2_2_0_inputs_ready;
wire SFC_4_VALID_2_2_0_stall_local;
wire SFC_4_VALID_2_2_0;

assign SFC_4_VALID_2_2_0_inputs_ready = local_bb6_c0_enter103_c0_eni2102_valid_out_2_NO_SHIFT_REG;
assign SFC_4_VALID_2_2_0 = local_bb6_c0_enter103_c0_eni2102_valid_bit_NO_SHIFT_REG;
assign SFC_4_VALID_2_2_0_valid_out = 1'b1;
assign local_bb6_c0_enter103_c0_eni2102_stall_in_2 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_19to20_bb6_add38_0_valid_out_NO_SHIFT_REG;
 logic rnode_19to20_bb6_add38_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_19to20_bb6_add38_0_NO_SHIFT_REG;
 logic rnode_19to20_bb6_add38_0_reg_20_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_19to20_bb6_add38_0_reg_20_NO_SHIFT_REG;
 logic rnode_19to20_bb6_add38_0_valid_out_reg_20_NO_SHIFT_REG;
 logic rnode_19to20_bb6_add38_0_stall_in_reg_20_NO_SHIFT_REG;
 logic rnode_19to20_bb6_add38_0_stall_out_reg_20_NO_SHIFT_REG;

acl_data_fifo rnode_19to20_bb6_add38_0_reg_20_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_19to20_bb6_add38_0_reg_20_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_19to20_bb6_add38_0_stall_in_reg_20_NO_SHIFT_REG),
	.valid_out(rnode_19to20_bb6_add38_0_valid_out_reg_20_NO_SHIFT_REG),
	.stall_out(rnode_19to20_bb6_add38_0_stall_out_reg_20_NO_SHIFT_REG),
	.data_in(rnode_1to19_bb6_add38_0_NO_SHIFT_REG),
	.data_out(rnode_19to20_bb6_add38_0_reg_20_NO_SHIFT_REG)
);

defparam rnode_19to20_bb6_add38_0_reg_20_fifo.DEPTH = 1;
defparam rnode_19to20_bb6_add38_0_reg_20_fifo.DATA_WIDTH = 32;
defparam rnode_19to20_bb6_add38_0_reg_20_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_19to20_bb6_add38_0_reg_20_fifo.IMPL = "ll_reg";

assign rnode_19to20_bb6_add38_0_reg_20_inputs_ready_NO_SHIFT_REG = rnode_1to19_bb6_add38_0_valid_out_NO_SHIFT_REG;
assign rnode_1to19_bb6_add38_0_stall_in_NO_SHIFT_REG = rnode_19to20_bb6_add38_0_stall_out_reg_20_NO_SHIFT_REG;
assign rnode_19to20_bb6_add38_0_NO_SHIFT_REG = rnode_19to20_bb6_add38_0_reg_20_NO_SHIFT_REG;
assign rnode_19to20_bb6_add38_0_stall_in_reg_20_NO_SHIFT_REG = rnode_19to20_bb6_add38_0_stall_in_NO_SHIFT_REG;
assign rnode_19to20_bb6_add38_0_valid_out_NO_SHIFT_REG = rnode_19to20_bb6_add38_0_valid_out_reg_20_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb6_div36_inputs_ready;
 reg local_bb6_div36_valid_out_NO_SHIFT_REG;
wire local_bb6_div36_stall_in;
wire local_bb6_div36_output_regs_ready;
wire [31:0] local_bb6_div36;
 reg local_bb6_div36_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb6_div36_valid_pipe_12_NO_SHIFT_REG;
wire local_bb6_div36_causedstall;

acl_fp_div_s5 fp_module_local_bb6_div36 (
	.clock(clock),
	.dataa(local_bb6_c0_ene1104),
	.datab(local_bb6_c0_ene2105),
	.enable(local_bb6_div36_output_regs_ready),
	.result(local_bb6_div36)
);


assign local_bb6_div36_inputs_ready = 1'b1;
assign local_bb6_div36_output_regs_ready = 1'b1;
assign local_bb6_c0_ene1104_stall_in = 1'b0;
assign local_bb6_c0_ene2105_stall_in = 1'b0;
assign local_bb6_div36_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_div36_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb6_div36_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_div36_output_regs_ready)
		begin
			local_bb6_div36_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb6_div36_valid_pipe_1_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_0_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_2_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_1_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_3_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_2_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_4_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_3_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_5_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_4_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_6_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_5_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_7_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_6_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_8_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_7_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_9_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_8_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_10_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_9_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_11_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_10_NO_SHIFT_REG;
			local_bb6_div36_valid_pipe_12_NO_SHIFT_REG <= local_bb6_div36_valid_pipe_11_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_div36_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_div36_output_regs_ready)
		begin
			local_bb6_div36_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb6_div36_stall_in))
			begin
				local_bb6_div36_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_2_3_0_inputs_ready;
 reg SFC_4_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_2_3_0_stall_in;
wire SFC_4_VALID_2_3_0_output_regs_ready;
 reg SFC_4_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_2_3_0_causedstall;

assign SFC_4_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_4_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_2_2_0_stall_in = 1'b0;
assign SFC_4_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_2_3_0_output_regs_ready)
		begin
			SFC_4_VALID_2_3_0_NO_SHIFT_REG <= SFC_4_VALID_2_2_0;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_idxprom39_stall_local;
wire [63:0] local_bb6_idxprom39;

assign local_bb6_idxprom39[63:32] = 32'h0;
assign local_bb6_idxprom39[31:0] = rnode_19to20_bb6_add38_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exi1106_valid_out;
wire local_bb6_c0_exi1106_stall_in;
wire local_bb6_c0_exi1106_inputs_ready;
wire local_bb6_c0_exi1106_stall_local;
wire [63:0] local_bb6_c0_exi1106;

assign local_bb6_c0_exi1106_inputs_ready = local_bb6_div36_valid_out_NO_SHIFT_REG;
assign local_bb6_c0_exi1106[31:0] = 32'bx;
assign local_bb6_c0_exi1106[63:32] = local_bb6_div36;
assign local_bb6_c0_exi1106_valid_out = 1'b1;
assign local_bb6_div36_stall_in = 1'b0;

// This section implements a registered operation.
// 
wire SFC_4_VALID_3_4_0_inputs_ready;
 reg SFC_4_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_3_4_0_stall_in;
wire SFC_4_VALID_3_4_0_output_regs_ready;
 reg SFC_4_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_3_4_0_causedstall;

assign SFC_4_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_4_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_2_3_0_stall_in = 1'b0;
assign SFC_4_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_3_4_0_output_regs_ready)
		begin
			SFC_4_VALID_3_4_0_NO_SHIFT_REG <= SFC_4_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_arrayidx40_valid_out;
wire local_bb6_arrayidx40_stall_in;
wire local_bb6_arrayidx40_inputs_ready;
wire local_bb6_arrayidx40_stall_local;
wire [63:0] local_bb6_arrayidx40;

assign local_bb6_arrayidx40_inputs_ready = rnode_19to20_bb6_add38_0_valid_out_NO_SHIFT_REG;
assign local_bb6_arrayidx40 = ((input_out & 64'hFFFFFFFFFFFFFC00) + ((local_bb6_idxprom39 & 64'hFFFFFFFF) << 6'h2));
assign local_bb6_arrayidx40_valid_out = local_bb6_arrayidx40_inputs_ready;
assign local_bb6_arrayidx40_stall_local = local_bb6_arrayidx40_stall_in;
assign rnode_19to20_bb6_add38_0_stall_in_NO_SHIFT_REG = (|local_bb6_arrayidx40_stall_local);

// This section implements a registered operation.
// 
wire SFC_4_VALID_4_5_0_inputs_ready;
 reg SFC_4_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_4_5_0_stall_in;
wire SFC_4_VALID_4_5_0_output_regs_ready;
 reg SFC_4_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_4_5_0_causedstall;

assign SFC_4_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_4_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_3_4_0_stall_in = 1'b0;
assign SFC_4_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_4_5_0_output_regs_ready)
		begin
			SFC_4_VALID_4_5_0_NO_SHIFT_REG <= SFC_4_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_20to21_bb6_arrayidx40_0_valid_out_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx40_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx40_0_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx40_0_reg_21_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx40_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx40_0_valid_out_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx40_0_stall_in_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx40_0_stall_out_reg_21_NO_SHIFT_REG;

acl_data_fifo rnode_20to21_bb6_arrayidx40_0_reg_21_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_20to21_bb6_arrayidx40_0_reg_21_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_20to21_bb6_arrayidx40_0_stall_in_reg_21_NO_SHIFT_REG),
	.valid_out(rnode_20to21_bb6_arrayidx40_0_valid_out_reg_21_NO_SHIFT_REG),
	.stall_out(rnode_20to21_bb6_arrayidx40_0_stall_out_reg_21_NO_SHIFT_REG),
	.data_in((local_bb6_arrayidx40 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_20to21_bb6_arrayidx40_0_reg_21_NO_SHIFT_REG)
);

defparam rnode_20to21_bb6_arrayidx40_0_reg_21_fifo.DEPTH = 2;
defparam rnode_20to21_bb6_arrayidx40_0_reg_21_fifo.DATA_WIDTH = 64;
defparam rnode_20to21_bb6_arrayidx40_0_reg_21_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_20to21_bb6_arrayidx40_0_reg_21_fifo.IMPL = "ll_reg";

assign rnode_20to21_bb6_arrayidx40_0_reg_21_inputs_ready_NO_SHIFT_REG = local_bb6_arrayidx40_valid_out;
assign local_bb6_arrayidx40_stall_in = rnode_20to21_bb6_arrayidx40_0_stall_out_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb6_arrayidx40_0_NO_SHIFT_REG = rnode_20to21_bb6_arrayidx40_0_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb6_arrayidx40_0_stall_in_reg_21_NO_SHIFT_REG = rnode_20to21_bb6_arrayidx40_0_stall_in_NO_SHIFT_REG;
assign rnode_20to21_bb6_arrayidx40_0_valid_out_NO_SHIFT_REG = rnode_20to21_bb6_arrayidx40_0_valid_out_reg_21_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_4_VALID_5_6_0_inputs_ready;
 reg SFC_4_VALID_5_6_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_5_6_0_stall_in;
wire SFC_4_VALID_5_6_0_output_regs_ready;
 reg SFC_4_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_5_6_0_causedstall;

assign SFC_4_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_4_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_4_5_0_stall_in = 1'b0;
assign SFC_4_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_5_6_0_output_regs_ready)
		begin
			SFC_4_VALID_5_6_0_NO_SHIFT_REG <= SFC_4_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_6_7_0_inputs_ready;
 reg SFC_4_VALID_6_7_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_6_7_0_stall_in;
wire SFC_4_VALID_6_7_0_output_regs_ready;
 reg SFC_4_VALID_6_7_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_6_7_0_causedstall;

assign SFC_4_VALID_6_7_0_inputs_ready = 1'b1;
assign SFC_4_VALID_6_7_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_5_6_0_stall_in = 1'b0;
assign SFC_4_VALID_6_7_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_6_7_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_6_7_0_output_regs_ready)
		begin
			SFC_4_VALID_6_7_0_NO_SHIFT_REG <= SFC_4_VALID_5_6_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_7_8_0_inputs_ready;
 reg SFC_4_VALID_7_8_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_7_8_0_stall_in;
wire SFC_4_VALID_7_8_0_output_regs_ready;
 reg SFC_4_VALID_7_8_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_7_8_0_causedstall;

assign SFC_4_VALID_7_8_0_inputs_ready = 1'b1;
assign SFC_4_VALID_7_8_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_6_7_0_stall_in = 1'b0;
assign SFC_4_VALID_7_8_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_7_8_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_7_8_0_output_regs_ready)
		begin
			SFC_4_VALID_7_8_0_NO_SHIFT_REG <= SFC_4_VALID_6_7_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_8_9_0_inputs_ready;
 reg SFC_4_VALID_8_9_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_8_9_0_stall_in;
wire SFC_4_VALID_8_9_0_output_regs_ready;
 reg SFC_4_VALID_8_9_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_8_9_0_causedstall;

assign SFC_4_VALID_8_9_0_inputs_ready = 1'b1;
assign SFC_4_VALID_8_9_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_7_8_0_stall_in = 1'b0;
assign SFC_4_VALID_8_9_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_8_9_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_8_9_0_output_regs_ready)
		begin
			SFC_4_VALID_8_9_0_NO_SHIFT_REG <= SFC_4_VALID_7_8_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_9_10_0_inputs_ready;
 reg SFC_4_VALID_9_10_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_9_10_0_stall_in;
wire SFC_4_VALID_9_10_0_output_regs_ready;
 reg SFC_4_VALID_9_10_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_9_10_0_causedstall;

assign SFC_4_VALID_9_10_0_inputs_ready = 1'b1;
assign SFC_4_VALID_9_10_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_8_9_0_stall_in = 1'b0;
assign SFC_4_VALID_9_10_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_9_10_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_9_10_0_output_regs_ready)
		begin
			SFC_4_VALID_9_10_0_NO_SHIFT_REG <= SFC_4_VALID_8_9_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_10_11_0_inputs_ready;
 reg SFC_4_VALID_10_11_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_10_11_0_stall_in;
wire SFC_4_VALID_10_11_0_output_regs_ready;
 reg SFC_4_VALID_10_11_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_10_11_0_causedstall;

assign SFC_4_VALID_10_11_0_inputs_ready = 1'b1;
assign SFC_4_VALID_10_11_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_9_10_0_stall_in = 1'b0;
assign SFC_4_VALID_10_11_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_10_11_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_10_11_0_output_regs_ready)
		begin
			SFC_4_VALID_10_11_0_NO_SHIFT_REG <= SFC_4_VALID_9_10_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_11_12_0_inputs_ready;
 reg SFC_4_VALID_11_12_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_11_12_0_stall_in;
wire SFC_4_VALID_11_12_0_output_regs_ready;
 reg SFC_4_VALID_11_12_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_11_12_0_causedstall;

assign SFC_4_VALID_11_12_0_inputs_ready = 1'b1;
assign SFC_4_VALID_11_12_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_10_11_0_stall_in = 1'b0;
assign SFC_4_VALID_11_12_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_11_12_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_11_12_0_output_regs_ready)
		begin
			SFC_4_VALID_11_12_0_NO_SHIFT_REG <= SFC_4_VALID_10_11_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_12_13_0_inputs_ready;
 reg SFC_4_VALID_12_13_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_12_13_0_stall_in;
wire SFC_4_VALID_12_13_0_output_regs_ready;
 reg SFC_4_VALID_12_13_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_12_13_0_causedstall;

assign SFC_4_VALID_12_13_0_inputs_ready = 1'b1;
assign SFC_4_VALID_12_13_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_11_12_0_stall_in = 1'b0;
assign SFC_4_VALID_12_13_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_12_13_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_12_13_0_output_regs_ready)
		begin
			SFC_4_VALID_12_13_0_NO_SHIFT_REG <= SFC_4_VALID_11_12_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_13_14_0_inputs_ready;
 reg SFC_4_VALID_13_14_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_13_14_0_stall_in;
wire SFC_4_VALID_13_14_0_output_regs_ready;
 reg SFC_4_VALID_13_14_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_13_14_0_causedstall;

assign SFC_4_VALID_13_14_0_inputs_ready = 1'b1;
assign SFC_4_VALID_13_14_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_12_13_0_stall_in = 1'b0;
assign SFC_4_VALID_13_14_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_13_14_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_13_14_0_output_regs_ready)
		begin
			SFC_4_VALID_13_14_0_NO_SHIFT_REG <= SFC_4_VALID_12_13_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_14_15_0_inputs_ready;
 reg SFC_4_VALID_14_15_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_14_15_0_stall_in;
wire SFC_4_VALID_14_15_0_output_regs_ready;
 reg SFC_4_VALID_14_15_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_14_15_0_causedstall;

assign SFC_4_VALID_14_15_0_inputs_ready = 1'b1;
assign SFC_4_VALID_14_15_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_13_14_0_stall_in = 1'b0;
assign SFC_4_VALID_14_15_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_14_15_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_14_15_0_output_regs_ready)
		begin
			SFC_4_VALID_14_15_0_NO_SHIFT_REG <= SFC_4_VALID_13_14_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_15_16_0_inputs_ready;
 reg SFC_4_VALID_15_16_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_15_16_0_stall_in;
wire SFC_4_VALID_15_16_0_output_regs_ready;
 reg SFC_4_VALID_15_16_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_15_16_0_causedstall;

assign SFC_4_VALID_15_16_0_inputs_ready = 1'b1;
assign SFC_4_VALID_15_16_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_14_15_0_stall_in = 1'b0;
assign SFC_4_VALID_15_16_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_15_16_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_15_16_0_output_regs_ready)
		begin
			SFC_4_VALID_15_16_0_NO_SHIFT_REG <= SFC_4_VALID_14_15_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb6_c0_exit107_c0_exi1106_inputs_ready;
 reg local_bb6_c0_exit107_c0_exi1106_valid_out_NO_SHIFT_REG;
wire local_bb6_c0_exit107_c0_exi1106_stall_in;
 reg [63:0] local_bb6_c0_exit107_c0_exi1106_NO_SHIFT_REG;
wire [63:0] local_bb6_c0_exit107_c0_exi1106_in;
wire local_bb6_c0_exit107_c0_exi1106_valid;
wire local_bb6_c0_exit107_c0_exi1106_causedstall;

acl_stall_free_sink local_bb6_c0_exit107_c0_exi1106_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb6_c0_exi1106),
	.data_out(local_bb6_c0_exit107_c0_exi1106_in),
	.input_accepted(local_bb6_c0_enter103_c0_eni2102_input_accepted),
	.valid_out(local_bb6_c0_exit107_c0_exi1106_valid),
	.stall_in(~(local_bb6_c0_exit107_c0_exi1106_output_regs_ready)),
	.stall_entry(local_bb6_c0_exit107_c0_exi1106_entry_stall),
	.valid_in(local_bb6_c0_exit107_c0_exi1106_valid_in),
	.IIphases(local_bb6_c0_exit107_c0_exi1106_phases),
	.inc_pipelined_thread(local_bb6_c0_enter103_c0_eni2102_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb6_c0_enter103_c0_eni2102_dec_pipelined_thread)
);

defparam local_bb6_c0_exit107_c0_exi1106_instance.DATA_WIDTH = 64;
defparam local_bb6_c0_exit107_c0_exi1106_instance.PIPELINE_DEPTH = 20;
defparam local_bb6_c0_exit107_c0_exi1106_instance.SHARINGII = 1;
defparam local_bb6_c0_exit107_c0_exi1106_instance.SCHEDULEII = 1;
defparam local_bb6_c0_exit107_c0_exi1106_instance.ALWAYS_THROTTLE = 0;

assign local_bb6_c0_exit107_c0_exi1106_inputs_ready = 1'b1;
assign local_bb6_c0_exit107_c0_exi1106_output_regs_ready = (&(~(local_bb6_c0_exit107_c0_exi1106_valid_out_NO_SHIFT_REG) | ~(local_bb6_c0_exit107_c0_exi1106_stall_in)));
assign local_bb6_c0_exit107_c0_exi1106_valid_in = SFC_4_VALID_15_16_0_NO_SHIFT_REG;
assign local_bb6_c0_exi1106_stall_in = 1'b0;
assign SFC_4_VALID_15_16_0_stall_in = 1'b0;
assign local_bb6_c0_exit107_c0_exi1106_causedstall = (1'b1 && (1'b0 && !(~(local_bb6_c0_exit107_c0_exi1106_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_exit107_c0_exi1106_NO_SHIFT_REG <= 'x;
		local_bb6_c0_exit107_c0_exi1106_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_c0_exit107_c0_exi1106_output_regs_ready)
		begin
			local_bb6_c0_exit107_c0_exi1106_NO_SHIFT_REG <= local_bb6_c0_exit107_c0_exi1106_in;
			local_bb6_c0_exit107_c0_exi1106_valid_out_NO_SHIFT_REG <= local_bb6_c0_exit107_c0_exi1106_valid;
		end
		else
		begin
			if (~(local_bb6_c0_exit107_c0_exi1106_stall_in))
			begin
				local_bb6_c0_exit107_c0_exi1106_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_c0_exe1108_valid_out;
wire local_bb6_c0_exe1108_stall_in;
wire local_bb6_c0_exe1108_inputs_ready;
wire local_bb6_c0_exe1108_stall_local;
wire [31:0] local_bb6_c0_exe1108;

assign local_bb6_c0_exe1108_inputs_ready = local_bb6_c0_exit107_c0_exi1106_valid_out_NO_SHIFT_REG;
assign local_bb6_c0_exe1108 = local_bb6_c0_exit107_c0_exi1106_NO_SHIFT_REG[63:32];
assign local_bb6_c0_exe1108_valid_out = local_bb6_c0_exe1108_inputs_ready;
assign local_bb6_c0_exe1108_stall_local = local_bb6_c0_exe1108_stall_in;
assign local_bb6_c0_exit107_c0_exi1106_stall_in = (|local_bb6_c0_exe1108_stall_local);

// This section implements a registered operation.
// 
wire local_bb6_st_c0_exe1108_inputs_ready;
 reg local_bb6_st_c0_exe1108_valid_out_NO_SHIFT_REG;
wire local_bb6_st_c0_exe1108_stall_in;
wire local_bb6_st_c0_exe1108_output_regs_ready;
wire local_bb6_st_c0_exe1108_fu_stall_out;
wire local_bb6_st_c0_exe1108_fu_valid_out;
wire [31:0] local_bb6_st_c0_exe1108_lsu_wackout;
 reg local_bb6_st_c0_exe1108_NO_SHIFT_REG;
wire local_bb6_st_c0_exe1108_causedstall;

lsu_top lsu_local_bb6_st_c0_exe1108 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb6_st_c0_exe1108_fu_stall_out),
	.i_valid(local_bb6_st_c0_exe1108_inputs_ready),
	.i_address((rnode_20to21_bb6_arrayidx40_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(local_bb6_c0_exe1108),
	.i_cmpdata(),
	.i_predicate(input_wii_var_),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb6_st_c0_exe1108_output_regs_ready)),
	.o_valid(local_bb6_st_c0_exe1108_fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(local_bb6_st_c0_exe1108_lsu_wackout),
	.i_atomic_op(3'h0),
	.o_active(local_bb6_st_c0_exe1108_active),
	.avm_address(avm_local_bb6_st_c0_exe1108_address),
	.avm_read(avm_local_bb6_st_c0_exe1108_read),
	.avm_readdata(avm_local_bb6_st_c0_exe1108_readdata),
	.avm_write(avm_local_bb6_st_c0_exe1108_write),
	.avm_writeack(avm_local_bb6_st_c0_exe1108_writeack),
	.avm_burstcount(avm_local_bb6_st_c0_exe1108_burstcount),
	.avm_writedata(avm_local_bb6_st_c0_exe1108_writedata),
	.avm_byteenable(avm_local_bb6_st_c0_exe1108_byteenable),
	.avm_waitrequest(avm_local_bb6_st_c0_exe1108_waitrequest),
	.avm_readdatavalid(avm_local_bb6_st_c0_exe1108_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb6_st_c0_exe1108.AWIDTH = 33;
defparam lsu_local_bb6_st_c0_exe1108.WIDTH_BYTES = 4;
defparam lsu_local_bb6_st_c0_exe1108.MWIDTH_BYTES = 64;
defparam lsu_local_bb6_st_c0_exe1108.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb6_st_c0_exe1108.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb6_st_c0_exe1108.READ = 0;
defparam lsu_local_bb6_st_c0_exe1108.ATOMIC = 0;
defparam lsu_local_bb6_st_c0_exe1108.WIDTH = 32;
defparam lsu_local_bb6_st_c0_exe1108.MWIDTH = 512;
defparam lsu_local_bb6_st_c0_exe1108.ATOMIC_WIDTH = 3;
defparam lsu_local_bb6_st_c0_exe1108.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb6_st_c0_exe1108.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb6_st_c0_exe1108.MEMORY_SIDE_MEM_LATENCY = 8;
defparam lsu_local_bb6_st_c0_exe1108.USE_WRITE_ACK = 1;
defparam lsu_local_bb6_st_c0_exe1108.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb6_st_c0_exe1108.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb6_st_c0_exe1108.NUMBER_BANKS = 1;
defparam lsu_local_bb6_st_c0_exe1108.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb6_st_c0_exe1108.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb6_st_c0_exe1108.USEINPUTFIFO = 0;
defparam lsu_local_bb6_st_c0_exe1108.USECACHING = 0;
defparam lsu_local_bb6_st_c0_exe1108.USEOUTPUTFIFO = 1;
defparam lsu_local_bb6_st_c0_exe1108.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb6_st_c0_exe1108.HIGH_FMAX = 1;
defparam lsu_local_bb6_st_c0_exe1108.ADDRSPACE = 1;
defparam lsu_local_bb6_st_c0_exe1108.STYLE = "BURST-COALESCED";
defparam lsu_local_bb6_st_c0_exe1108.USE_BYTE_EN = 0;

assign local_bb6_st_c0_exe1108_inputs_ready = (local_bb6_c0_exe1108_valid_out & rnode_20to21_bb6_arrayidx40_0_valid_out_NO_SHIFT_REG & rnode_20to21_var__0_valid_out_NO_SHIFT_REG);
assign local_bb6_st_c0_exe1108_output_regs_ready = (&(~(local_bb6_st_c0_exe1108_valid_out_NO_SHIFT_REG) | ~(local_bb6_st_c0_exe1108_stall_in)));
assign local_bb6_c0_exe1108_stall_in = (local_bb6_st_c0_exe1108_fu_stall_out | ~(local_bb6_st_c0_exe1108_inputs_ready));
assign rnode_20to21_bb6_arrayidx40_0_stall_in_NO_SHIFT_REG = (local_bb6_st_c0_exe1108_fu_stall_out | ~(local_bb6_st_c0_exe1108_inputs_ready));
assign rnode_20to21_var__0_stall_in_NO_SHIFT_REG = (local_bb6_st_c0_exe1108_fu_stall_out | ~(local_bb6_st_c0_exe1108_inputs_ready));
assign local_bb6_st_c0_exe1108_causedstall = (local_bb6_st_c0_exe1108_inputs_ready && (local_bb6_st_c0_exe1108_fu_stall_out && !(~(local_bb6_st_c0_exe1108_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_st_c0_exe1108_NO_SHIFT_REG <= 'x;
		local_bb6_st_c0_exe1108_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_st_c0_exe1108_output_regs_ready)
		begin
			local_bb6_st_c0_exe1108_NO_SHIFT_REG <= local_bb6_st_c0_exe1108_lsu_wackout;
			local_bb6_st_c0_exe1108_valid_out_NO_SHIFT_REG <= local_bb6_st_c0_exe1108_fu_valid_out;
		end
		else
		begin
			if (~(local_bb6_st_c0_exe1108_stall_in))
			begin
				local_bb6_st_c0_exe1108_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_181to181_bb6_st_c0_exe1108_valid_out_0;
wire rstag_181to181_bb6_st_c0_exe1108_stall_in_0;
wire rstag_181to181_bb6_st_c0_exe1108_valid_out_1;
wire rstag_181to181_bb6_st_c0_exe1108_stall_in_1;
wire rstag_181to181_bb6_st_c0_exe1108_inputs_ready;
wire rstag_181to181_bb6_st_c0_exe1108_stall_local;
 reg rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG;
wire rstag_181to181_bb6_st_c0_exe1108_combined_valid;
 reg rstag_181to181_bb6_st_c0_exe1108_staging_reg_NO_SHIFT_REG;
wire rstag_181to181_bb6_st_c0_exe1108;
 reg rstag_181to181_bb6_st_c0_exe1108_consumed_0_NO_SHIFT_REG;
 reg rstag_181to181_bb6_st_c0_exe1108_consumed_1_NO_SHIFT_REG;
wire [3:0] rci_rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_181;

assign rstag_181to181_bb6_st_c0_exe1108_inputs_ready = local_bb6_st_c0_exe1108_valid_out_NO_SHIFT_REG;
assign rstag_181to181_bb6_st_c0_exe1108 = (rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG ? rstag_181to181_bb6_st_c0_exe1108_staging_reg_NO_SHIFT_REG : local_bb6_st_c0_exe1108_NO_SHIFT_REG);
assign rstag_181to181_bb6_st_c0_exe1108_combined_valid = (rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG | rstag_181to181_bb6_st_c0_exe1108_inputs_ready);
assign rstag_181to181_bb6_st_c0_exe1108_stall_local = ((rstag_181to181_bb6_st_c0_exe1108_stall_in_0 & ~(rstag_181to181_bb6_st_c0_exe1108_consumed_0_NO_SHIFT_REG)) | (rstag_181to181_bb6_st_c0_exe1108_stall_in_1 & ~(rstag_181to181_bb6_st_c0_exe1108_consumed_1_NO_SHIFT_REG)));
assign rstag_181to181_bb6_st_c0_exe1108_valid_out_0 = (rstag_181to181_bb6_st_c0_exe1108_combined_valid & ~(rstag_181to181_bb6_st_c0_exe1108_consumed_0_NO_SHIFT_REG));
assign rstag_181to181_bb6_st_c0_exe1108_valid_out_1 = (rstag_181to181_bb6_st_c0_exe1108_combined_valid & ~(rstag_181to181_bb6_st_c0_exe1108_consumed_1_NO_SHIFT_REG));
assign local_bb6_st_c0_exe1108_stall_in = (|rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG);
assign rci_rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_181[0] = rstag_181to181_bb6_st_c0_exe1108;
assign rci_rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_181[1] = rcnode_1to181_rc6_c0_exe895_0_NO_SHIFT_REG[0];
assign rci_rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_181[2] = rcnode_1to181_rc6_c0_exe895_0_NO_SHIFT_REG[1];
assign rci_rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_181[3] = rcnode_1to181_rc6_c0_exe895_0_NO_SHIFT_REG[2];

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_181to181_bb6_st_c0_exe1108_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_181to181_bb6_st_c0_exe1108_stall_local)
		begin
			if (~(rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG))
			begin
				rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG <= rstag_181to181_bb6_st_c0_exe1108_inputs_ready;
			end
		end
		else
		begin
			rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_181to181_bb6_st_c0_exe1108_staging_valid_NO_SHIFT_REG))
		begin
			rstag_181to181_bb6_st_c0_exe1108_staging_reg_NO_SHIFT_REG <= local_bb6_st_c0_exe1108_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_181to181_bb6_st_c0_exe1108_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_181to181_bb6_st_c0_exe1108_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_181to181_bb6_st_c0_exe1108_consumed_0_NO_SHIFT_REG <= (rstag_181to181_bb6_st_c0_exe1108_combined_valid & (rstag_181to181_bb6_st_c0_exe1108_consumed_0_NO_SHIFT_REG | ~(rstag_181to181_bb6_st_c0_exe1108_stall_in_0)) & rstag_181to181_bb6_st_c0_exe1108_stall_local);
		rstag_181to181_bb6_st_c0_exe1108_consumed_1_NO_SHIFT_REG <= (rstag_181to181_bb6_st_c0_exe1108_combined_valid & (rstag_181to181_bb6_st_c0_exe1108_consumed_1_NO_SHIFT_REG | ~(rstag_181to181_bb6_st_c0_exe1108_stall_in_1)) & rstag_181to181_bb6_st_c0_exe1108_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_181to182_rc0_bb6_st_c0_exe1108_0_valid_out_NO_SHIFT_REG;
 logic rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_in_NO_SHIFT_REG;
 logic [3:0] rcnode_181to182_rc0_bb6_st_c0_exe1108_0_NO_SHIFT_REG;
 logic rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [3:0] rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_NO_SHIFT_REG;
 logic rcnode_181to182_rc0_bb6_st_c0_exe1108_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_out_0_reg_182_IP_NO_SHIFT_REG;
 logic rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_out_0_reg_182_NO_SHIFT_REG;

acl_data_fifo rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rcnode_181to182_rc0_bb6_st_c0_exe1108_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_out_0_reg_182_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_181),
	.data_out(rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_NO_SHIFT_REG)
);

defparam rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_fifo.DEPTH = 1;
defparam rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_fifo.DATA_WIDTH = 4;
defparam rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_fifo.IMPL = "ll_reg";

assign rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_inputs_ready_NO_SHIFT_REG = (rcnode_1to181_rc6_c0_exe895_0_valid_out_NO_SHIFT_REG & rstag_181to181_bb6_st_c0_exe1108_valid_out_0);
assign rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_out_0_reg_182_NO_SHIFT_REG = (~(rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_inputs_ready_NO_SHIFT_REG) | rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_out_0_reg_182_IP_NO_SHIFT_REG);
assign rcnode_1to181_rc6_c0_exe895_0_stall_in_NO_SHIFT_REG = rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_out_0_reg_182_NO_SHIFT_REG;
assign rstag_181to181_bb6_st_c0_exe1108_stall_in_0 = rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_out_0_reg_182_NO_SHIFT_REG;
assign rcnode_181to182_rc0_bb6_st_c0_exe1108_0_NO_SHIFT_REG = rcnode_181to182_rc0_bb6_st_c0_exe1108_0_reg_182_NO_SHIFT_REG;
assign rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_in_reg_182_NO_SHIFT_REG = rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_in_NO_SHIFT_REG;
assign rcnode_181to182_rc0_bb6_st_c0_exe1108_0_valid_out_NO_SHIFT_REG = rcnode_181to182_rc0_bb6_st_c0_exe1108_0_valid_out_reg_182_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb6_memdep_phi_push11_memdep__inputs_ready;
 reg local_bb6_memdep_phi_push11_memdep__valid_out_NO_SHIFT_REG;
wire local_bb6_memdep_phi_push11_memdep__stall_in;
wire local_bb6_memdep_phi_push11_memdep__output_regs_ready;
wire local_bb6_memdep_phi_push11_memdep__result;
wire local_bb6_memdep_phi_push11_memdep__fu_valid_out;
wire local_bb6_memdep_phi_push11_memdep__fu_stall_out;
 reg local_bb6_memdep_phi_push11_memdep__NO_SHIFT_REG;
wire local_bb6_memdep_phi_push11_memdep__causedstall;

acl_push local_bb6_memdep_phi_push11_memdep__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_180to181_c0_exe1299_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rstag_181to181_bb6_st_c0_exe1108),
	.stall_out(local_bb6_memdep_phi_push11_memdep__fu_stall_out),
	.valid_in(local_bb6_memdep_phi_push11_memdep__inputs_ready),
	.valid_out(local_bb6_memdep_phi_push11_memdep__fu_valid_out),
	.stall_in(~(local_bb6_memdep_phi_push11_memdep__output_regs_ready)),
	.data_out(local_bb6_memdep_phi_push11_memdep__result),
	.feedback_out(feedback_data_out_11),
	.feedback_valid_out(feedback_valid_out_11),
	.feedback_stall_in(feedback_stall_in_11)
);

defparam local_bb6_memdep_phi_push11_memdep__feedback.STALLFREE = 0;
defparam local_bb6_memdep_phi_push11_memdep__feedback.DATA_WIDTH = 1;
defparam local_bb6_memdep_phi_push11_memdep__feedback.FIFO_DEPTH = 3;
defparam local_bb6_memdep_phi_push11_memdep__feedback.MIN_FIFO_LATENCY = 3;
defparam local_bb6_memdep_phi_push11_memdep__feedback.STYLE = "REGULAR";

assign local_bb6_memdep_phi_push11_memdep__inputs_ready = (rnode_180to181_c0_exe1299_0_valid_out_NO_SHIFT_REG & rstag_181to181_bb6_st_c0_exe1108_valid_out_1);
assign local_bb6_memdep_phi_push11_memdep__output_regs_ready = (&(~(local_bb6_memdep_phi_push11_memdep__valid_out_NO_SHIFT_REG) | ~(local_bb6_memdep_phi_push11_memdep__stall_in)));
assign rnode_180to181_c0_exe1299_0_stall_in_NO_SHIFT_REG = (local_bb6_memdep_phi_push11_memdep__fu_stall_out | ~(local_bb6_memdep_phi_push11_memdep__inputs_ready));
assign rstag_181to181_bb6_st_c0_exe1108_stall_in_1 = (local_bb6_memdep_phi_push11_memdep__fu_stall_out | ~(local_bb6_memdep_phi_push11_memdep__inputs_ready));
assign local_bb6_memdep_phi_push11_memdep__causedstall = (local_bb6_memdep_phi_push11_memdep__inputs_ready && (local_bb6_memdep_phi_push11_memdep__fu_stall_out && !(~(local_bb6_memdep_phi_push11_memdep__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_memdep_phi_push11_memdep__NO_SHIFT_REG <= 'x;
		local_bb6_memdep_phi_push11_memdep__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_memdep_phi_push11_memdep__output_regs_ready)
		begin
			local_bb6_memdep_phi_push11_memdep__NO_SHIFT_REG <= local_bb6_memdep_phi_push11_memdep__result;
			local_bb6_memdep_phi_push11_memdep__valid_out_NO_SHIFT_REG <= local_bb6_memdep_phi_push11_memdep__fu_valid_out;
		end
		else
		begin
			if (~(local_bb6_memdep_phi_push11_memdep__stall_in))
			begin
				local_bb6_memdep_phi_push11_memdep__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg lvb_c0_exe895_0_reg_NO_SHIFT_REG;
 reg lvb_c0_exe996_0_reg_NO_SHIFT_REG;
 reg lvb_bb6_st_c0_exe1108_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb6_memdep_phi_push11_memdep__valid_out_NO_SHIFT_REG & rcnode_181to182_rc0_bb6_st_c0_exe1108_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb6_memdep_phi_push11_memdep__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_181to182_rc0_bb6_st_c0_exe1108_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_c0_exe895_0 = lvb_c0_exe895_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe895_1 = lvb_c0_exe895_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe996_0 = lvb_c0_exe996_0_reg_NO_SHIFT_REG;
assign lvb_c0_exe996_1 = lvb_c0_exe996_0_reg_NO_SHIFT_REG;
assign lvb_bb6_st_c0_exe1108_0 = lvb_bb6_st_c0_exe1108_0_reg_NO_SHIFT_REG;
assign lvb_bb6_st_c0_exe1108_1 = lvb_bb6_st_c0_exe1108_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_c0_exe895_0_reg_NO_SHIFT_REG <= 'x;
		lvb_c0_exe996_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb6_st_c0_exe1108_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_c0_exe895_0_reg_NO_SHIFT_REG <= rcnode_181to182_rc0_bb6_st_c0_exe1108_0_NO_SHIFT_REG[1];
			lvb_c0_exe996_0_reg_NO_SHIFT_REG <= rcnode_181to182_rc0_bb6_st_c0_exe1108_0_NO_SHIFT_REG[2];
			lvb_bb6_st_c0_exe1108_0_reg_NO_SHIFT_REG <= rcnode_181to182_rc0_bb6_st_c0_exe1108_0_NO_SHIFT_REG[0];
			branch_compare_result_NO_SHIFT_REG <= rcnode_181to182_rc0_bb6_st_c0_exe1108_0_NO_SHIFT_REG[3];
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_7
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_wii_div,
		input [31:0] 		input_wii_div1,
		input 		input_wii_cmp19,
		input [31:0] 		input_wii_add7,
		input [31:0] 		input_wii_sub20,
		input [31:0] 		input_wii_sub22,
		input 		input_wii_var_,
		input 		input_wii_var__u64,
		input 		input_wii_var__u65,
		input 		input_wii_var__u66,
		input 		valid_in,
		output 		stall_out,
		input 		input_c0_exe895,
		input 		input_c0_exe996,
		input 		input_st_c0_exe1108,
		output 		valid_out_0,
		input 		stall_in_0,
		output 		valid_out_1,
		input 		stall_in_1,
		input [31:0] 		workgroup_size,
		input 		start,
		output 		feedback_valid_out_9,
		input 		feedback_stall_in_9,
		output 		feedback_data_out_9
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe895_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe996_staging_reg_NO_SHIFT_REG;
 reg input_st_c0_exe1108_staging_reg_NO_SHIFT_REG;
 reg local_lvm_c0_exe895_NO_SHIFT_REG;
 reg local_lvm_c0_exe996_NO_SHIFT_REG;
 reg local_lvm_st_c0_exe1108_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_c0_exe895_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe996_staging_reg_NO_SHIFT_REG <= 'x;
		input_st_c0_exe1108_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_c0_exe895_staging_reg_NO_SHIFT_REG <= input_c0_exe895;
				input_c0_exe996_staging_reg_NO_SHIFT_REG <= input_c0_exe996;
				input_st_c0_exe1108_staging_reg_NO_SHIFT_REG <= input_st_c0_exe1108;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_c0_exe895_NO_SHIFT_REG <= input_c0_exe895_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe996_NO_SHIFT_REG <= input_c0_exe996_staging_reg_NO_SHIFT_REG;
					local_lvm_st_c0_exe1108_NO_SHIFT_REG <= input_st_c0_exe1108_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_c0_exe895_NO_SHIFT_REG <= input_c0_exe895;
					local_lvm_c0_exe996_NO_SHIFT_REG <= input_c0_exe996;
					local_lvm_st_c0_exe1108_NO_SHIFT_REG <= input_st_c0_exe1108;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb7_memdep_phi1_push9_memdep__inputs_ready;
 reg local_bb7_memdep_phi1_push9_memdep__valid_out_NO_SHIFT_REG;
wire local_bb7_memdep_phi1_push9_memdep__stall_in;
wire local_bb7_memdep_phi1_push9_memdep__output_regs_ready;
wire local_bb7_memdep_phi1_push9_memdep__result;
wire local_bb7_memdep_phi1_push9_memdep__fu_valid_out;
wire local_bb7_memdep_phi1_push9_memdep__fu_stall_out;
 reg local_bb7_memdep_phi1_push9_memdep__NO_SHIFT_REG;
wire local_bb7_memdep_phi1_push9_memdep__causedstall;

acl_push local_bb7_memdep_phi1_push9_memdep__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_c0_exe996_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_lvm_st_c0_exe1108_NO_SHIFT_REG),
	.stall_out(local_bb7_memdep_phi1_push9_memdep__fu_stall_out),
	.valid_in(local_bb7_memdep_phi1_push9_memdep__inputs_ready),
	.valid_out(local_bb7_memdep_phi1_push9_memdep__fu_valid_out),
	.stall_in(~(local_bb7_memdep_phi1_push9_memdep__output_regs_ready)),
	.data_out(local_bb7_memdep_phi1_push9_memdep__result),
	.feedback_out(feedback_data_out_9),
	.feedback_valid_out(feedback_valid_out_9),
	.feedback_stall_in(feedback_stall_in_9)
);

defparam local_bb7_memdep_phi1_push9_memdep__feedback.STALLFREE = 0;
defparam local_bb7_memdep_phi1_push9_memdep__feedback.DATA_WIDTH = 1;
defparam local_bb7_memdep_phi1_push9_memdep__feedback.FIFO_DEPTH = 3;
defparam local_bb7_memdep_phi1_push9_memdep__feedback.MIN_FIFO_LATENCY = 3;
defparam local_bb7_memdep_phi1_push9_memdep__feedback.STYLE = "REGULAR";

assign local_bb7_memdep_phi1_push9_memdep__inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb7_memdep_phi1_push9_memdep__output_regs_ready = (&(~(local_bb7_memdep_phi1_push9_memdep__valid_out_NO_SHIFT_REG) | ~(local_bb7_memdep_phi1_push9_memdep__stall_in)));
assign merge_node_stall_in_0 = (local_bb7_memdep_phi1_push9_memdep__fu_stall_out | ~(local_bb7_memdep_phi1_push9_memdep__inputs_ready));
assign local_bb7_memdep_phi1_push9_memdep__causedstall = (local_bb7_memdep_phi1_push9_memdep__inputs_ready && (local_bb7_memdep_phi1_push9_memdep__fu_stall_out && !(~(local_bb7_memdep_phi1_push9_memdep__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb7_memdep_phi1_push9_memdep__NO_SHIFT_REG <= 'x;
		local_bb7_memdep_phi1_push9_memdep__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb7_memdep_phi1_push9_memdep__output_regs_ready)
		begin
			local_bb7_memdep_phi1_push9_memdep__NO_SHIFT_REG <= local_bb7_memdep_phi1_push9_memdep__result;
			local_bb7_memdep_phi1_push9_memdep__valid_out_NO_SHIFT_REG <= local_bb7_memdep_phi1_push9_memdep__fu_valid_out;
		end
		else
		begin
			if (~(local_bb7_memdep_phi1_push9_memdep__stall_in))
			begin
				local_bb7_memdep_phi1_push9_memdep__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_c0_exe895_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_c0_exe895_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_c0_exe895_0_NO_SHIFT_REG;
 logic rnode_1to2_c0_exe895_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_c0_exe895_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_c0_exe895_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_c0_exe895_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_c0_exe895_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_c0_exe895_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_c0_exe895_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_c0_exe895_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_c0_exe895_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_c0_exe895_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_lvm_c0_exe895_NO_SHIFT_REG),
	.data_out(rnode_1to2_c0_exe895_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_c0_exe895_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_c0_exe895_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_c0_exe895_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_c0_exe895_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_c0_exe895_0_reg_2_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign merge_node_stall_in_1 = rnode_1to2_c0_exe895_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_c0_exe895_0_NO_SHIFT_REG = rnode_1to2_c0_exe895_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_c0_exe895_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_c0_exe895_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_c0_exe895_0_valid_out_NO_SHIFT_REG = rnode_1to2_c0_exe895_0_valid_out_reg_2_NO_SHIFT_REG;

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;

assign branch_var__inputs_ready = (local_bb7_memdep_phi1_push9_memdep__valid_out_NO_SHIFT_REG & rnode_1to2_c0_exe895_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb7_memdep_phi1_push9_memdep__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to2_c0_exe895_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			branch_compare_result_NO_SHIFT_REG <= rnode_1to2_c0_exe895_0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_basic_block_8
	(
		input 		clock,
		input 		resetn,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in;
 reg merge_node_valid_out_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = (|(merge_node_stall_in & merge_node_valid_out_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in))
			begin
				merge_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
wire branch_var__output_regs_ready;

assign branch_var__inputs_ready = merge_node_valid_out_NO_SHIFT_REG;
assign branch_var__output_regs_ready = ~(stall_in);
assign merge_node_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out = branch_var__inputs_ready;

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_function
	(
		input 		clock,
		input 		resetn,
		output 		stall_out,
		input 		valid_in,
		output 		valid_out,
		input 		stall_in,
		input [511:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [32:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [511:0] 		avm_local_bb2_ld__writedata,
		output [63:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		input [511:0] 		avm_local_bb4_ld__readdata,
		input 		avm_local_bb4_ld__readdatavalid,
		input 		avm_local_bb4_ld__waitrequest,
		output [32:0] 		avm_local_bb4_ld__address,
		output 		avm_local_bb4_ld__read,
		output 		avm_local_bb4_ld__write,
		input 		avm_local_bb4_ld__writeack,
		output [511:0] 		avm_local_bb4_ld__writedata,
		output [63:0] 		avm_local_bb4_ld__byteenable,
		output [4:0] 		avm_local_bb4_ld__burstcount,
		input [511:0] 		avm_local_bb6_st_c0_exe1108_readdata,
		input 		avm_local_bb6_st_c0_exe1108_readdatavalid,
		input 		avm_local_bb6_st_c0_exe1108_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe1108_address,
		output 		avm_local_bb6_st_c0_exe1108_read,
		output 		avm_local_bb6_st_c0_exe1108_write,
		input 		avm_local_bb6_st_c0_exe1108_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe1108_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe1108_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe1108_burstcount,
		input 		start,
		input [31:0] 		input_inSize_x,
		input [31:0] 		input_inSize_y,
		input [31:0] 		input_r,
		input 		clock2x,
		input [63:0] 		input_in,
		input [31:0] 		input_e_d,
		input [63:0] 		input_out,
		output reg 		has_a_write_pending,
		output reg 		has_a_lsu_active
	);


wire [31:0] workgroup_size;
wire [31:0] cur_cycle;
wire bb_0_stall_out;
wire bb_0_valid_out;
wire [31:0] bb_0_lvb_bb0_div;
wire [31:0] bb_0_lvb_bb0_div1;
wire bb_0_lvb_bb0_cmp19;
wire [31:0] bb_0_lvb_bb0_add7;
wire [31:0] bb_0_lvb_bb0_sub20;
wire [31:0] bb_0_lvb_bb0_sub22;
wire bb_0_lvb_bb0_var_;
wire bb_0_lvb_bb0_var__u0;
wire bb_0_lvb_bb0_var__u1;
wire bb_0_lvb_bb0_var__u2;
wire bb_1_stall_out_0;
wire bb_1_stall_out_1;
wire bb_1_valid_out;
wire [31:0] bb_1_lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0;
wire [31:0] bb_1_lvb_bb1_mul37;
wire bb_1_lvb_bb1_notcmp11;
wire bb_1_lvb_bb1_notexitcond14_;
wire bb_1_lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0;
wire bb_1_feedback_stall_out_8;
wire bb_1_feedback_stall_out_9;
wire bb_1_feedback_stall_out_6;
wire bb_1_feedback_stall_out_7;
wire bb_1_acl_pipelined_valid;
wire bb_1_acl_pipelined_exiting_valid;
wire bb_1_acl_pipelined_exiting_stall;
wire bb_1_feedback_valid_out_8;
wire [31:0] bb_1_feedback_data_out_8;
wire bb_1_feedback_valid_out_7;
wire bb_1_feedback_data_out_7;
wire bb_2_stall_out_0;
wire bb_2_stall_out_1;
wire bb_2_valid_out;
wire [31:0] bb_2_lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819;
wire [31:0] bb_2_lvb_bb2_mul5;
wire [63:0] bb_2_lvb_bb2_indvars_iv_pop10_acl_pop_i64_0;
wire [31:0] bb_2_lvb_bb2_var_;
wire bb_2_lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931;
wire bb_2_lvb_bb2_memdep_phi1_or;
wire [31:0] bb_2_lvb_bb2_ld_;
wire bb_2_lvb_bb2_notcmp;
wire bb_2_lvb_bb2_notexitcond9_;
wire [31:0] bb_2_lvb_bb2_mul3722_pop13_mul3722;
wire bb_2_lvb_bb2_notcmp1125_pop14_notcmp1125;
wire bb_2_lvb_bb2_notexitcond1428_pop15_notexitcond1428;
wire bb_2_feedback_stall_out_12;
wire bb_2_feedback_stall_out_10;
wire bb_2_feedback_stall_out_4;
wire bb_2_feedback_stall_out_5;
wire bb_2_acl_pipelined_valid;
wire bb_2_acl_pipelined_exiting_valid;
wire bb_2_acl_pipelined_exiting_stall;
wire bb_2_feedback_stall_out_11;
wire bb_2_feedback_stall_out_16;
wire bb_2_feedback_stall_out_13;
wire bb_2_feedback_stall_out_14;
wire bb_2_feedback_stall_out_15;
wire bb_2_feedback_valid_out_10;
wire [63:0] bb_2_feedback_data_out_10;
wire bb_2_feedback_valid_out_5;
wire bb_2_feedback_data_out_5;
wire bb_2_feedback_valid_out_12;
wire [31:0] bb_2_feedback_data_out_12;
wire bb_2_feedback_valid_out_16;
wire bb_2_feedback_data_out_16;
wire bb_2_feedback_valid_out_13;
wire [31:0] bb_2_feedback_data_out_13;
wire bb_2_feedback_valid_out_14;
wire bb_2_feedback_data_out_14;
wire bb_2_feedback_valid_out_15;
wire bb_2_feedback_data_out_15;
wire bb_2_local_bb2_ld__active;
wire bb_3_stall_out_0;
wire bb_3_stall_out_1;
wire bb_3_valid_out;
wire bb_3_lvb_forked16;
wire [31:0] bb_3_lvb_bb3_c0_exe1;
wire [31:0] bb_3_lvb_bb3_c0_exe2;
wire bb_3_lvb_bb3_c0_exe3;
wire bb_3_lvb_bb3_c0_exe4;
wire [31:0] bb_3_lvb_bb3_c0_exe5;
wire [31:0] bb_3_lvb_bb3_c0_exe6;
wire bb_3_lvb_bb3_c0_exe7;
wire bb_3_lvb_bb3_c0_exe8;
wire bb_3_lvb_bb3_c0_exe9;
wire [63:0] bb_3_lvb_bb3_c0_exe10;
wire [31:0] bb_3_lvb_bb3_c0_exe11;
wire bb_3_lvb_bb3_c0_exe12;
wire [31:0] bb_3_lvb_bb3_c0_exe13;
wire bb_3_lvb_bb3_c0_exe14;
wire bb_3_lvb_bb3_c0_exe15;
wire bb_3_feedback_stall_out_17;
wire bb_3_feedback_stall_out_23;
wire bb_3_feedback_stall_out_2;
wire bb_3_feedback_stall_out_3;
wire bb_3_acl_pipelined_valid;
wire bb_3_acl_pipelined_exiting_valid;
wire bb_3_acl_pipelined_exiting_stall;
wire bb_3_feedback_stall_out_18;
wire bb_3_feedback_stall_out_19;
wire bb_3_feedback_stall_out_20;
wire bb_3_feedback_stall_out_21;
wire bb_3_feedback_stall_out_22;
wire bb_3_feedback_stall_out_24;
wire bb_3_feedback_stall_out_25;
wire bb_3_feedback_stall_out_26;
wire bb_3_feedback_stall_out_27;
wire bb_3_feedback_stall_out_28;
wire bb_3_feedback_stall_out_29;
wire bb_3_feedback_valid_out_3;
wire bb_3_feedback_data_out_3;
wire bb_3_feedback_valid_out_17;
wire [31:0] bb_3_feedback_data_out_17;
wire bb_3_feedback_valid_out_23;
wire [31:0] bb_3_feedback_data_out_23;
wire bb_3_feedback_valid_out_18;
wire [31:0] bb_3_feedback_data_out_18;
wire bb_3_feedback_valid_out_19;
wire [31:0] bb_3_feedback_data_out_19;
wire bb_3_feedback_valid_out_20;
wire bb_3_feedback_data_out_20;
wire bb_3_feedback_valid_out_21;
wire bb_3_feedback_data_out_21;
wire bb_3_feedback_valid_out_22;
wire bb_3_feedback_data_out_22;
wire bb_3_feedback_valid_out_24;
wire [63:0] bb_3_feedback_data_out_24;
wire bb_3_feedback_valid_out_25;
wire [31:0] bb_3_feedback_data_out_25;
wire bb_3_feedback_valid_out_26;
wire bb_3_feedback_data_out_26;
wire bb_3_feedback_valid_out_27;
wire [31:0] bb_3_feedback_data_out_27;
wire bb_3_feedback_valid_out_28;
wire bb_3_feedback_data_out_28;
wire bb_3_feedback_valid_out_29;
wire bb_3_feedback_data_out_29;
wire bb_4_stall_out_0;
wire bb_4_stall_out_1;
wire bb_4_valid_out_0;
wire [447:0] bb_4_lvb_bb4_c0_exit87_c0_exi1386_0;
wire [31:0] bb_4_lvb_bb4_c0_exe794_0;
wire bb_4_lvb_bb4_c0_exe895_0;
wire bb_4_lvb_bb4_c0_exe996_0;
wire [63:0] bb_4_lvb_bb4_c0_exe1097_0;
wire bb_4_lvb_bb4_c0_exe1198_0;
wire bb_4_lvb_bb4_c0_exe1299_0;
wire [31:0] bb_4_lvb_bb4_c1_exe1_0;
wire [31:0] bb_4_lvb_bb4_c1_exe2_0;
wire bb_4_valid_out_1;
wire [447:0] bb_4_lvb_bb4_c0_exit87_c0_exi1386_1;
wire [31:0] bb_4_lvb_bb4_c0_exe794_1;
wire bb_4_lvb_bb4_c0_exe895_1;
wire bb_4_lvb_bb4_c0_exe996_1;
wire [63:0] bb_4_lvb_bb4_c0_exe1097_1;
wire bb_4_lvb_bb4_c0_exe1198_1;
wire bb_4_lvb_bb4_c0_exe1299_1;
wire [31:0] bb_4_lvb_bb4_c1_exe1_1;
wire [31:0] bb_4_lvb_bb4_c1_exe2_1;
wire bb_4_feedback_stall_out_30;
wire bb_4_feedback_stall_out_40;
wire bb_4_feedback_stall_out_0;
wire bb_4_feedback_stall_out_1;
wire bb_4_acl_pipelined_valid;
wire bb_4_acl_pipelined_exiting_valid;
wire bb_4_acl_pipelined_exiting_stall;
wire bb_4_feedback_stall_out_46;
wire bb_4_feedback_stall_out_45;
wire bb_4_feedback_stall_out_41;
wire bb_4_feedback_stall_out_42;
wire bb_4_feedback_stall_out_33;
wire bb_4_feedback_stall_out_34;
wire bb_4_feedback_stall_out_35;
wire bb_4_feedback_stall_out_36;
wire bb_4_feedback_stall_out_37;
wire bb_4_feedback_stall_out_38;
wire bb_4_feedback_stall_out_39;
wire bb_4_feedback_stall_out_43;
wire bb_4_feedback_stall_out_44;
wire bb_4_feedback_stall_out_47;
wire bb_4_feedback_valid_out_1;
wire bb_4_feedback_data_out_1;
wire bb_4_feedback_valid_out_30;
wire [31:0] bb_4_feedback_data_out_30;
wire bb_4_feedback_valid_out_45;
wire bb_4_feedback_data_out_45;
wire bb_4_feedback_valid_out_42;
wire [31:0] bb_4_feedback_data_out_42;
wire bb_4_feedback_valid_out_41;
wire bb_4_feedback_data_out_41;
wire bb_4_feedback_valid_out_40;
wire [31:0] bb_4_feedback_data_out_40;
wire bb_4_feedback_valid_out_33;
wire [31:0] bb_4_feedback_data_out_33;
wire bb_4_feedback_valid_out_34;
wire [31:0] bb_4_feedback_data_out_34;
wire bb_4_feedback_valid_out_35;
wire bb_4_feedback_data_out_35;
wire bb_4_feedback_valid_out_36;
wire bb_4_feedback_data_out_36;
wire bb_4_feedback_valid_out_37;
wire bb_4_feedback_data_out_37;
wire bb_4_feedback_valid_out_38;
wire [31:0] bb_4_feedback_data_out_38;
wire bb_4_feedback_valid_out_39;
wire [63:0] bb_4_feedback_data_out_39;
wire bb_4_feedback_valid_out_43;
wire bb_4_feedback_data_out_43;
wire bb_4_feedback_valid_out_44;
wire bb_4_feedback_data_out_44;
wire bb_4_feedback_valid_out_47;
wire bb_4_feedback_data_out_47;
wire bb_4_feedback_valid_out_46;
wire [31:0] bb_4_feedback_data_out_46;
wire bb_4_local_bb4_ld__active;
wire bb_4_feedback_stall_out_48;
wire bb_4_feedback_valid_out_48;
wire bb_4_feedback_data_out_48;
wire bb_4_feedback_stall_out_31;
wire bb_4_feedback_stall_out_32;
wire bb_4_feedback_valid_out_32;
wire [31:0] bb_4_feedback_data_out_32;
wire bb_4_feedback_valid_out_31;
wire [31:0] bb_4_feedback_data_out_31;
wire bb_5_stall_out;
wire bb_5_valid_out_0;
wire [31:0] bb_5_lvb_c0_exe794_0;
wire bb_5_lvb_c0_exe895_0;
wire bb_5_lvb_c0_exe996_0;
wire [63:0] bb_5_lvb_c0_exe1097_0;
wire bb_5_lvb_c0_exe1198_0;
wire bb_5_lvb_c0_exe1299_0;
wire [31:0] bb_5_lvb_c1_exe1_0;
wire [31:0] bb_5_lvb_c1_exe2_0;
wire bb_5_valid_out_1;
wire [31:0] bb_5_lvb_c0_exe794_1;
wire bb_5_lvb_c0_exe895_1;
wire bb_5_lvb_c0_exe996_1;
wire [63:0] bb_5_lvb_c0_exe1097_1;
wire bb_5_lvb_c0_exe1198_1;
wire bb_5_lvb_c0_exe1299_1;
wire [31:0] bb_5_lvb_c1_exe1_1;
wire [31:0] bb_5_lvb_c1_exe2_1;
wire bb_6_stall_out;
wire bb_6_valid_out_0;
wire bb_6_lvb_c0_exe895_0;
wire bb_6_lvb_c0_exe996_0;
wire bb_6_lvb_bb6_st_c0_exe1108_0;
wire bb_6_valid_out_1;
wire bb_6_lvb_c0_exe895_1;
wire bb_6_lvb_c0_exe996_1;
wire bb_6_lvb_bb6_st_c0_exe1108_1;
wire bb_6_local_bb6_st_c0_exe1108_active;
wire bb_6_feedback_valid_out_11;
wire bb_6_feedback_data_out_11;
wire bb_7_stall_out;
wire bb_7_valid_out_0;
wire bb_7_valid_out_1;
wire bb_7_feedback_valid_out_9;
wire bb_7_feedback_data_out_9;
wire bb_8_stall_out;
wire bb_8_valid_out;
wire feedback_stall_7;
wire feedback_valid_7;
wire feedback_data_7;
wire feedback_stall_8;
wire feedback_valid_8;
wire [31:0] feedback_data_8;
wire feedback_stall_5;
wire feedback_valid_5;
wire feedback_data_5;
wire feedback_stall_16;
wire feedback_valid_16;
wire feedback_data_16;
wire feedback_stall_12;
wire feedback_valid_12;
wire [31:0] feedback_data_12;
wire feedback_stall_10;
wire feedback_valid_10;
wire [63:0] feedback_data_10;
wire feedback_stall_13;
wire feedback_valid_13;
wire [31:0] feedback_data_13;
wire feedback_stall_14;
wire feedback_valid_14;
wire feedback_data_14;
wire feedback_stall_15;
wire feedback_valid_15;
wire feedback_data_15;
wire feedback_stall_3;
wire feedback_valid_3;
wire feedback_data_3;
wire feedback_stall_23;
wire feedback_valid_23;
wire [31:0] feedback_data_23;
wire feedback_stall_17;
wire feedback_valid_17;
wire [31:0] feedback_data_17;
wire feedback_stall_18;
wire feedback_valid_18;
wire [31:0] feedback_data_18;
wire feedback_stall_19;
wire feedback_valid_19;
wire [31:0] feedback_data_19;
wire feedback_stall_20;
wire feedback_valid_20;
wire feedback_data_20;
wire feedback_stall_21;
wire feedback_valid_21;
wire feedback_data_21;
wire feedback_stall_22;
wire feedback_valid_22;
wire feedback_data_22;
wire feedback_stall_24;
wire feedback_valid_24;
wire [63:0] feedback_data_24;
wire feedback_stall_25;
wire feedback_valid_25;
wire [31:0] feedback_data_25;
wire feedback_stall_26;
wire feedback_valid_26;
wire feedback_data_26;
wire feedback_stall_27;
wire feedback_valid_27;
wire [31:0] feedback_data_27;
wire feedback_stall_28;
wire feedback_valid_28;
wire feedback_data_28;
wire feedback_stall_29;
wire feedback_valid_29;
wire feedback_data_29;
wire feedback_stall_1;
wire feedback_valid_1;
wire feedback_data_1;
wire feedback_stall_46;
wire feedback_valid_46;
wire [31:0] feedback_data_46;
wire feedback_stall_45;
wire feedback_valid_45;
wire feedback_data_45;
wire feedback_stall_42;
wire feedback_valid_42;
wire [31:0] feedback_data_42;
wire feedback_stall_41;
wire feedback_valid_41;
wire feedback_data_41;
wire feedback_stall_40;
wire feedback_valid_40;
wire [31:0] feedback_data_40;
wire feedback_stall_30;
wire feedback_valid_30;
wire [31:0] feedback_data_30;
wire feedback_stall_33;
wire feedback_valid_33;
wire [31:0] feedback_data_33;
wire feedback_stall_34;
wire feedback_valid_34;
wire [31:0] feedback_data_34;
wire feedback_stall_35;
wire feedback_valid_35;
wire feedback_data_35;
wire feedback_stall_36;
wire feedback_valid_36;
wire feedback_data_36;
wire feedback_stall_37;
wire feedback_valid_37;
wire feedback_data_37;
wire feedback_stall_38;
wire feedback_valid_38;
wire [31:0] feedback_data_38;
wire feedback_stall_39;
wire feedback_valid_39;
wire [63:0] feedback_data_39;
wire feedback_stall_43;
wire feedback_valid_43;
wire feedback_data_43;
wire feedback_stall_44;
wire feedback_valid_44;
wire feedback_data_44;
wire feedback_stall_47;
wire feedback_valid_47;
wire feedback_data_47;
wire feedback_stall_48;
wire feedback_valid_48;
wire feedback_data_48;
wire feedback_stall_32;
wire feedback_valid_32;
wire [31:0] feedback_data_32;
wire feedback_stall_31;
wire feedback_valid_31;
wire [31:0] feedback_data_31;
wire feedback_stall_11;
wire feedback_valid_11;
wire feedback_data_11;
wire feedback_stall_9;
wire feedback_valid_9;
wire feedback_data_9;
wire loop_limiter_1_stall_out;
wire loop_limiter_1_valid_out;
wire loop_limiter_2_stall_out;
wire loop_limiter_2_valid_out;
wire loop_limiter_3_stall_out;
wire loop_limiter_3_valid_out;
wire writes_pending;
wire [2:0] lsus_active;

AOChalfSampleRobustImageKernel_basic_block_0 AOChalfSampleRobustImageKernel_basic_block_0 (
	.clock(clock),
	.resetn(resetn),
	.start(start),
	.input_inSize_x(input_inSize_x),
	.input_inSize_y(input_inSize_y),
	.input_r(input_r),
	.valid_in(valid_in),
	.stall_out(bb_0_stall_out),
	.valid_out(bb_0_valid_out),
	.stall_in(bb_1_stall_out_1),
	.lvb_bb0_div(bb_0_lvb_bb0_div),
	.lvb_bb0_div1(bb_0_lvb_bb0_div1),
	.lvb_bb0_cmp19(bb_0_lvb_bb0_cmp19),
	.lvb_bb0_add7(bb_0_lvb_bb0_add7),
	.lvb_bb0_sub20(bb_0_lvb_bb0_sub20),
	.lvb_bb0_sub22(bb_0_lvb_bb0_sub22),
	.lvb_bb0_var_(bb_0_lvb_bb0_var_),
	.lvb_bb0_var__u0(bb_0_lvb_bb0_var__u0),
	.lvb_bb0_var__u1(bb_0_lvb_bb0_var__u1),
	.lvb_bb0_var__u2(bb_0_lvb_bb0_var__u2),
	.workgroup_size(workgroup_size)
);


AOChalfSampleRobustImageKernel_basic_block_1 AOChalfSampleRobustImageKernel_basic_block_1 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_div(bb_0_lvb_bb0_div),
	.input_wii_div1(bb_0_lvb_bb0_div1),
	.input_wii_cmp19(bb_0_lvb_bb0_cmp19),
	.input_wii_add7(bb_0_lvb_bb0_add7),
	.input_wii_sub20(bb_0_lvb_bb0_sub20),
	.input_wii_sub22(bb_0_lvb_bb0_sub22),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u3(bb_0_lvb_bb0_var__u0),
	.input_wii_var__u4(bb_0_lvb_bb0_var__u1),
	.input_wii_var__u5(bb_0_lvb_bb0_var__u2),
	.valid_in_0(bb_1_acl_pipelined_valid),
	.stall_out_0(bb_1_stall_out_0),
	.input_forked17_0(1'b0),
	.valid_in_1(bb_0_valid_out),
	.stall_out_1(bb_1_stall_out_1),
	.input_forked17_1(1'b1),
	.valid_out(bb_1_valid_out),
	.stall_in(loop_limiter_1_stall_out),
	.lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0(bb_1_lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0),
	.lvb_bb1_mul37(bb_1_lvb_bb1_mul37),
	.lvb_bb1_notcmp11(bb_1_lvb_bb1_notcmp11),
	.lvb_bb1_notexitcond14_(bb_1_lvb_bb1_notexitcond14_),
	.lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0(bb_1_lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_in_8(feedback_valid_8),
	.feedback_stall_out_8(feedback_stall_8),
	.feedback_data_in_8(feedback_data_8),
	.feedback_valid_in_9(feedback_valid_9),
	.feedback_stall_out_9(feedback_stall_9),
	.feedback_data_in_9(feedback_data_9),
	.feedback_stall_out_6(bb_1_feedback_stall_out_6),
	.feedback_valid_in_7(feedback_valid_7),
	.feedback_stall_out_7(feedback_stall_7),
	.feedback_data_in_7(feedback_data_7),
	.acl_pipelined_valid(bb_1_acl_pipelined_valid),
	.acl_pipelined_stall(bb_1_stall_out_0),
	.acl_pipelined_exiting_valid(bb_1_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_1_acl_pipelined_exiting_stall),
	.feedback_valid_out_8(feedback_valid_8),
	.feedback_stall_in_8(feedback_stall_8),
	.feedback_data_out_8(feedback_data_8),
	.feedback_valid_out_7(feedback_valid_7),
	.feedback_stall_in_7(feedback_stall_7),
	.feedback_data_out_7(feedback_data_7)
);


AOChalfSampleRobustImageKernel_basic_block_2 AOChalfSampleRobustImageKernel_basic_block_2 (
	.clock(clock),
	.resetn(resetn),
	.input_inSize_x(input_inSize_x),
	.input_in(input_in),
	.input_wii_div(bb_0_lvb_bb0_div),
	.input_wii_div1(bb_0_lvb_bb0_div1),
	.input_wii_cmp19(bb_0_lvb_bb0_cmp19),
	.input_wii_add7(bb_0_lvb_bb0_add7),
	.input_wii_sub20(bb_0_lvb_bb0_sub20),
	.input_wii_sub22(bb_0_lvb_bb0_sub22),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u6(bb_0_lvb_bb0_var__u0),
	.input_wii_var__u7(bb_0_lvb_bb0_var__u1),
	.input_wii_var__u8(bb_0_lvb_bb0_var__u2),
	.valid_in_0(bb_2_acl_pipelined_valid),
	.stall_out_0(bb_2_stall_out_0),
	.input_forked18_0(1'b0),
	.input_pixel_y_020_pop819_0('x),
	.input_mul3722_0('x),
	.input_notcmp1125_0('x),
	.input_notexitcond1428_0('x),
	.input_memdep_phi1_pop931_0('x),
	.valid_in_1(loop_limiter_1_valid_out),
	.stall_out_1(bb_2_stall_out_1),
	.input_forked18_1(1'b1),
	.input_pixel_y_020_pop819_1(bb_1_lvb_bb1_pixel_y_020_pop8_acl_pop_i32_0),
	.input_mul3722_1(bb_1_lvb_bb1_mul37),
	.input_notcmp1125_1(bb_1_lvb_bb1_notcmp11),
	.input_notexitcond1428_1(bb_1_lvb_bb1_notexitcond14_),
	.input_memdep_phi1_pop931_1(bb_1_lvb_bb1_memdep_phi1_pop9_acl_pop_i1_0),
	.valid_out(bb_2_valid_out),
	.stall_in(loop_limiter_2_stall_out),
	.lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819(bb_2_lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819),
	.lvb_bb2_mul5(bb_2_lvb_bb2_mul5),
	.lvb_bb2_indvars_iv_pop10_acl_pop_i64_0(bb_2_lvb_bb2_indvars_iv_pop10_acl_pop_i64_0),
	.lvb_bb2_var_(bb_2_lvb_bb2_var_),
	.lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931(bb_2_lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931),
	.lvb_bb2_memdep_phi1_or(bb_2_lvb_bb2_memdep_phi1_or),
	.lvb_bb2_ld_(bb_2_lvb_bb2_ld_),
	.lvb_bb2_notcmp(bb_2_lvb_bb2_notcmp),
	.lvb_bb2_notexitcond9_(bb_2_lvb_bb2_notexitcond9_),
	.lvb_bb2_mul3722_pop13_mul3722(bb_2_lvb_bb2_mul3722_pop13_mul3722),
	.lvb_bb2_notcmp1125_pop14_notcmp1125(bb_2_lvb_bb2_notcmp1125_pop14_notcmp1125),
	.lvb_bb2_notexitcond1428_pop15_notexitcond1428(bb_2_lvb_bb2_notexitcond1428_pop15_notexitcond1428),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_in_12(feedback_valid_12),
	.feedback_stall_out_12(feedback_stall_12),
	.feedback_data_in_12(feedback_data_12),
	.feedback_valid_in_10(feedback_valid_10),
	.feedback_stall_out_10(feedback_stall_10),
	.feedback_data_in_10(feedback_data_10),
	.feedback_stall_out_4(bb_2_feedback_stall_out_4),
	.feedback_valid_in_5(feedback_valid_5),
	.feedback_stall_out_5(feedback_stall_5),
	.feedback_data_in_5(feedback_data_5),
	.acl_pipelined_valid(bb_2_acl_pipelined_valid),
	.acl_pipelined_stall(bb_2_stall_out_0),
	.acl_pipelined_exiting_valid(bb_2_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_2_acl_pipelined_exiting_stall),
	.feedback_valid_in_11(feedback_valid_11),
	.feedback_stall_out_11(feedback_stall_11),
	.feedback_data_in_11(feedback_data_11),
	.feedback_valid_in_16(feedback_valid_16),
	.feedback_stall_out_16(feedback_stall_16),
	.feedback_data_in_16(feedback_data_16),
	.feedback_valid_in_13(feedback_valid_13),
	.feedback_stall_out_13(feedback_stall_13),
	.feedback_data_in_13(feedback_data_13),
	.feedback_valid_in_14(feedback_valid_14),
	.feedback_stall_out_14(feedback_stall_14),
	.feedback_data_in_14(feedback_data_14),
	.feedback_valid_in_15(feedback_valid_15),
	.feedback_stall_out_15(feedback_stall_15),
	.feedback_data_in_15(feedback_data_15),
	.feedback_valid_out_10(feedback_valid_10),
	.feedback_stall_in_10(feedback_stall_10),
	.feedback_data_out_10(feedback_data_10),
	.feedback_valid_out_5(feedback_valid_5),
	.feedback_stall_in_5(feedback_stall_5),
	.feedback_data_out_5(feedback_data_5),
	.feedback_valid_out_12(feedback_valid_12),
	.feedback_stall_in_12(feedback_stall_12),
	.feedback_data_out_12(feedback_data_12),
	.feedback_valid_out_16(feedback_valid_16),
	.feedback_stall_in_16(feedback_stall_16),
	.feedback_data_out_16(feedback_data_16),
	.feedback_valid_out_13(feedback_valid_13),
	.feedback_stall_in_13(feedback_stall_13),
	.feedback_data_out_13(feedback_data_13),
	.feedback_valid_out_14(feedback_valid_14),
	.feedback_stall_in_14(feedback_stall_14),
	.feedback_data_out_14(feedback_data_14),
	.feedback_valid_out_15(feedback_valid_15),
	.feedback_stall_in_15(feedback_stall_15),
	.feedback_data_out_15(feedback_data_15),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__burstcount),
	.local_bb2_ld__active(bb_2_local_bb2_ld__active),
	.clock2x(clock2x)
);


AOChalfSampleRobustImageKernel_basic_block_3 AOChalfSampleRobustImageKernel_basic_block_3 (
	.clock(clock),
	.resetn(resetn),
	.input_inSize_x(input_inSize_x),
	.input_r(input_r),
	.input_wii_div(bb_0_lvb_bb0_div),
	.input_wii_div1(bb_0_lvb_bb0_div1),
	.input_wii_cmp19(bb_0_lvb_bb0_cmp19),
	.input_wii_add7(bb_0_lvb_bb0_add7),
	.input_wii_sub20(bb_0_lvb_bb0_sub20),
	.input_wii_sub22(bb_0_lvb_bb0_sub22),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u12(bb_0_lvb_bb0_var__u0),
	.input_wii_var__u13(bb_0_lvb_bb0_var__u1),
	.input_wii_var__u14(bb_0_lvb_bb0_var__u2),
	.valid_in_0(bb_3_acl_pipelined_valid),
	.stall_out_0(bb_3_stall_out_0),
	.input_forked16_0(1'b0),
	.input_pixel_y_020_pop820_0('x),
	.input_mul3723_0('x),
	.input_notcmp1126_0('x),
	.input_notexitcond1429_0('x),
	.input_memdep_phi1_pop932_0('x),
	.input_mul534_0('x),
	.input_indvars_iv_pop1036_0('x),
	.input_var__u15_0('x),
	.input_memdep_phi1_or38_0('x),
	.input_var__u16_0('x),
	.input_notcmp40_0('x),
	.input_notexitcond942_0('x),
	.valid_in_1(loop_limiter_2_valid_out),
	.stall_out_1(bb_3_stall_out_1),
	.input_forked16_1(1'b1),
	.input_pixel_y_020_pop820_1(bb_2_lvb_bb2_pixel_y_020_pop819_pop12_pixel_y_020_pop819),
	.input_mul3723_1(bb_2_lvb_bb2_mul3722_pop13_mul3722),
	.input_notcmp1126_1(bb_2_lvb_bb2_notcmp1125_pop14_notcmp1125),
	.input_notexitcond1429_1(bb_2_lvb_bb2_notexitcond1428_pop15_notexitcond1428),
	.input_memdep_phi1_pop932_1(bb_2_lvb_bb2_memdep_phi1_pop931_pop16_memdep_phi1_pop931),
	.input_mul534_1(bb_2_lvb_bb2_mul5),
	.input_indvars_iv_pop1036_1(bb_2_lvb_bb2_indvars_iv_pop10_acl_pop_i64_0),
	.input_var__u15_1(bb_2_lvb_bb2_var_),
	.input_memdep_phi1_or38_1(bb_2_lvb_bb2_memdep_phi1_or),
	.input_var__u16_1(bb_2_lvb_bb2_ld_),
	.input_notcmp40_1(bb_2_lvb_bb2_notcmp),
	.input_notexitcond942_1(bb_2_lvb_bb2_notexitcond9_),
	.valid_out(bb_3_valid_out),
	.stall_in(loop_limiter_3_stall_out),
	.lvb_forked16(bb_3_lvb_forked16),
	.lvb_bb3_c0_exe1(bb_3_lvb_bb3_c0_exe1),
	.lvb_bb3_c0_exe2(bb_3_lvb_bb3_c0_exe2),
	.lvb_bb3_c0_exe3(bb_3_lvb_bb3_c0_exe3),
	.lvb_bb3_c0_exe4(bb_3_lvb_bb3_c0_exe4),
	.lvb_bb3_c0_exe5(bb_3_lvb_bb3_c0_exe5),
	.lvb_bb3_c0_exe6(bb_3_lvb_bb3_c0_exe6),
	.lvb_bb3_c0_exe7(bb_3_lvb_bb3_c0_exe7),
	.lvb_bb3_c0_exe8(bb_3_lvb_bb3_c0_exe8),
	.lvb_bb3_c0_exe9(bb_3_lvb_bb3_c0_exe9),
	.lvb_bb3_c0_exe10(bb_3_lvb_bb3_c0_exe10),
	.lvb_bb3_c0_exe11(bb_3_lvb_bb3_c0_exe11),
	.lvb_bb3_c0_exe12(bb_3_lvb_bb3_c0_exe12),
	.lvb_bb3_c0_exe13(bb_3_lvb_bb3_c0_exe13),
	.lvb_bb3_c0_exe14(bb_3_lvb_bb3_c0_exe14),
	.lvb_bb3_c0_exe15(bb_3_lvb_bb3_c0_exe15),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_in_17(feedback_valid_17),
	.feedback_stall_out_17(feedback_stall_17),
	.feedback_data_in_17(feedback_data_17),
	.feedback_valid_in_23(feedback_valid_23),
	.feedback_stall_out_23(feedback_stall_23),
	.feedback_data_in_23(feedback_data_23),
	.feedback_stall_out_2(bb_3_feedback_stall_out_2),
	.feedback_valid_in_3(feedback_valid_3),
	.feedback_stall_out_3(feedback_stall_3),
	.feedback_data_in_3(feedback_data_3),
	.acl_pipelined_valid(bb_3_acl_pipelined_valid),
	.acl_pipelined_stall(bb_3_stall_out_0),
	.acl_pipelined_exiting_valid(bb_3_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_3_acl_pipelined_exiting_stall),
	.feedback_valid_in_18(feedback_valid_18),
	.feedback_stall_out_18(feedback_stall_18),
	.feedback_data_in_18(feedback_data_18),
	.feedback_valid_in_19(feedback_valid_19),
	.feedback_stall_out_19(feedback_stall_19),
	.feedback_data_in_19(feedback_data_19),
	.feedback_valid_in_20(feedback_valid_20),
	.feedback_stall_out_20(feedback_stall_20),
	.feedback_data_in_20(feedback_data_20),
	.feedback_valid_in_21(feedback_valid_21),
	.feedback_stall_out_21(feedback_stall_21),
	.feedback_data_in_21(feedback_data_21),
	.feedback_valid_in_22(feedback_valid_22),
	.feedback_stall_out_22(feedback_stall_22),
	.feedback_data_in_22(feedback_data_22),
	.feedback_valid_in_24(feedback_valid_24),
	.feedback_stall_out_24(feedback_stall_24),
	.feedback_data_in_24(feedback_data_24),
	.feedback_valid_in_25(feedback_valid_25),
	.feedback_stall_out_25(feedback_stall_25),
	.feedback_data_in_25(feedback_data_25),
	.feedback_valid_in_26(feedback_valid_26),
	.feedback_stall_out_26(feedback_stall_26),
	.feedback_data_in_26(feedback_data_26),
	.feedback_valid_in_27(feedback_valid_27),
	.feedback_stall_out_27(feedback_stall_27),
	.feedback_data_in_27(feedback_data_27),
	.feedback_valid_in_28(feedback_valid_28),
	.feedback_stall_out_28(feedback_stall_28),
	.feedback_data_in_28(feedback_data_28),
	.feedback_valid_in_29(feedback_valid_29),
	.feedback_stall_out_29(feedback_stall_29),
	.feedback_data_in_29(feedback_data_29),
	.feedback_valid_out_3(feedback_valid_3),
	.feedback_stall_in_3(feedback_stall_3),
	.feedback_data_out_3(feedback_data_3),
	.feedback_valid_out_17(feedback_valid_17),
	.feedback_stall_in_17(feedback_stall_17),
	.feedback_data_out_17(feedback_data_17),
	.feedback_valid_out_23(feedback_valid_23),
	.feedback_stall_in_23(feedback_stall_23),
	.feedback_data_out_23(feedback_data_23),
	.feedback_valid_out_18(feedback_valid_18),
	.feedback_stall_in_18(feedback_stall_18),
	.feedback_data_out_18(feedback_data_18),
	.feedback_valid_out_19(feedback_valid_19),
	.feedback_stall_in_19(feedback_stall_19),
	.feedback_data_out_19(feedback_data_19),
	.feedback_valid_out_20(feedback_valid_20),
	.feedback_stall_in_20(feedback_stall_20),
	.feedback_data_out_20(feedback_data_20),
	.feedback_valid_out_21(feedback_valid_21),
	.feedback_stall_in_21(feedback_stall_21),
	.feedback_data_out_21(feedback_data_21),
	.feedback_valid_out_22(feedback_valid_22),
	.feedback_stall_in_22(feedback_stall_22),
	.feedback_data_out_22(feedback_data_22),
	.feedback_valid_out_24(feedback_valid_24),
	.feedback_stall_in_24(feedback_stall_24),
	.feedback_data_out_24(feedback_data_24),
	.feedback_valid_out_25(feedback_valid_25),
	.feedback_stall_in_25(feedback_stall_25),
	.feedback_data_out_25(feedback_data_25),
	.feedback_valid_out_26(feedback_valid_26),
	.feedback_stall_in_26(feedback_stall_26),
	.feedback_data_out_26(feedback_data_26),
	.feedback_valid_out_27(feedback_valid_27),
	.feedback_stall_in_27(feedback_stall_27),
	.feedback_data_out_27(feedback_data_27),
	.feedback_valid_out_28(feedback_valid_28),
	.feedback_stall_in_28(feedback_stall_28),
	.feedback_data_out_28(feedback_data_28),
	.feedback_valid_out_29(feedback_valid_29),
	.feedback_stall_in_29(feedback_stall_29),
	.feedback_data_out_29(feedback_data_29)
);


AOChalfSampleRobustImageKernel_basic_block_4 AOChalfSampleRobustImageKernel_basic_block_4 (
	.clock(clock),
	.resetn(resetn),
	.input_in(input_in),
	.input_r(input_r),
	.input_e_d(input_e_d),
	.input_wii_div(bb_0_lvb_bb0_div),
	.input_wii_div1(bb_0_lvb_bb0_div1),
	.input_wii_cmp19(bb_0_lvb_bb0_cmp19),
	.input_wii_add7(bb_0_lvb_bb0_add7),
	.input_wii_sub20(bb_0_lvb_bb0_sub20),
	.input_wii_sub22(bb_0_lvb_bb0_sub22),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u17(bb_0_lvb_bb0_var__u0),
	.input_wii_var__u18(bb_0_lvb_bb0_var__u1),
	.input_wii_var__u19(bb_0_lvb_bb0_var__u2),
	.valid_in_0(bb_4_acl_pipelined_valid),
	.stall_out_0(bb_4_stall_out_0),
	.input_forked_0(1'b0),
	.input_pixel_y_020_pop821_0('x),
	.input_mul3724_0('x),
	.input_notcmp1127_0('x),
	.input_notexitcond1430_0('x),
	.input_memdep_phi1_pop933_0('x),
	.input_mul535_0('x),
	.input_indvars_iv_pop1037_0('x),
	.input_var__u20_0('x),
	.input_memdep_phi1_or39_0('x),
	.input_var__u21_0('x),
	.input_notcmp41_0('x),
	.input_notexitcond943_0('x),
	.input_forked1644_0('x),
	.input_mul2445_0('x),
	.input_var__u22_0('x),
	.input_notexitcond546_0('x),
	.valid_in_1(loop_limiter_3_valid_out),
	.stall_out_1(bb_4_stall_out_1),
	.input_forked_1(1'b1),
	.input_pixel_y_020_pop821_1(bb_3_lvb_bb3_c0_exe5),
	.input_mul3724_1(bb_3_lvb_bb3_c0_exe6),
	.input_notcmp1127_1(bb_3_lvb_bb3_c0_exe7),
	.input_notexitcond1430_1(bb_3_lvb_bb3_c0_exe8),
	.input_memdep_phi1_pop933_1(bb_3_lvb_bb3_c0_exe9),
	.input_mul535_1(bb_3_lvb_bb3_c0_exe1),
	.input_indvars_iv_pop1037_1(bb_3_lvb_bb3_c0_exe10),
	.input_var__u20_1(bb_3_lvb_bb3_c0_exe11),
	.input_memdep_phi1_or39_1(bb_3_lvb_bb3_c0_exe12),
	.input_var__u21_1(bb_3_lvb_bb3_c0_exe13),
	.input_notcmp41_1(bb_3_lvb_bb3_c0_exe14),
	.input_notexitcond943_1(bb_3_lvb_bb3_c0_exe15),
	.input_forked1644_1(bb_3_lvb_forked16),
	.input_mul2445_1(bb_3_lvb_bb3_c0_exe2),
	.input_var__u22_1(bb_3_lvb_bb3_c0_exe3),
	.input_notexitcond546_1(bb_3_lvb_bb3_c0_exe4),
	.valid_out_0(bb_4_valid_out_0),
	.stall_in_0(bb_5_stall_out),
	.lvb_bb4_c0_exit87_c0_exi1386_0(bb_4_lvb_bb4_c0_exit87_c0_exi1386_0),
	.lvb_bb4_c0_exe794_0(bb_4_lvb_bb4_c0_exe794_0),
	.lvb_bb4_c0_exe895_0(bb_4_lvb_bb4_c0_exe895_0),
	.lvb_bb4_c0_exe996_0(bb_4_lvb_bb4_c0_exe996_0),
	.lvb_bb4_c0_exe1097_0(bb_4_lvb_bb4_c0_exe1097_0),
	.lvb_bb4_c0_exe1198_0(bb_4_lvb_bb4_c0_exe1198_0),
	.lvb_bb4_c0_exe1299_0(bb_4_lvb_bb4_c0_exe1299_0),
	.lvb_bb4_c1_exe1_0(bb_4_lvb_bb4_c1_exe1_0),
	.lvb_bb4_c1_exe2_0(bb_4_lvb_bb4_c1_exe2_0),
	.valid_out_1(bb_4_valid_out_1),
	.stall_in_1(1'b0),
	.lvb_bb4_c0_exit87_c0_exi1386_1(bb_4_lvb_bb4_c0_exit87_c0_exi1386_1),
	.lvb_bb4_c0_exe794_1(bb_4_lvb_bb4_c0_exe794_1),
	.lvb_bb4_c0_exe895_1(bb_4_lvb_bb4_c0_exe895_1),
	.lvb_bb4_c0_exe996_1(bb_4_lvb_bb4_c0_exe996_1),
	.lvb_bb4_c0_exe1097_1(bb_4_lvb_bb4_c0_exe1097_1),
	.lvb_bb4_c0_exe1198_1(bb_4_lvb_bb4_c0_exe1198_1),
	.lvb_bb4_c0_exe1299_1(bb_4_lvb_bb4_c0_exe1299_1),
	.lvb_bb4_c1_exe1_1(bb_4_lvb_bb4_c1_exe1_1),
	.lvb_bb4_c1_exe2_1(bb_4_lvb_bb4_c1_exe2_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_in_30(feedback_valid_30),
	.feedback_stall_out_30(feedback_stall_30),
	.feedback_data_in_30(feedback_data_30),
	.feedback_valid_in_40(feedback_valid_40),
	.feedback_stall_out_40(feedback_stall_40),
	.feedback_data_in_40(feedback_data_40),
	.feedback_stall_out_0(bb_4_feedback_stall_out_0),
	.feedback_valid_in_1(feedback_valid_1),
	.feedback_stall_out_1(feedback_stall_1),
	.feedback_data_in_1(feedback_data_1),
	.acl_pipelined_valid(bb_4_acl_pipelined_valid),
	.acl_pipelined_stall(bb_4_stall_out_0),
	.acl_pipelined_exiting_valid(bb_4_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_4_acl_pipelined_exiting_stall),
	.feedback_valid_in_46(feedback_valid_46),
	.feedback_stall_out_46(feedback_stall_46),
	.feedback_data_in_46(feedback_data_46),
	.feedback_valid_in_45(feedback_valid_45),
	.feedback_stall_out_45(feedback_stall_45),
	.feedback_data_in_45(feedback_data_45),
	.feedback_valid_in_41(feedback_valid_41),
	.feedback_stall_out_41(feedback_stall_41),
	.feedback_data_in_41(feedback_data_41),
	.feedback_valid_in_42(feedback_valid_42),
	.feedback_stall_out_42(feedback_stall_42),
	.feedback_data_in_42(feedback_data_42),
	.feedback_valid_in_33(feedback_valid_33),
	.feedback_stall_out_33(feedback_stall_33),
	.feedback_data_in_33(feedback_data_33),
	.feedback_valid_in_34(feedback_valid_34),
	.feedback_stall_out_34(feedback_stall_34),
	.feedback_data_in_34(feedback_data_34),
	.feedback_valid_in_35(feedback_valid_35),
	.feedback_stall_out_35(feedback_stall_35),
	.feedback_data_in_35(feedback_data_35),
	.feedback_valid_in_36(feedback_valid_36),
	.feedback_stall_out_36(feedback_stall_36),
	.feedback_data_in_36(feedback_data_36),
	.feedback_valid_in_37(feedback_valid_37),
	.feedback_stall_out_37(feedback_stall_37),
	.feedback_data_in_37(feedback_data_37),
	.feedback_valid_in_38(feedback_valid_38),
	.feedback_stall_out_38(feedback_stall_38),
	.feedback_data_in_38(feedback_data_38),
	.feedback_valid_in_39(feedback_valid_39),
	.feedback_stall_out_39(feedback_stall_39),
	.feedback_data_in_39(feedback_data_39),
	.feedback_valid_in_43(feedback_valid_43),
	.feedback_stall_out_43(feedback_stall_43),
	.feedback_data_in_43(feedback_data_43),
	.feedback_valid_in_44(feedback_valid_44),
	.feedback_stall_out_44(feedback_stall_44),
	.feedback_data_in_44(feedback_data_44),
	.feedback_valid_in_47(feedback_valid_47),
	.feedback_stall_out_47(feedback_stall_47),
	.feedback_data_in_47(feedback_data_47),
	.feedback_valid_out_1(feedback_valid_1),
	.feedback_stall_in_1(feedback_stall_1),
	.feedback_data_out_1(feedback_data_1),
	.feedback_valid_out_30(feedback_valid_30),
	.feedback_stall_in_30(feedback_stall_30),
	.feedback_data_out_30(feedback_data_30),
	.feedback_valid_out_45(feedback_valid_45),
	.feedback_stall_in_45(feedback_stall_45),
	.feedback_data_out_45(feedback_data_45),
	.feedback_valid_out_42(feedback_valid_42),
	.feedback_stall_in_42(feedback_stall_42),
	.feedback_data_out_42(feedback_data_42),
	.feedback_valid_out_41(feedback_valid_41),
	.feedback_stall_in_41(feedback_stall_41),
	.feedback_data_out_41(feedback_data_41),
	.feedback_valid_out_40(feedback_valid_40),
	.feedback_stall_in_40(feedback_stall_40),
	.feedback_data_out_40(feedback_data_40),
	.feedback_valid_out_33(feedback_valid_33),
	.feedback_stall_in_33(feedback_stall_33),
	.feedback_data_out_33(feedback_data_33),
	.feedback_valid_out_34(feedback_valid_34),
	.feedback_stall_in_34(feedback_stall_34),
	.feedback_data_out_34(feedback_data_34),
	.feedback_valid_out_35(feedback_valid_35),
	.feedback_stall_in_35(feedback_stall_35),
	.feedback_data_out_35(feedback_data_35),
	.feedback_valid_out_36(feedback_valid_36),
	.feedback_stall_in_36(feedback_stall_36),
	.feedback_data_out_36(feedback_data_36),
	.feedback_valid_out_37(feedback_valid_37),
	.feedback_stall_in_37(feedback_stall_37),
	.feedback_data_out_37(feedback_data_37),
	.feedback_valid_out_38(feedback_valid_38),
	.feedback_stall_in_38(feedback_stall_38),
	.feedback_data_out_38(feedback_data_38),
	.feedback_valid_out_39(feedback_valid_39),
	.feedback_stall_in_39(feedback_stall_39),
	.feedback_data_out_39(feedback_data_39),
	.feedback_valid_out_43(feedback_valid_43),
	.feedback_stall_in_43(feedback_stall_43),
	.feedback_data_out_43(feedback_data_43),
	.feedback_valid_out_44(feedback_valid_44),
	.feedback_stall_in_44(feedback_stall_44),
	.feedback_data_out_44(feedback_data_44),
	.feedback_valid_out_47(feedback_valid_47),
	.feedback_stall_in_47(feedback_stall_47),
	.feedback_data_out_47(feedback_data_47),
	.feedback_valid_out_46(feedback_valid_46),
	.feedback_stall_in_46(feedback_stall_46),
	.feedback_data_out_46(feedback_data_46),
	.avm_local_bb4_ld__readdata(avm_local_bb4_ld__readdata),
	.avm_local_bb4_ld__readdatavalid(avm_local_bb4_ld__readdatavalid),
	.avm_local_bb4_ld__waitrequest(avm_local_bb4_ld__waitrequest),
	.avm_local_bb4_ld__address(avm_local_bb4_ld__address),
	.avm_local_bb4_ld__read(avm_local_bb4_ld__read),
	.avm_local_bb4_ld__write(avm_local_bb4_ld__write),
	.avm_local_bb4_ld__writeack(avm_local_bb4_ld__writeack),
	.avm_local_bb4_ld__writedata(avm_local_bb4_ld__writedata),
	.avm_local_bb4_ld__byteenable(avm_local_bb4_ld__byteenable),
	.avm_local_bb4_ld__burstcount(avm_local_bb4_ld__burstcount),
	.local_bb4_ld__active(bb_4_local_bb4_ld__active),
	.clock2x(clock2x),
	.feedback_valid_in_48(feedback_valid_48),
	.feedback_stall_out_48(feedback_stall_48),
	.feedback_data_in_48(feedback_data_48),
	.feedback_valid_out_48(feedback_valid_48),
	.feedback_stall_in_48(feedback_stall_48),
	.feedback_data_out_48(feedback_data_48),
	.feedback_valid_in_31(feedback_valid_31),
	.feedback_stall_out_31(feedback_stall_31),
	.feedback_data_in_31(feedback_data_31),
	.feedback_valid_in_32(feedback_valid_32),
	.feedback_stall_out_32(feedback_stall_32),
	.feedback_data_in_32(feedback_data_32),
	.feedback_valid_out_32(feedback_valid_32),
	.feedback_stall_in_32(feedback_stall_32),
	.feedback_data_out_32(feedback_data_32),
	.feedback_valid_out_31(feedback_valid_31),
	.feedback_stall_in_31(feedback_stall_31),
	.feedback_data_out_31(feedback_data_31)
);


AOChalfSampleRobustImageKernel_basic_block_5 AOChalfSampleRobustImageKernel_basic_block_5 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_div(bb_0_lvb_bb0_div),
	.input_wii_div1(bb_0_lvb_bb0_div1),
	.input_wii_cmp19(bb_0_lvb_bb0_cmp19),
	.input_wii_add7(bb_0_lvb_bb0_add7),
	.input_wii_sub20(bb_0_lvb_bb0_sub20),
	.input_wii_sub22(bb_0_lvb_bb0_sub22),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u58(bb_0_lvb_bb0_var__u0),
	.input_wii_var__u59(bb_0_lvb_bb0_var__u1),
	.input_wii_var__u60(bb_0_lvb_bb0_var__u2),
	.valid_in(bb_4_valid_out_0),
	.stall_out(bb_5_stall_out),
	.input_c0_exit87_c0_exi1386(bb_4_lvb_bb4_c0_exit87_c0_exi1386_0),
	.input_c0_exe794(bb_4_lvb_bb4_c0_exe794_0),
	.input_c0_exe895(bb_4_lvb_bb4_c0_exe895_0),
	.input_c0_exe996(bb_4_lvb_bb4_c0_exe996_0),
	.input_c0_exe1097(bb_4_lvb_bb4_c0_exe1097_0),
	.input_c0_exe1198(bb_4_lvb_bb4_c0_exe1198_0),
	.input_c0_exe1299(bb_4_lvb_bb4_c0_exe1299_0),
	.input_c1_exe1(bb_4_lvb_bb4_c1_exe1_0),
	.input_c1_exe2(bb_4_lvb_bb4_c1_exe2_0),
	.valid_out_0(bb_5_valid_out_0),
	.stall_in_0(bb_6_stall_out),
	.lvb_c0_exe794_0(bb_5_lvb_c0_exe794_0),
	.lvb_c0_exe895_0(bb_5_lvb_c0_exe895_0),
	.lvb_c0_exe996_0(bb_5_lvb_c0_exe996_0),
	.lvb_c0_exe1097_0(bb_5_lvb_c0_exe1097_0),
	.lvb_c0_exe1198_0(bb_5_lvb_c0_exe1198_0),
	.lvb_c0_exe1299_0(bb_5_lvb_c0_exe1299_0),
	.lvb_c1_exe1_0(bb_5_lvb_c1_exe1_0),
	.lvb_c1_exe2_0(bb_5_lvb_c1_exe2_0),
	.valid_out_1(bb_5_valid_out_1),
	.stall_in_1(1'b0),
	.lvb_c0_exe794_1(bb_5_lvb_c0_exe794_1),
	.lvb_c0_exe895_1(bb_5_lvb_c0_exe895_1),
	.lvb_c0_exe996_1(bb_5_lvb_c0_exe996_1),
	.lvb_c0_exe1097_1(bb_5_lvb_c0_exe1097_1),
	.lvb_c0_exe1198_1(bb_5_lvb_c0_exe1198_1),
	.lvb_c0_exe1299_1(bb_5_lvb_c0_exe1299_1),
	.lvb_c1_exe1_1(bb_5_lvb_c1_exe1_1),
	.lvb_c1_exe2_1(bb_5_lvb_c1_exe2_1),
	.workgroup_size(workgroup_size),
	.start(start)
);


AOChalfSampleRobustImageKernel_basic_block_6 AOChalfSampleRobustImageKernel_basic_block_6 (
	.clock(clock),
	.resetn(resetn),
	.input_out(input_out),
	.input_wii_div(bb_0_lvb_bb0_div),
	.input_wii_div1(bb_0_lvb_bb0_div1),
	.input_wii_cmp19(bb_0_lvb_bb0_cmp19),
	.input_wii_add7(bb_0_lvb_bb0_add7),
	.input_wii_sub20(bb_0_lvb_bb0_sub20),
	.input_wii_sub22(bb_0_lvb_bb0_sub22),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u61(bb_0_lvb_bb0_var__u0),
	.input_wii_var__u62(bb_0_lvb_bb0_var__u1),
	.input_wii_var__u63(bb_0_lvb_bb0_var__u2),
	.valid_in(bb_5_valid_out_0),
	.stall_out(bb_6_stall_out),
	.input_c0_exe794(bb_5_lvb_c0_exe794_0),
	.input_c0_exe895(bb_5_lvb_c0_exe895_0),
	.input_c0_exe996(bb_5_lvb_c0_exe996_0),
	.input_c0_exe1097(bb_5_lvb_c0_exe1097_0),
	.input_c0_exe1198(bb_5_lvb_c0_exe1198_0),
	.input_c0_exe1299(bb_5_lvb_c0_exe1299_0),
	.input_c1_exe1(bb_5_lvb_c1_exe1_0),
	.input_c1_exe2(bb_5_lvb_c1_exe2_0),
	.valid_out_0(bb_6_valid_out_0),
	.stall_in_0(bb_7_stall_out),
	.lvb_c0_exe895_0(bb_6_lvb_c0_exe895_0),
	.lvb_c0_exe996_0(bb_6_lvb_c0_exe996_0),
	.lvb_bb6_st_c0_exe1108_0(bb_6_lvb_bb6_st_c0_exe1108_0),
	.valid_out_1(bb_6_valid_out_1),
	.stall_in_1(1'b0),
	.lvb_c0_exe895_1(bb_6_lvb_c0_exe895_1),
	.lvb_c0_exe996_1(bb_6_lvb_c0_exe996_1),
	.lvb_bb6_st_c0_exe1108_1(bb_6_lvb_bb6_st_c0_exe1108_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.avm_local_bb6_st_c0_exe1108_readdata(avm_local_bb6_st_c0_exe1108_readdata),
	.avm_local_bb6_st_c0_exe1108_readdatavalid(avm_local_bb6_st_c0_exe1108_readdatavalid),
	.avm_local_bb6_st_c0_exe1108_waitrequest(avm_local_bb6_st_c0_exe1108_waitrequest),
	.avm_local_bb6_st_c0_exe1108_address(avm_local_bb6_st_c0_exe1108_address),
	.avm_local_bb6_st_c0_exe1108_read(avm_local_bb6_st_c0_exe1108_read),
	.avm_local_bb6_st_c0_exe1108_write(avm_local_bb6_st_c0_exe1108_write),
	.avm_local_bb6_st_c0_exe1108_writeack(avm_local_bb6_st_c0_exe1108_writeack),
	.avm_local_bb6_st_c0_exe1108_writedata(avm_local_bb6_st_c0_exe1108_writedata),
	.avm_local_bb6_st_c0_exe1108_byteenable(avm_local_bb6_st_c0_exe1108_byteenable),
	.avm_local_bb6_st_c0_exe1108_burstcount(avm_local_bb6_st_c0_exe1108_burstcount),
	.local_bb6_st_c0_exe1108_active(bb_6_local_bb6_st_c0_exe1108_active),
	.clock2x(clock2x),
	.feedback_valid_out_11(feedback_valid_11),
	.feedback_stall_in_11(feedback_stall_11),
	.feedback_data_out_11(feedback_data_11)
);


AOChalfSampleRobustImageKernel_basic_block_7 AOChalfSampleRobustImageKernel_basic_block_7 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_div(bb_0_lvb_bb0_div),
	.input_wii_div1(bb_0_lvb_bb0_div1),
	.input_wii_cmp19(bb_0_lvb_bb0_cmp19),
	.input_wii_add7(bb_0_lvb_bb0_add7),
	.input_wii_sub20(bb_0_lvb_bb0_sub20),
	.input_wii_sub22(bb_0_lvb_bb0_sub22),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u64(bb_0_lvb_bb0_var__u0),
	.input_wii_var__u65(bb_0_lvb_bb0_var__u1),
	.input_wii_var__u66(bb_0_lvb_bb0_var__u2),
	.valid_in(bb_6_valid_out_0),
	.stall_out(bb_7_stall_out),
	.input_c0_exe895(bb_6_lvb_c0_exe895_0),
	.input_c0_exe996(bb_6_lvb_c0_exe996_0),
	.input_st_c0_exe1108(bb_6_lvb_bb6_st_c0_exe1108_0),
	.valid_out_0(bb_7_valid_out_0),
	.stall_in_0(bb_8_stall_out),
	.valid_out_1(bb_7_valid_out_1),
	.stall_in_1(1'b0),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_out_9(feedback_valid_9),
	.feedback_stall_in_9(feedback_stall_9),
	.feedback_data_out_9(feedback_data_9)
);


AOChalfSampleRobustImageKernel_basic_block_8 AOChalfSampleRobustImageKernel_basic_block_8 (
	.clock(clock),
	.resetn(resetn),
	.valid_in(bb_7_valid_out_0),
	.stall_out(bb_8_stall_out),
	.valid_out(bb_8_valid_out),
	.stall_in(stall_in),
	.workgroup_size(workgroup_size),
	.start(start)
);


acl_loop_limiter loop_limiter_1 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_1_valid_out),
	.i_stall(bb_2_stall_out_1),
	.i_valid_exit(bb_2_acl_pipelined_exiting_valid),
	.i_stall_exit(bb_2_acl_pipelined_exiting_stall),
	.o_valid(loop_limiter_1_valid_out),
	.o_stall(loop_limiter_1_stall_out)
);

defparam loop_limiter_1.ENTRY_WIDTH = 1;
defparam loop_limiter_1.EXIT_WIDTH = 1;
defparam loop_limiter_1.THRESHOLD = 2;

acl_loop_limiter loop_limiter_2 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_2_valid_out),
	.i_stall(bb_3_stall_out_1),
	.i_valid_exit(bb_3_acl_pipelined_exiting_valid),
	.i_stall_exit(bb_3_acl_pipelined_exiting_stall),
	.o_valid(loop_limiter_2_valid_out),
	.o_stall(loop_limiter_2_stall_out)
);

defparam loop_limiter_2.ENTRY_WIDTH = 1;
defparam loop_limiter_2.EXIT_WIDTH = 1;
defparam loop_limiter_2.THRESHOLD = 1;

acl_loop_limiter loop_limiter_3 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_3_valid_out),
	.i_stall(bb_4_stall_out_1),
	.i_valid_exit(bb_4_acl_pipelined_exiting_valid),
	.i_stall_exit(bb_4_acl_pipelined_exiting_stall),
	.o_valid(loop_limiter_3_valid_out),
	.o_stall(loop_limiter_3_stall_out)
);

defparam loop_limiter_3.ENTRY_WIDTH = 1;
defparam loop_limiter_3.EXIT_WIDTH = 1;
defparam loop_limiter_3.THRESHOLD = 1;

AOChalfSampleRobustImageKernel_sys_cycle_time system_cycle_time_module (
	.clock(clock),
	.resetn(resetn),
	.cur_cycle(cur_cycle)
);


assign workgroup_size = 32'h1;
assign valid_out = bb_8_valid_out;
assign stall_out = bb_0_stall_out;
assign writes_pending = bb_6_local_bb6_st_c0_exe1108_active;
assign lsus_active[0] = bb_2_local_bb2_ld__active;
assign lsus_active[1] = bb_4_local_bb4_ld__active;
assign lsus_active[2] = bb_6_local_bb6_st_c0_exe1108_active;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		has_a_write_pending <= 1'b0;
		has_a_lsu_active <= 1'b0;
	end
	else
	begin
		has_a_write_pending <= (|writes_pending);
		has_a_lsu_active <= (|lsus_active);
	end
end

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_function_wrapper
	(
		input 		clock,
		input 		resetn,
		input 		clock2x,
		input 		local_router_hang,
		input 		avs_cra_read,
		input 		avs_cra_write,
		input [4:0] 		avs_cra_address,
		input [63:0] 		avs_cra_writedata,
		input [7:0] 		avs_cra_byteenable,
		output reg [63:0] 		avs_cra_readdata,
		output reg 		avs_cra_readdatavalid,
		output 		cra_irq,
		input [511:0] 		avm_local_bb2_ld__inst0_readdata,
		input 		avm_local_bb2_ld__inst0_readdatavalid,
		input 		avm_local_bb2_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb2_ld__inst0_address,
		output 		avm_local_bb2_ld__inst0_read,
		output 		avm_local_bb2_ld__inst0_write,
		input 		avm_local_bb2_ld__inst0_writeack,
		output [511:0] 		avm_local_bb2_ld__inst0_writedata,
		output [63:0] 		avm_local_bb2_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb4_ld__inst0_readdata,
		input 		avm_local_bb4_ld__inst0_readdatavalid,
		input 		avm_local_bb4_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb4_ld__inst0_address,
		output 		avm_local_bb4_ld__inst0_read,
		output 		avm_local_bb4_ld__inst0_write,
		input 		avm_local_bb4_ld__inst0_writeack,
		output [511:0] 		avm_local_bb4_ld__inst0_writedata,
		output [63:0] 		avm_local_bb4_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb4_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb6_st_c0_exe1108_inst0_readdata,
		input 		avm_local_bb6_st_c0_exe1108_inst0_readdatavalid,
		input 		avm_local_bb6_st_c0_exe1108_inst0_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe1108_inst0_address,
		output 		avm_local_bb6_st_c0_exe1108_inst0_read,
		output 		avm_local_bb6_st_c0_exe1108_inst0_write,
		input 		avm_local_bb6_st_c0_exe1108_inst0_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe1108_inst0_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe1108_inst0_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe1108_inst0_burstcount
	);

// Responsible for interfacing a kernel with the outside world. It comprises a
// slave interface to specify the kernel arguments and retain kernel status. 

// This section of the wrapper implements the slave interface.
// twoXclock_consumer uses clock2x, even if nobody inside the kernel does. Keeps interface to acl_iface consistent for all kernels.
 reg start_NO_SHIFT_REG;
 reg started_NO_SHIFT_REG;
wire finish;
 reg [31:0] status_NO_SHIFT_REG;
wire has_a_write_pending;
wire has_a_lsu_active;
 reg [255:0] kernel_arguments_NO_SHIFT_REG;
 reg twoXclock_consumer_NO_SHIFT_REG /* synthesis  preserve  noprune  */;
 reg [31:0] workgroup_size_NO_SHIFT_REG;
 reg [31:0] global_size_NO_SHIFT_REG[2:0];
 reg [31:0] num_groups_NO_SHIFT_REG[2:0];
 reg [31:0] local_size_NO_SHIFT_REG[2:0];
 reg [31:0] work_dim_NO_SHIFT_REG;
 reg [31:0] global_offset_NO_SHIFT_REG[2:0];
 reg [63:0] profile_data_NO_SHIFT_REG;
 reg [31:0] profile_ctrl_NO_SHIFT_REG;
 reg [63:0] profile_start_cycle_NO_SHIFT_REG;
 reg [63:0] profile_stop_cycle_NO_SHIFT_REG;
wire dispatched_all_groups;
wire [31:0] group_id_tmp[2:0];
wire [31:0] global_id_base_out[2:0];
wire start_out;
wire [31:0] local_id[0:0][2:0];
wire [31:0] global_id[0:0][2:0];
wire [31:0] group_id[0:0][2:0];
wire iter_valid_in;
wire iter_stall_out;
wire stall_in;
wire stall_out;
wire valid_in;
wire valid_out;

always @(posedge clock2x or negedge resetn)
begin
	if (~(resetn))
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b1;
	end
end



// Work group dispatcher is responsible for issuing work-groups to id iterator(s)
acl_work_group_dispatcher group_dispatcher (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.num_groups(num_groups_NO_SHIFT_REG),
	.local_size(local_size_NO_SHIFT_REG),
	.stall_in(iter_stall_out),
	.valid_out(iter_valid_in),
	.group_id_out(group_id_tmp),
	.global_id_base_out(global_id_base_out),
	.start_out(start_out),
	.dispatched_all_groups(dispatched_all_groups)
);

defparam group_dispatcher.NUM_COPIES = 1;
defparam group_dispatcher.RUN_FOREVER = 0;


// This section of the wrapper implements an Avalon Slave Interface used to configure a kernel invocation.
// The few words words contain the status and the workgroup size registers.
// The remaining addressable space is reserved for kernel arguments.
 reg [63:0] cra_readdata_st1_NO_SHIFT_REG;
 reg [4:0] cra_addr_st1_NO_SHIFT_REG;
 reg cra_read_st1_NO_SHIFT_REG;
wire [63:0] bitenable;

assign bitenable[7:0] = (avs_cra_byteenable[0] ? 8'hFF : 8'h0);
assign bitenable[15:8] = (avs_cra_byteenable[1] ? 8'hFF : 8'h0);
assign bitenable[23:16] = (avs_cra_byteenable[2] ? 8'hFF : 8'h0);
assign bitenable[31:24] = (avs_cra_byteenable[3] ? 8'hFF : 8'h0);
assign bitenable[39:32] = (avs_cra_byteenable[4] ? 8'hFF : 8'h0);
assign bitenable[47:40] = (avs_cra_byteenable[5] ? 8'hFF : 8'h0);
assign bitenable[55:48] = (avs_cra_byteenable[6] ? 8'hFF : 8'h0);
assign bitenable[63:56] = (avs_cra_byteenable[7] ? 8'hFF : 8'h0);
assign cra_irq = (status_NO_SHIFT_REG[1] | status_NO_SHIFT_REG[3]);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		start_NO_SHIFT_REG <= 1'b0;
		started_NO_SHIFT_REG <= 1'b0;
		kernel_arguments_NO_SHIFT_REG <= 256'h0;
		status_NO_SHIFT_REG <= 32'h30000;
		profile_ctrl_NO_SHIFT_REG <= 32'h4;
		profile_start_cycle_NO_SHIFT_REG <= 64'h0;
		profile_stop_cycle_NO_SHIFT_REG <= 64'hFFFFFFFFFFFFFFFF;
		work_dim_NO_SHIFT_REG <= 32'h0;
		workgroup_size_NO_SHIFT_REG <= 32'h0;
		global_size_NO_SHIFT_REG[0] <= 32'h0;
		global_size_NO_SHIFT_REG[1] <= 32'h0;
		global_size_NO_SHIFT_REG[2] <= 32'h0;
		num_groups_NO_SHIFT_REG[0] <= 32'h0;
		num_groups_NO_SHIFT_REG[1] <= 32'h0;
		num_groups_NO_SHIFT_REG[2] <= 32'h0;
		local_size_NO_SHIFT_REG[0] <= 32'h0;
		local_size_NO_SHIFT_REG[1] <= 32'h0;
		local_size_NO_SHIFT_REG[2] <= 32'h0;
		global_offset_NO_SHIFT_REG[0] <= 32'h0;
		global_offset_NO_SHIFT_REG[1] <= 32'h0;
		global_offset_NO_SHIFT_REG[2] <= 32'h0;
	end
	else
	begin
		if (avs_cra_write)
		begin
			case (avs_cra_address)
				5'h0:
				begin
					status_NO_SHIFT_REG[31:16] <= 16'h3;
					status_NO_SHIFT_REG[15:0] <= ((status_NO_SHIFT_REG[15:0] & ~(bitenable[15:0])) | (avs_cra_writedata[15:0] & bitenable[15:0]));
				end

				5'h1:
				begin
					profile_ctrl_NO_SHIFT_REG <= ((profile_ctrl_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h3:
				begin
					profile_start_cycle_NO_SHIFT_REG[31:0] <= ((profile_start_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_start_cycle_NO_SHIFT_REG[63:32] <= ((profile_start_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h4:
				begin
					profile_stop_cycle_NO_SHIFT_REG[31:0] <= ((profile_stop_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_stop_cycle_NO_SHIFT_REG[63:32] <= ((profile_stop_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h5:
				begin
					work_dim_NO_SHIFT_REG <= ((work_dim_NO_SHIFT_REG & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					workgroup_size_NO_SHIFT_REG <= ((workgroup_size_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h6:
				begin
					global_size_NO_SHIFT_REG[0] <= ((global_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_size_NO_SHIFT_REG[1] <= ((global_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h7:
				begin
					global_size_NO_SHIFT_REG[2] <= ((global_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[0] <= ((num_groups_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h8:
				begin
					num_groups_NO_SHIFT_REG[1] <= ((num_groups_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[2] <= ((num_groups_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h9:
				begin
					local_size_NO_SHIFT_REG[0] <= ((local_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					local_size_NO_SHIFT_REG[1] <= ((local_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hA:
				begin
					local_size_NO_SHIFT_REG[2] <= ((local_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[0] <= ((global_offset_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hB:
				begin
					global_offset_NO_SHIFT_REG[1] <= ((global_offset_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[2] <= ((global_offset_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hC:
				begin
					kernel_arguments_NO_SHIFT_REG[31:0] <= ((kernel_arguments_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[63:32] <= ((kernel_arguments_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hD:
				begin
					kernel_arguments_NO_SHIFT_REG[95:64] <= ((kernel_arguments_NO_SHIFT_REG[95:64] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[127:96] <= ((kernel_arguments_NO_SHIFT_REG[127:96] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hE:
				begin
					kernel_arguments_NO_SHIFT_REG[159:128] <= ((kernel_arguments_NO_SHIFT_REG[159:128] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[191:160] <= ((kernel_arguments_NO_SHIFT_REG[191:160] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hF:
				begin
					kernel_arguments_NO_SHIFT_REG[223:192] <= ((kernel_arguments_NO_SHIFT_REG[223:192] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[255:224] <= ((kernel_arguments_NO_SHIFT_REG[255:224] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				default:
				begin
				end

			endcase
		end
		else
		begin
			if (status_NO_SHIFT_REG[0])
			begin
				start_NO_SHIFT_REG <= 1'b1;
			end
			if (start_NO_SHIFT_REG)
			begin
				status_NO_SHIFT_REG[0] <= 1'b0;
				started_NO_SHIFT_REG <= 1'b1;
			end
			if (started_NO_SHIFT_REG)
			begin
				start_NO_SHIFT_REG <= 1'b0;
			end
			if (finish)
			begin
				status_NO_SHIFT_REG[1] <= 1'b1;
				started_NO_SHIFT_REG <= 1'b0;
			end
		end
		status_NO_SHIFT_REG[11] <= 1'b0;
		status_NO_SHIFT_REG[12] <= (|has_a_lsu_active);
		status_NO_SHIFT_REG[13] <= (|has_a_write_pending);
		status_NO_SHIFT_REG[14] <= (|valid_in);
		status_NO_SHIFT_REG[15] <= started_NO_SHIFT_REG;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cra_read_st1_NO_SHIFT_REG <= 1'b0;
		cra_addr_st1_NO_SHIFT_REG <= 5'h0;
		cra_readdata_st1_NO_SHIFT_REG <= 64'h0;
	end
	else
	begin
		cra_read_st1_NO_SHIFT_REG <= avs_cra_read;
		cra_addr_st1_NO_SHIFT_REG <= avs_cra_address;
		case (avs_cra_address)
			5'h0:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= status_NO_SHIFT_REG;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			5'h1:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= 'x;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			5'h2:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			5'h3:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			5'h4:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			default:
			begin
				cra_readdata_st1_NO_SHIFT_REG <= status_NO_SHIFT_REG;
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		avs_cra_readdatavalid <= 1'b0;
		avs_cra_readdata <= 64'h0;
	end
	else
	begin
		avs_cra_readdatavalid <= cra_read_st1_NO_SHIFT_REG;
		case (cra_addr_st1_NO_SHIFT_REG)
			5'h2:
			begin
				avs_cra_readdata[63:0] <= profile_data_NO_SHIFT_REG;
			end

			default:
			begin
				avs_cra_readdata <= cra_readdata_st1_NO_SHIFT_REG;
			end

		endcase
	end
end


// Handshaking signals used to control data through the pipeline

// Determine when the kernel is finished.
acl_kernel_finish_detector kernel_finish_detector (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.wg_size(workgroup_size_NO_SHIFT_REG),
	.wg_dispatch_valid_out(iter_valid_in),
	.wg_dispatch_stall_in(iter_stall_out),
	.dispatched_all_groups(dispatched_all_groups),
	.kernel_copy_valid_out(valid_out),
	.kernel_copy_stall_in(stall_in),
	.pending_writes(has_a_write_pending),
	.finish(finish)
);

defparam kernel_finish_detector.TESSELLATION_SIZE = 0;
defparam kernel_finish_detector.NUM_COPIES = 1;
defparam kernel_finish_detector.WG_SIZE_W = 32;

assign stall_in = 1'b0;

// Creating ID iterator and kernel instance for every requested kernel copy

// ID iterator is responsible for iterating over all local ids for given work-groups
acl_id_iterator id_iter_inst0 (
	.clock(clock),
	.resetn(resetn),
	.start(start_out),
	.valid_in(iter_valid_in),
	.stall_out(iter_stall_out),
	.stall_in(stall_out),
	.valid_out(valid_in),
	.group_id_in(group_id_tmp),
	.global_id_base_in(global_id_base_out),
	.local_size(local_size_NO_SHIFT_REG),
	.global_size(global_size_NO_SHIFT_REG),
	.local_id(local_id[0]),
	.global_id(global_id[0]),
	.group_id(group_id[0])
);



// This section instantiates a kernel function block
AOChalfSampleRobustImageKernel_function AOChalfSampleRobustImageKernel_function_inst0 (
	.clock(clock),
	.resetn(resetn),
	.stall_out(stall_out),
	.valid_in(valid_in),
	.valid_out(valid_out),
	.stall_in(stall_in),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__inst0_readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__inst0_readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__inst0_waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__inst0_address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__inst0_read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__inst0_write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__inst0_writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__inst0_writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__inst0_byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__inst0_burstcount),
	.avm_local_bb4_ld__readdata(avm_local_bb4_ld__inst0_readdata),
	.avm_local_bb4_ld__readdatavalid(avm_local_bb4_ld__inst0_readdatavalid),
	.avm_local_bb4_ld__waitrequest(avm_local_bb4_ld__inst0_waitrequest),
	.avm_local_bb4_ld__address(avm_local_bb4_ld__inst0_address),
	.avm_local_bb4_ld__read(avm_local_bb4_ld__inst0_read),
	.avm_local_bb4_ld__write(avm_local_bb4_ld__inst0_write),
	.avm_local_bb4_ld__writeack(avm_local_bb4_ld__inst0_writeack),
	.avm_local_bb4_ld__writedata(avm_local_bb4_ld__inst0_writedata),
	.avm_local_bb4_ld__byteenable(avm_local_bb4_ld__inst0_byteenable),
	.avm_local_bb4_ld__burstcount(avm_local_bb4_ld__inst0_burstcount),
	.avm_local_bb6_st_c0_exe1108_readdata(avm_local_bb6_st_c0_exe1108_inst0_readdata),
	.avm_local_bb6_st_c0_exe1108_readdatavalid(avm_local_bb6_st_c0_exe1108_inst0_readdatavalid),
	.avm_local_bb6_st_c0_exe1108_waitrequest(avm_local_bb6_st_c0_exe1108_inst0_waitrequest),
	.avm_local_bb6_st_c0_exe1108_address(avm_local_bb6_st_c0_exe1108_inst0_address),
	.avm_local_bb6_st_c0_exe1108_read(avm_local_bb6_st_c0_exe1108_inst0_read),
	.avm_local_bb6_st_c0_exe1108_write(avm_local_bb6_st_c0_exe1108_inst0_write),
	.avm_local_bb6_st_c0_exe1108_writeack(avm_local_bb6_st_c0_exe1108_inst0_writeack),
	.avm_local_bb6_st_c0_exe1108_writedata(avm_local_bb6_st_c0_exe1108_inst0_writedata),
	.avm_local_bb6_st_c0_exe1108_byteenable(avm_local_bb6_st_c0_exe1108_inst0_byteenable),
	.avm_local_bb6_st_c0_exe1108_burstcount(avm_local_bb6_st_c0_exe1108_inst0_burstcount),
	.start(start_out),
	.input_inSize_x(kernel_arguments_NO_SHIFT_REG[159:128]),
	.input_inSize_y(kernel_arguments_NO_SHIFT_REG[191:160]),
	.input_r(kernel_arguments_NO_SHIFT_REG[255:224]),
	.clock2x(clock2x),
	.input_in(kernel_arguments_NO_SHIFT_REG[127:64]),
	.input_e_d(kernel_arguments_NO_SHIFT_REG[223:192]),
	.input_out(kernel_arguments_NO_SHIFT_REG[63:0]),
	.has_a_write_pending(has_a_write_pending),
	.has_a_lsu_active(has_a_lsu_active)
);



endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOChalfSampleRobustImageKernel_sys_cycle_time
	(
		input 		clock,
		input 		resetn,
		output [31:0] 		cur_cycle
	);


 reg [31:0] cur_count_NO_SHIFT_REG;

assign cur_cycle = cur_count_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cur_count_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		cur_count_NO_SHIFT_REG <= (cur_count_NO_SHIFT_REG + 32'h1);
	end
end

endmodule

