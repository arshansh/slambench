// (C) 1992-2015 Altera Corporation. All rights reserved.                         
// Your use of Altera Corporation's design tools, logic functions and other       
// software and tools, and its AMPP partner logic functions, and any output       
// files any of the foregoing (including device programming or simulation         
// files), and any associated documentation or information are expressly subject  
// to the terms and conditions of the Altera Program License Subscription         
// Agreement, Altera MegaCore Function License Agreement, or other applicable     
// license agreement, including, without limitation, that your use is for the     
// sole purpose of programming logic devices manufactured by Altera and sold by   
// Altera or its authorized distributors.  Please refer to the applicable         
// agreement for further details.                                                 
    

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_0
	(
		input 		clock,
		input 		resetn,
		input 		start,
		input [31:0] 		input_r,
		input [31:0] 		input_global_size_0,
		input [31:0] 		input_global_size_1,
		input [31:0] 		input_e_d,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out,
		input 		stall_in,
		output 		lvb_bb0_cmp1526,
		output [31:0] 		lvb_bb0_sub24,
		output [31:0] 		lvb_bb0_sub27,
		output [31:0] 		lvb_bb0_mul48,
		output [63:0] 		lvb_bb0_var_,
		output [63:0] 		lvb_bb0_var__u0,
		input [31:0] 		workgroup_size
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub_inputs_ready;
 reg local_bb0_sub_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub_valid_out_0_NO_SHIFT_REG;
wire local_bb0_sub_stall_in_0;
 reg local_bb0_sub_valid_out_1_NO_SHIFT_REG;
wire local_bb0_sub_stall_in_1;
wire local_bb0_sub_output_regs_ready;
 reg [31:0] local_bb0_sub_NO_SHIFT_REG;
wire local_bb0_sub_causedstall;

assign local_bb0_sub_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb0_sub_output_regs_ready = (~(local_bb0_sub_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_sub_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_sub_stall_in_0)) & (~(local_bb0_sub_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_sub_stall_in_1))));
assign merge_node_stall_in_0 = (~(local_bb0_sub_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub_output_regs_ready) | ~(local_bb0_sub_inputs_ready)));
assign local_bb0_sub_causedstall = (local_bb0_sub_inputs_ready && (~(local_bb0_sub_output_regs_ready) && !(~(local_bb0_sub_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub_NO_SHIFT_REG <= 'x;
		local_bb0_sub_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_sub_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub_NO_SHIFT_REG <= 'x;
			local_bb0_sub_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_sub_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub_output_regs_ready)
			begin
				local_bb0_sub_NO_SHIFT_REG <= (32'h0 - input_r);
				local_bb0_sub_valid_out_0_NO_SHIFT_REG <= local_bb0_sub_inputs_ready;
				local_bb0_sub_valid_out_1_NO_SHIFT_REG <= local_bb0_sub_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub_stall_in_0))
				begin
					local_bb0_sub_valid_out_0_NO_SHIFT_REG <= local_bb0_sub_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_sub_stall_in_1))
				begin
					local_bb0_sub_valid_out_1_NO_SHIFT_REG <= local_bb0_sub_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub_inputs_ready)
			begin
				local_bb0_sub_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub24_inputs_ready;
 reg local_bb0_sub24_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub24_valid_out_NO_SHIFT_REG;
wire local_bb0_sub24_stall_in;
wire local_bb0_sub24_output_regs_ready;
 reg [31:0] local_bb0_sub24_NO_SHIFT_REG;
wire local_bb0_sub24_causedstall;

assign local_bb0_sub24_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign local_bb0_sub24_output_regs_ready = (~(local_bb0_sub24_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_sub24_valid_out_NO_SHIFT_REG) | ~(local_bb0_sub24_stall_in))));
assign merge_node_stall_in_2 = (~(local_bb0_sub24_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub24_output_regs_ready) | ~(local_bb0_sub24_inputs_ready)));
assign local_bb0_sub24_causedstall = (local_bb0_sub24_inputs_ready && (~(local_bb0_sub24_output_regs_ready) && !(~(local_bb0_sub24_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub24_NO_SHIFT_REG <= 'x;
		local_bb0_sub24_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub24_NO_SHIFT_REG <= 'x;
			local_bb0_sub24_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub24_output_regs_ready)
			begin
				local_bb0_sub24_NO_SHIFT_REG <= (input_global_size_0 + 32'hFFFFFFFF);
				local_bb0_sub24_valid_out_NO_SHIFT_REG <= local_bb0_sub24_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub24_stall_in))
				begin
					local_bb0_sub24_valid_out_NO_SHIFT_REG <= local_bb0_sub24_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub24_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub24_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub24_inputs_ready)
			begin
				local_bb0_sub24_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_sub27_inputs_ready;
 reg local_bb0_sub27_wii_reg_NO_SHIFT_REG;
 reg local_bb0_sub27_valid_out_NO_SHIFT_REG;
wire local_bb0_sub27_stall_in;
wire local_bb0_sub27_output_regs_ready;
 reg [31:0] local_bb0_sub27_NO_SHIFT_REG;
wire local_bb0_sub27_causedstall;

assign local_bb0_sub27_inputs_ready = merge_node_valid_out_3_NO_SHIFT_REG;
assign local_bb0_sub27_output_regs_ready = (~(local_bb0_sub27_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_sub27_valid_out_NO_SHIFT_REG) | ~(local_bb0_sub27_stall_in))));
assign merge_node_stall_in_3 = (~(local_bb0_sub27_wii_reg_NO_SHIFT_REG) & (~(local_bb0_sub27_output_regs_ready) | ~(local_bb0_sub27_inputs_ready)));
assign local_bb0_sub27_causedstall = (local_bb0_sub27_inputs_ready && (~(local_bb0_sub27_output_regs_ready) && !(~(local_bb0_sub27_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub27_NO_SHIFT_REG <= 'x;
		local_bb0_sub27_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub27_NO_SHIFT_REG <= 'x;
			local_bb0_sub27_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub27_output_regs_ready)
			begin
				local_bb0_sub27_NO_SHIFT_REG <= (input_global_size_1 + 32'hFFFFFFFF);
				local_bb0_sub27_valid_out_NO_SHIFT_REG <= local_bb0_sub27_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_sub27_stall_in))
				begin
					local_bb0_sub27_valid_out_NO_SHIFT_REG <= local_bb0_sub27_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_sub27_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_sub27_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_sub27_inputs_ready)
			begin
				local_bb0_sub27_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u1_inputs_ready;
 reg local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u1_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u1_stall_in;
wire local_bb0_var__u1_output_regs_ready;
 reg [31:0] local_bb0_var__u1_NO_SHIFT_REG;
wire local_bb0_var__u1_causedstall;

assign local_bb0_var__u1_inputs_ready = merge_node_valid_out_4_NO_SHIFT_REG;
assign local_bb0_var__u1_output_regs_ready = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u1_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u1_stall_in))));
assign merge_node_stall_in_4 = (~(local_bb0_var__u1_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u1_output_regs_ready) | ~(local_bb0_var__u1_inputs_ready)));
assign local_bb0_var__u1_causedstall = (local_bb0_var__u1_inputs_ready && (~(local_bb0_var__u1_output_regs_ready) && !(~(local_bb0_var__u1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_NO_SHIFT_REG <= 'x;
		local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_NO_SHIFT_REG <= 'x;
			local_bb0_var__u1_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_output_regs_ready)
			begin
				local_bb0_var__u1_NO_SHIFT_REG <= input_e_d;
				local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u1_stall_in))
				begin
					local_bb0_var__u1_valid_out_NO_SHIFT_REG <= local_bb0_var__u1_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u1_inputs_ready)
			begin
				local_bb0_var__u1_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__u0_inputs_ready;
 reg local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__u0_valid_out_NO_SHIFT_REG;
wire local_bb0_var__u0_stall_in;
wire local_bb0_var__u0_output_regs_ready;
 reg [63:0] local_bb0_var__u0_NO_SHIFT_REG;
wire local_bb0_var__u0_causedstall;

assign local_bb0_var__u0_inputs_ready = merge_node_valid_out_6_NO_SHIFT_REG;
assign local_bb0_var__u0_output_regs_ready = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__u0_valid_out_NO_SHIFT_REG) | ~(local_bb0_var__u0_stall_in))));
assign merge_node_stall_in_6 = (~(local_bb0_var__u0_wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__u0_output_regs_ready) | ~(local_bb0_var__u0_inputs_ready)));
assign local_bb0_var__u0_causedstall = (local_bb0_var__u0_inputs_ready && (~(local_bb0_var__u0_output_regs_ready) && !(~(local_bb0_var__u0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_NO_SHIFT_REG <= 'x;
		local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_NO_SHIFT_REG <= 'x;
			local_bb0_var__u0_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_output_regs_ready)
			begin
				local_bb0_var__u0_NO_SHIFT_REG <= $signed(input_r);
				local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__u0_stall_in))
				begin
					local_bb0_var__u0_valid_out_NO_SHIFT_REG <= local_bb0_var__u0_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__u0_inputs_ready)
			begin
				local_bb0_var__u0_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp1526_inputs_ready;
 reg local_bb0_cmp1526_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp1526_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp1526_stall_in;
wire local_bb0_cmp1526_output_regs_ready;
 reg local_bb0_cmp1526_NO_SHIFT_REG;
wire local_bb0_cmp1526_causedstall;

assign local_bb0_cmp1526_inputs_ready = (local_bb0_sub_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign local_bb0_cmp1526_output_regs_ready = (~(local_bb0_cmp1526_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp1526_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp1526_stall_in))));
assign local_bb0_sub_stall_in_0 = (~(local_bb0_cmp1526_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp1526_output_regs_ready) | ~(local_bb0_cmp1526_inputs_ready)));
assign merge_node_stall_in_1 = (~(local_bb0_cmp1526_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp1526_output_regs_ready) | ~(local_bb0_cmp1526_inputs_ready)));
assign local_bb0_cmp1526_causedstall = (local_bb0_cmp1526_inputs_ready && (~(local_bb0_cmp1526_output_regs_ready) && !(~(local_bb0_cmp1526_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp1526_NO_SHIFT_REG <= 'x;
		local_bb0_cmp1526_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp1526_NO_SHIFT_REG <= 'x;
			local_bb0_cmp1526_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp1526_output_regs_ready)
			begin
				local_bb0_cmp1526_NO_SHIFT_REG <= ($signed(local_bb0_sub_NO_SHIFT_REG) > $signed(input_r));
				local_bb0_cmp1526_valid_out_NO_SHIFT_REG <= local_bb0_cmp1526_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp1526_stall_in))
				begin
					local_bb0_cmp1526_valid_out_NO_SHIFT_REG <= local_bb0_cmp1526_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp1526_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp1526_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp1526_inputs_ready)
			begin
				local_bb0_cmp1526_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_var__inputs_ready;
 reg local_bb0_var__wii_reg_NO_SHIFT_REG;
 reg local_bb0_var__valid_out_NO_SHIFT_REG;
wire local_bb0_var__stall_in;
wire local_bb0_var__output_regs_ready;
 reg [63:0] local_bb0_var__NO_SHIFT_REG;
wire local_bb0_var__causedstall;

assign local_bb0_var__inputs_ready = local_bb0_sub_valid_out_1_NO_SHIFT_REG;
assign local_bb0_var__output_regs_ready = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_var__valid_out_NO_SHIFT_REG) | ~(local_bb0_var__stall_in))));
assign local_bb0_sub_stall_in_1 = (~(local_bb0_var__wii_reg_NO_SHIFT_REG) & (~(local_bb0_var__output_regs_ready) | ~(local_bb0_var__inputs_ready)));
assign local_bb0_var__causedstall = (local_bb0_var__inputs_ready && (~(local_bb0_var__output_regs_ready) && !(~(local_bb0_var__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__NO_SHIFT_REG <= 'x;
		local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__NO_SHIFT_REG <= 'x;
			local_bb0_var__valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__output_regs_ready)
			begin
				local_bb0_var__NO_SHIFT_REG <= $signed(local_bb0_sub_NO_SHIFT_REG);
				local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__inputs_ready;
			end
			else
			begin
				if (~(local_bb0_var__stall_in))
				begin
					local_bb0_var__valid_out_NO_SHIFT_REG <= local_bb0_var__wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_var__inputs_ready)
			begin
				local_bb0_var__wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_2to2_bb0_var__u1_valid_out_0;
wire rstag_2to2_bb0_var__u1_stall_in_0;
wire rstag_2to2_bb0_var__u1_valid_out_1;
wire rstag_2to2_bb0_var__u1_stall_in_1;
wire rstag_2to2_bb0_var__u1_valid_out_2;
wire rstag_2to2_bb0_var__u1_stall_in_2;
wire rstag_2to2_bb0_var__u1_inputs_ready;
wire rstag_2to2_bb0_var__u1_stall_local;
 reg rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG;
wire rstag_2to2_bb0_var__u1_combined_valid;
 reg [31:0] rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_2to2_bb0_var__u1;
 reg rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG;
 reg rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG;
 reg rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG;

assign rstag_2to2_bb0_var__u1_inputs_ready = local_bb0_var__u1_valid_out_NO_SHIFT_REG;
assign rstag_2to2_bb0_var__u1 = (rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG ? rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG : local_bb0_var__u1_NO_SHIFT_REG);
assign rstag_2to2_bb0_var__u1_combined_valid = (rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG | rstag_2to2_bb0_var__u1_inputs_ready);
assign rstag_2to2_bb0_var__u1_stall_local = ((rstag_2to2_bb0_var__u1_stall_in_0 & ~(rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG)) | (rstag_2to2_bb0_var__u1_stall_in_1 & ~(rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG)) | (rstag_2to2_bb0_var__u1_stall_in_2 & ~(rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG)));
assign rstag_2to2_bb0_var__u1_valid_out_0 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG));
assign rstag_2to2_bb0_var__u1_valid_out_1 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG));
assign rstag_2to2_bb0_var__u1_valid_out_2 = (rstag_2to2_bb0_var__u1_combined_valid & ~(rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG));
assign local_bb0_var__u1_stall_in = (|rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_2to2_bb0_var__u1_stall_local)
			begin
				if (~(rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG))
				begin
					rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= rstag_2to2_bb0_var__u1_inputs_ready;
				end
			end
			else
			begin
				rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_2to2_bb0_var__u1_staging_valid_NO_SHIFT_REG))
		begin
			rstag_2to2_bb0_var__u1_staging_reg_NO_SHIFT_REG <= local_bb0_var__u1_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_0_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_0)) & rstag_2to2_bb0_var__u1_stall_local);
			rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_1_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_1)) & rstag_2to2_bb0_var__u1_stall_local);
			rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1_combined_valid & (rstag_2to2_bb0_var__u1_consumed_2_NO_SHIFT_REG | ~(rstag_2to2_bb0_var__u1_stall_in_2)) & rstag_2to2_bb0_var__u1_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and33_i_inputs_ready;
 reg local_bb0_and33_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and33_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and33_i_stall_in;
wire local_bb0_and33_i_output_regs_ready;
 reg [31:0] local_bb0_and33_i_NO_SHIFT_REG;
wire local_bb0_and33_i_causedstall;

assign local_bb0_and33_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_0;
assign local_bb0_and33_i_output_regs_ready = (~(local_bb0_and33_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and33_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and33_i_stall_in))));
assign rstag_2to2_bb0_var__u1_stall_in_0 = (~(local_bb0_and33_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and33_i_output_regs_ready) | ~(local_bb0_and33_i_inputs_ready)));
assign local_bb0_and33_i_causedstall = (local_bb0_and33_i_inputs_ready && (~(local_bb0_and33_i_output_regs_ready) && !(~(local_bb0_and33_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and33_i_NO_SHIFT_REG <= 'x;
		local_bb0_and33_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and33_i_NO_SHIFT_REG <= 'x;
			local_bb0_and33_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and33_i_output_regs_ready)
			begin
				local_bb0_and33_i_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1 & 32'h807FFFFF);
				local_bb0_and33_i_valid_out_NO_SHIFT_REG <= local_bb0_and33_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and33_i_stall_in))
				begin
					local_bb0_and33_i_valid_out_NO_SHIFT_REG <= local_bb0_and33_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and33_i_inputs_ready)
			begin
				local_bb0_and33_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_and2_i_valid_out;
wire local_bb0_and2_i_stall_in;
wire local_bb0_and2_i_inputs_ready;
wire local_bb0_and2_i_stall_local;
wire [31:0] local_bb0_and2_i;

assign local_bb0_and2_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_1;
assign local_bb0_and2_i = (rstag_2to2_bb0_var__u1 & 32'h7FFFFF);
assign local_bb0_and2_i_valid_out = local_bb0_and2_i_inputs_ready;
assign local_bb0_and2_i_stall_local = local_bb0_and2_i_stall_in;
assign rstag_2to2_bb0_var__u1_stall_in_1 = (|local_bb0_and2_i_stall_local);

// This section implements a registered operation.
// 
wire local_bb0_shr_i_inputs_ready;
 reg local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_shr_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_shr_i_stall_in_0;
 reg local_bb0_shr_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_shr_i_stall_in_1;
wire local_bb0_shr_i_output_regs_ready;
 reg [31:0] local_bb0_shr_i_NO_SHIFT_REG;
wire local_bb0_shr_i_causedstall;

assign local_bb0_shr_i_inputs_ready = rstag_2to2_bb0_var__u1_valid_out_2;
assign local_bb0_shr_i_output_regs_ready = (~(local_bb0_shr_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_shr_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_shr_i_stall_in_0)) & (~(local_bb0_shr_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_shr_i_stall_in_1))));
assign rstag_2to2_bb0_var__u1_stall_in_2 = (~(local_bb0_shr_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_shr_i_output_regs_ready) | ~(local_bb0_shr_i_inputs_ready)));
assign local_bb0_shr_i_causedstall = (local_bb0_shr_i_inputs_ready && (~(local_bb0_shr_i_output_regs_ready) && !(~(local_bb0_shr_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_shr_i_NO_SHIFT_REG <= 'x;
		local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_shr_i_NO_SHIFT_REG <= 'x;
			local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_shr_i_output_regs_ready)
			begin
				local_bb0_shr_i_NO_SHIFT_REG <= (rstag_2to2_bb0_var__u1 >> 32'h17);
				local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= local_bb0_shr_i_inputs_ready;
				local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= local_bb0_shr_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_shr_i_stall_in_0))
				begin
					local_bb0_shr_i_valid_out_0_NO_SHIFT_REG <= local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_shr_i_stall_in_1))
				begin
					local_bb0_shr_i_valid_out_1_NO_SHIFT_REG <= local_bb0_shr_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_shr_i_inputs_ready)
			begin
				local_bb0_shr_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_lnot6_i_inputs_ready;
 reg local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_lnot6_i_valid_out_NO_SHIFT_REG;
wire local_bb0_lnot6_i_stall_in;
wire local_bb0_lnot6_i_output_regs_ready;
 reg local_bb0_lnot6_i_NO_SHIFT_REG;
wire local_bb0_lnot6_i_causedstall;

assign local_bb0_lnot6_i_inputs_ready = local_bb0_and2_i_valid_out;
assign local_bb0_lnot6_i_output_regs_ready = (~(local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_lnot6_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_lnot6_i_stall_in))));
assign local_bb0_and2_i_stall_in = (~(local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_lnot6_i_output_regs_ready) | ~(local_bb0_lnot6_i_inputs_ready)));
assign local_bb0_lnot6_i_causedstall = (local_bb0_lnot6_i_inputs_ready && (~(local_bb0_lnot6_i_output_regs_ready) && !(~(local_bb0_lnot6_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_lnot6_i_NO_SHIFT_REG <= 'x;
		local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_lnot6_i_NO_SHIFT_REG <= 'x;
			local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_lnot6_i_output_regs_ready)
			begin
				local_bb0_lnot6_i_NO_SHIFT_REG <= ((local_bb0_and2_i & 32'h7FFFFF) != 32'h0);
				local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= local_bb0_lnot6_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_lnot6_i_stall_in))
				begin
					local_bb0_lnot6_i_valid_out_NO_SHIFT_REG <= local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_lnot6_i_inputs_ready)
			begin
				local_bb0_lnot6_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and1_i_inputs_ready;
 reg local_bb0_and1_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and1_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and1_i_stall_in;
wire local_bb0_and1_i_output_regs_ready;
 reg [31:0] local_bb0_and1_i_NO_SHIFT_REG;
wire local_bb0_and1_i_causedstall;

assign local_bb0_and1_i_inputs_ready = local_bb0_shr_i_valid_out_0_NO_SHIFT_REG;
assign local_bb0_and1_i_output_regs_ready = (~(local_bb0_and1_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and1_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and1_i_stall_in))));
assign local_bb0_shr_i_stall_in_0 = (~(local_bb0_and1_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and1_i_output_regs_ready) | ~(local_bb0_and1_i_inputs_ready)));
assign local_bb0_and1_i_causedstall = (local_bb0_and1_i_inputs_ready && (~(local_bb0_and1_i_output_regs_ready) && !(~(local_bb0_and1_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and1_i_NO_SHIFT_REG <= 'x;
		local_bb0_and1_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and1_i_NO_SHIFT_REG <= 'x;
			local_bb0_and1_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and1_i_output_regs_ready)
			begin
				local_bb0_and1_i_NO_SHIFT_REG <= ((local_bb0_shr_i_NO_SHIFT_REG & 32'h1FF) & 32'hFF);
				local_bb0_and1_i_valid_out_NO_SHIFT_REG <= local_bb0_and1_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and1_i_stall_in))
				begin
					local_bb0_and1_i_valid_out_NO_SHIFT_REG <= local_bb0_and1_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and1_i_inputs_ready)
			begin
				local_bb0_and1_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_4to4_bb0_and1_i_valid_out_0;
wire rstag_4to4_bb0_and1_i_stall_in_0;
wire rstag_4to4_bb0_and1_i_valid_out_1;
wire rstag_4to4_bb0_and1_i_stall_in_1;
wire rstag_4to4_bb0_and1_i_valid_out_2;
wire rstag_4to4_bb0_and1_i_stall_in_2;
wire rstag_4to4_bb0_and1_i_inputs_ready;
wire rstag_4to4_bb0_and1_i_stall_local;
 reg rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG;
wire rstag_4to4_bb0_and1_i_combined_valid;
 reg [31:0] rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_4to4_bb0_and1_i;
 reg rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG;
 reg rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG;
 reg rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG;

assign rstag_4to4_bb0_and1_i_inputs_ready = local_bb0_and1_i_valid_out_NO_SHIFT_REG;
assign rstag_4to4_bb0_and1_i = (rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG ? rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG : (local_bb0_and1_i_NO_SHIFT_REG & 32'hFF));
assign rstag_4to4_bb0_and1_i_combined_valid = (rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG | rstag_4to4_bb0_and1_i_inputs_ready);
assign rstag_4to4_bb0_and1_i_stall_local = ((rstag_4to4_bb0_and1_i_stall_in_0 & ~(rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG)) | (rstag_4to4_bb0_and1_i_stall_in_1 & ~(rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG)) | (rstag_4to4_bb0_and1_i_stall_in_2 & ~(rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG)));
assign rstag_4to4_bb0_and1_i_valid_out_0 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG));
assign rstag_4to4_bb0_and1_i_valid_out_1 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG));
assign rstag_4to4_bb0_and1_i_valid_out_2 = (rstag_4to4_bb0_and1_i_combined_valid & ~(rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG));
assign local_bb0_and1_i_stall_in = (|rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_4to4_bb0_and1_i_stall_local)
			begin
				if (~(rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= rstag_4to4_bb0_and1_i_inputs_ready;
				end
			end
			else
			begin
				rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_4to4_bb0_and1_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_4to4_bb0_and1_i_staging_reg_NO_SHIFT_REG <= (local_bb0_and1_i_NO_SHIFT_REG & 32'hFF);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_0_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_0)) & rstag_4to4_bb0_and1_i_stall_local);
			rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_1_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_1)) & rstag_4to4_bb0_and1_i_stall_local);
			rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG <= (rstag_4to4_bb0_and1_i_combined_valid & (rstag_4to4_bb0_and1_i_consumed_2_NO_SHIFT_REG | ~(rstag_4to4_bb0_and1_i_stall_in_2)) & rstag_4to4_bb0_and1_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp10_i_inputs_ready;
 reg local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_cmp10_i_stall_in_0;
 reg local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_cmp10_i_stall_in_1;
wire local_bb0_cmp10_i_output_regs_ready;
 reg local_bb0_cmp10_i_NO_SHIFT_REG;
wire local_bb0_cmp10_i_causedstall;

assign local_bb0_cmp10_i_inputs_ready = rstag_4to4_bb0_and1_i_valid_out_1;
assign local_bb0_cmp10_i_output_regs_ready = (~(local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_cmp10_i_stall_in_0)) & (~(local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_cmp10_i_stall_in_1))));
assign rstag_4to4_bb0_and1_i_stall_in_1 = (~(local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp10_i_output_regs_ready) | ~(local_bb0_cmp10_i_inputs_ready)));
assign local_bb0_cmp10_i_causedstall = (local_bb0_cmp10_i_inputs_ready && (~(local_bb0_cmp10_i_output_regs_ready) && !(~(local_bb0_cmp10_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp10_i_NO_SHIFT_REG <= 'x;
		local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp10_i_NO_SHIFT_REG <= 'x;
			local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp10_i_output_regs_ready)
			begin
				local_bb0_cmp10_i_NO_SHIFT_REG <= ((rstag_4to4_bb0_and1_i & 32'hFF) == 32'h0);
				local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp10_i_inputs_ready;
				local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp10_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp10_i_stall_in_0))
				begin
					local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_cmp10_i_stall_in_1))
				begin
					local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp10_i_inputs_ready)
			begin
				local_bb0_cmp10_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp_i_inputs_ready;
 reg local_bb0_cmp_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp_i_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp_i_stall_in;
wire local_bb0_cmp_i_output_regs_ready;
 reg local_bb0_cmp_i_NO_SHIFT_REG;
wire local_bb0_cmp_i_causedstall;

assign local_bb0_cmp_i_inputs_ready = rstag_4to4_bb0_and1_i_valid_out_2;
assign local_bb0_cmp_i_output_regs_ready = (~(local_bb0_cmp_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp_i_stall_in))));
assign rstag_4to4_bb0_and1_i_stall_in_2 = (~(local_bb0_cmp_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp_i_output_regs_ready) | ~(local_bb0_cmp_i_inputs_ready)));
assign local_bb0_cmp_i_causedstall = (local_bb0_cmp_i_inputs_ready && (~(local_bb0_cmp_i_output_regs_ready) && !(~(local_bb0_cmp_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp_i_NO_SHIFT_REG <= 'x;
		local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp_i_NO_SHIFT_REG <= 'x;
			local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp_i_output_regs_ready)
			begin
				local_bb0_cmp_i_NO_SHIFT_REG <= ((rstag_4to4_bb0_and1_i & 32'hFF) == 32'hFF);
				local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= local_bb0_cmp_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp_i_stall_in))
				begin
					local_bb0_cmp_i_valid_out_NO_SHIFT_REG <= local_bb0_cmp_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp_i_inputs_ready)
			begin
				local_bb0_cmp_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_not_cmp10_i_valid_out;
wire local_bb0_not_cmp10_i_stall_in;
wire local_bb0_not_cmp10_i_inputs_ready;
wire local_bb0_not_cmp10_i_stall_local;
wire local_bb0_not_cmp10_i;

assign local_bb0_not_cmp10_i_inputs_ready = local_bb0_cmp10_i_valid_out_1_NO_SHIFT_REG;
assign local_bb0_not_cmp10_i = (local_bb0_cmp10_i_NO_SHIFT_REG ^ 1'b1);
assign local_bb0_not_cmp10_i_valid_out = local_bb0_not_cmp10_i_inputs_ready;
assign local_bb0_not_cmp10_i_stall_local = local_bb0_not_cmp10_i_stall_in;
assign local_bb0_cmp10_i_stall_in_1 = (|local_bb0_not_cmp10_i_stall_local);

// This section implements a staging register.
// 
wire rstag_5to5_bb0_cmp_i_valid_out_0;
wire rstag_5to5_bb0_cmp_i_stall_in_0;
wire rstag_5to5_bb0_cmp_i_valid_out_1;
wire rstag_5to5_bb0_cmp_i_stall_in_1;
wire rstag_5to5_bb0_cmp_i_valid_out_2;
wire rstag_5to5_bb0_cmp_i_stall_in_2;
wire rstag_5to5_bb0_cmp_i_valid_out_3;
wire rstag_5to5_bb0_cmp_i_stall_in_3;
wire rstag_5to5_bb0_cmp_i_inputs_ready;
wire rstag_5to5_bb0_cmp_i_stall_local;
 reg rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb0_cmp_i_combined_valid;
 reg rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG;
wire rstag_5to5_bb0_cmp_i;
 reg rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG;
 reg rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG;

assign rstag_5to5_bb0_cmp_i_inputs_ready = local_bb0_cmp_i_valid_out_NO_SHIFT_REG;
assign rstag_5to5_bb0_cmp_i = (rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG : local_bb0_cmp_i_NO_SHIFT_REG);
assign rstag_5to5_bb0_cmp_i_combined_valid = (rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG | rstag_5to5_bb0_cmp_i_inputs_ready);
assign rstag_5to5_bb0_cmp_i_stall_local = ((rstag_5to5_bb0_cmp_i_stall_in_0 & ~(rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_1 & ~(rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_2 & ~(rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG)) | (rstag_5to5_bb0_cmp_i_stall_in_3 & ~(rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG)));
assign rstag_5to5_bb0_cmp_i_valid_out_0 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_1 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_2 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG));
assign rstag_5to5_bb0_cmp_i_valid_out_3 = (rstag_5to5_bb0_cmp_i_combined_valid & ~(rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG));
assign local_bb0_cmp_i_stall_in = (|rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_5to5_bb0_cmp_i_stall_local)
			begin
				if (~(rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb0_cmp_i_inputs_ready;
				end
			end
			else
			begin
				rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_5to5_bb0_cmp_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb0_cmp_i_staging_reg_NO_SHIFT_REG <= local_bb0_cmp_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= 1'b0;
			rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_0_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_0)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_1_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_1)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_2_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_2)) & rstag_5to5_bb0_cmp_i_stall_local);
			rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i_combined_valid & (rstag_5to5_bb0_cmp_i_consumed_3_NO_SHIFT_REG | ~(rstag_5to5_bb0_cmp_i_stall_in_3)) & rstag_5to5_bb0_cmp_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_conv22_i_inputs_ready;
 reg local_bb0_conv22_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_conv22_i_valid_out_NO_SHIFT_REG;
wire local_bb0_conv22_i_stall_in;
wire local_bb0_conv22_i_output_regs_ready;
 reg [31:0] local_bb0_conv22_i_NO_SHIFT_REG;
wire local_bb0_conv22_i_causedstall;

assign local_bb0_conv22_i_inputs_ready = rstag_5to5_bb0_cmp_i_valid_out_0;
assign local_bb0_conv22_i_output_regs_ready = (~(local_bb0_conv22_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_conv22_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_conv22_i_stall_in))));
assign rstag_5to5_bb0_cmp_i_stall_in_0 = (~(local_bb0_conv22_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_conv22_i_output_regs_ready) | ~(local_bb0_conv22_i_inputs_ready)));
assign local_bb0_conv22_i_causedstall = (local_bb0_conv22_i_inputs_ready && (~(local_bb0_conv22_i_output_regs_ready) && !(~(local_bb0_conv22_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_conv22_i_NO_SHIFT_REG <= 'x;
		local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_conv22_i_NO_SHIFT_REG <= 'x;
			local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_conv22_i_output_regs_ready)
			begin
				local_bb0_conv22_i_NO_SHIFT_REG <= rstag_5to5_bb0_cmp_i;
				local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= local_bb0_conv22_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_conv22_i_stall_in))
				begin
					local_bb0_conv22_i_valid_out_NO_SHIFT_REG <= local_bb0_conv22_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_conv22_i_inputs_ready)
			begin
				local_bb0_conv22_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__7_i_inputs_ready;
 reg local_bb0__7_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__7_i_valid_out_NO_SHIFT_REG;
wire local_bb0__7_i_stall_in;
wire local_bb0__7_i_output_regs_ready;
 reg local_bb0__7_i_NO_SHIFT_REG;
wire local_bb0__7_i_causedstall;

assign local_bb0__7_i_inputs_ready = (local_bb0_not_cmp10_i_valid_out & rstag_5to5_bb0_cmp_i_valid_out_1);
assign local_bb0__7_i_output_regs_ready = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__7_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__7_i_stall_in))));
assign local_bb0_not_cmp10_i_stall_in = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__7_i_output_regs_ready) | ~(local_bb0__7_i_inputs_ready)));
assign rstag_5to5_bb0_cmp_i_stall_in_1 = (~(local_bb0__7_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__7_i_output_regs_ready) | ~(local_bb0__7_i_inputs_ready)));
assign local_bb0__7_i_causedstall = (local_bb0__7_i_inputs_ready && (~(local_bb0__7_i_output_regs_ready) && !(~(local_bb0__7_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__7_i_NO_SHIFT_REG <= 'x;
		local_bb0__7_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__7_i_NO_SHIFT_REG <= 'x;
			local_bb0__7_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__7_i_output_regs_ready)
			begin
				local_bb0__7_i_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i | local_bb0_not_cmp10_i);
				local_bb0__7_i_valid_out_NO_SHIFT_REG <= local_bb0__7_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__7_i_stall_in))
				begin
					local_bb0__7_i_valid_out_NO_SHIFT_REG <= local_bb0__7_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__7_i_inputs_ready)
			begin
				local_bb0__7_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_not_cmp_i_valid_out;
wire local_bb0_not_cmp_i_stall_in;
wire local_bb0_not_cmp_i_inputs_ready;
wire local_bb0_not_cmp_i_stall_local;
wire local_bb0_not_cmp_i;

assign local_bb0_not_cmp_i_inputs_ready = rstag_5to5_bb0_cmp_i_valid_out_2;
assign local_bb0_not_cmp_i = (rstag_5to5_bb0_cmp_i ^ 1'b1);
assign local_bb0_not_cmp_i_valid_out = local_bb0_not_cmp_i_inputs_ready;
assign local_bb0_not_cmp_i_stall_local = local_bb0_not_cmp_i_stall_in;
assign rstag_5to5_bb0_cmp_i_stall_in_2 = (|local_bb0_not_cmp_i_stall_local);

// This section implements a registered operation.
// 
wire local_bb0___i_inputs_ready;
 reg local_bb0___i_wii_reg_NO_SHIFT_REG;
 reg local_bb0___i_valid_out_0_NO_SHIFT_REG;
wire local_bb0___i_stall_in_0;
 reg local_bb0___i_valid_out_1_NO_SHIFT_REG;
wire local_bb0___i_stall_in_1;
wire local_bb0___i_output_regs_ready;
 reg local_bb0___i_NO_SHIFT_REG;
wire local_bb0___i_causedstall;

assign local_bb0___i_inputs_ready = (local_bb0_lnot6_i_valid_out_NO_SHIFT_REG & rstag_5to5_bb0_cmp_i_valid_out_3);
assign local_bb0___i_output_regs_ready = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0___i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0___i_stall_in_0)) & (~(local_bb0___i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0___i_stall_in_1))));
assign local_bb0_lnot6_i_stall_in = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & (~(local_bb0___i_output_regs_ready) | ~(local_bb0___i_inputs_ready)));
assign rstag_5to5_bb0_cmp_i_stall_in_3 = (~(local_bb0___i_wii_reg_NO_SHIFT_REG) & (~(local_bb0___i_output_regs_ready) | ~(local_bb0___i_inputs_ready)));
assign local_bb0___i_causedstall = (local_bb0___i_inputs_ready && (~(local_bb0___i_output_regs_ready) && !(~(local_bb0___i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0___i_NO_SHIFT_REG <= 'x;
		local_bb0___i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0___i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0___i_NO_SHIFT_REG <= 'x;
			local_bb0___i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0___i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0___i_output_regs_ready)
			begin
				local_bb0___i_NO_SHIFT_REG <= (rstag_5to5_bb0_cmp_i & local_bb0_lnot6_i_NO_SHIFT_REG);
				local_bb0___i_valid_out_0_NO_SHIFT_REG <= local_bb0___i_inputs_ready;
				local_bb0___i_valid_out_1_NO_SHIFT_REG <= local_bb0___i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0___i_stall_in_0))
				begin
					local_bb0___i_valid_out_0_NO_SHIFT_REG <= local_bb0___i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0___i_stall_in_1))
				begin
					local_bb0___i_valid_out_1_NO_SHIFT_REG <= local_bb0___i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0___i_inputs_ready)
			begin
				local_bb0___i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_6to6_bb0__7_i_valid_out_0;
wire rstag_6to6_bb0__7_i_stall_in_0;
wire rstag_6to6_bb0__7_i_valid_out_1;
wire rstag_6to6_bb0__7_i_stall_in_1;
wire rstag_6to6_bb0__7_i_inputs_ready;
wire rstag_6to6_bb0__7_i_stall_local;
 reg rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG;
wire rstag_6to6_bb0__7_i_combined_valid;
 reg rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG;
wire rstag_6to6_bb0__7_i;
 reg rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG;
 reg rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG;

assign rstag_6to6_bb0__7_i_inputs_ready = local_bb0__7_i_valid_out_NO_SHIFT_REG;
assign rstag_6to6_bb0__7_i = (rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG ? rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG : local_bb0__7_i_NO_SHIFT_REG);
assign rstag_6to6_bb0__7_i_combined_valid = (rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG | rstag_6to6_bb0__7_i_inputs_ready);
assign rstag_6to6_bb0__7_i_stall_local = ((rstag_6to6_bb0__7_i_stall_in_0 & ~(rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG)) | (rstag_6to6_bb0__7_i_stall_in_1 & ~(rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG)));
assign rstag_6to6_bb0__7_i_valid_out_0 = (rstag_6to6_bb0__7_i_combined_valid & ~(rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG));
assign rstag_6to6_bb0__7_i_valid_out_1 = (rstag_6to6_bb0__7_i_combined_valid & ~(rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__7_i_stall_in = (|rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_6to6_bb0__7_i_stall_local)
			begin
				if (~(rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= rstag_6to6_bb0__7_i_inputs_ready;
				end
			end
			else
			begin
				rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_6to6_bb0__7_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_6to6_bb0__7_i_staging_reg_NO_SHIFT_REG <= local_bb0__7_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG <= (rstag_6to6_bb0__7_i_combined_valid & (rstag_6to6_bb0__7_i_consumed_0_NO_SHIFT_REG | ~(rstag_6to6_bb0__7_i_stall_in_0)) & rstag_6to6_bb0__7_i_stall_local);
			rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG <= (rstag_6to6_bb0__7_i_combined_valid & (rstag_6to6_bb0__7_i_consumed_1_NO_SHIFT_REG | ~(rstag_6to6_bb0__7_i_stall_in_1)) & rstag_6to6_bb0__7_i_stall_local);
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__4_i_inputs_ready;
 reg local_bb0__4_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__4_i_valid_out_NO_SHIFT_REG;
wire local_bb0__4_i_stall_in;
wire local_bb0__4_i_output_regs_ready;
 reg local_bb0__4_i_NO_SHIFT_REG;
wire local_bb0__4_i_causedstall;

assign local_bb0__4_i_inputs_ready = (local_bb0_cmp10_i_valid_out_0_NO_SHIFT_REG & local_bb0_not_cmp_i_valid_out);
assign local_bb0__4_i_output_regs_ready = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__4_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__4_i_stall_in))));
assign local_bb0_cmp10_i_stall_in_0 = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__4_i_output_regs_ready) | ~(local_bb0__4_i_inputs_ready)));
assign local_bb0_not_cmp_i_stall_in = (~(local_bb0__4_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__4_i_output_regs_ready) | ~(local_bb0__4_i_inputs_ready)));
assign local_bb0__4_i_causedstall = (local_bb0__4_i_inputs_ready && (~(local_bb0__4_i_output_regs_ready) && !(~(local_bb0__4_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__4_i_NO_SHIFT_REG <= 'x;
		local_bb0__4_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__4_i_NO_SHIFT_REG <= 'x;
			local_bb0__4_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__4_i_output_regs_ready)
			begin
				local_bb0__4_i_NO_SHIFT_REG <= (local_bb0_cmp10_i_NO_SHIFT_REG & local_bb0_not_cmp_i);
				local_bb0__4_i_valid_out_NO_SHIFT_REG <= local_bb0__4_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__4_i_stall_in))
				begin
					local_bb0__4_i_valid_out_NO_SHIFT_REG <= local_bb0__4_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__4_i_inputs_ready)
			begin
				local_bb0__4_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_conv44_i_stall_local;
wire [31:0] local_bb0_conv44_i;

assign local_bb0_conv44_i[31:1] = 31'h0;
assign local_bb0_conv44_i[0] = local_bb0___i_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb0_cond50_i_stall_local;
wire [31:0] local_bb0_cond50_i;

assign local_bb0_cond50_i = (local_bb0___i_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements a registered operation.
// 
wire local_bb0__12_i_inputs_ready;
 reg local_bb0__12_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__12_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0__12_i_stall_in_0;
 reg local_bb0__12_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0__12_i_stall_in_1;
wire local_bb0__12_i_output_regs_ready;
 reg local_bb0__12_i_NO_SHIFT_REG;
wire local_bb0__12_i_causedstall;

assign local_bb0__12_i_inputs_ready = rstag_6to6_bb0__7_i_valid_out_0;
assign local_bb0__12_i_output_regs_ready = (~(local_bb0__12_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0__12_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0__12_i_stall_in_0)) & (~(local_bb0__12_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0__12_i_stall_in_1))));
assign rstag_6to6_bb0__7_i_stall_in_0 = (~(local_bb0__12_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__12_i_output_regs_ready) | ~(local_bb0__12_i_inputs_ready)));
assign local_bb0__12_i_causedstall = (local_bb0__12_i_inputs_ready && (~(local_bb0__12_i_output_regs_ready) && !(~(local_bb0__12_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__12_i_NO_SHIFT_REG <= 'x;
		local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__12_i_NO_SHIFT_REG <= 'x;
			local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__12_i_output_regs_ready)
			begin
				local_bb0__12_i_NO_SHIFT_REG <= (1'b0 & rstag_6to6_bb0__7_i);
				local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= local_bb0__12_i_inputs_ready;
				local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= local_bb0__12_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__12_i_stall_in_0))
				begin
					local_bb0__12_i_valid_out_0_NO_SHIFT_REG <= local_bb0__12_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0__12_i_stall_in_1))
				begin
					local_bb0__12_i_valid_out_1_NO_SHIFT_REG <= local_bb0__12_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__12_i_inputs_ready)
			begin
				local_bb0__12_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__8_i_inputs_ready;
 reg local_bb0__8_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__8_i_valid_out_NO_SHIFT_REG;
wire local_bb0__8_i_stall_in;
wire local_bb0__8_i_output_regs_ready;
 reg local_bb0__8_i_NO_SHIFT_REG;
wire local_bb0__8_i_causedstall;

assign local_bb0__8_i_inputs_ready = rstag_6to6_bb0__7_i_valid_out_1;
assign local_bb0__8_i_output_regs_ready = (~(local_bb0__8_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__8_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__8_i_stall_in))));
assign rstag_6to6_bb0__7_i_stall_in_1 = (~(local_bb0__8_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__8_i_output_regs_ready) | ~(local_bb0__8_i_inputs_ready)));
assign local_bb0__8_i_causedstall = (local_bb0__8_i_inputs_ready && (~(local_bb0__8_i_output_regs_ready) && !(~(local_bb0__8_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__8_i_NO_SHIFT_REG <= 'x;
		local_bb0__8_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__8_i_NO_SHIFT_REG <= 'x;
			local_bb0__8_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__8_i_output_regs_ready)
			begin
				local_bb0__8_i_NO_SHIFT_REG <= (1'b1 & rstag_6to6_bb0__7_i);
				local_bb0__8_i_valid_out_NO_SHIFT_REG <= local_bb0__8_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__8_i_stall_in))
				begin
					local_bb0__8_i_valid_out_NO_SHIFT_REG <= local_bb0__8_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__8_i_inputs_ready)
			begin
				local_bb0__8_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_7to7_bb0__4_i_valid_out_0;
wire rstag_7to7_bb0__4_i_stall_in_0;
wire rstag_7to7_bb0__4_i_valid_out_1;
wire rstag_7to7_bb0__4_i_stall_in_1;
wire rstag_7to7_bb0__4_i_inputs_ready;
wire rstag_7to7_bb0__4_i_stall_local;
 reg rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG;
wire rstag_7to7_bb0__4_i_combined_valid;
 reg rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG;
wire rstag_7to7_bb0__4_i;
 reg rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG;
 reg rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG;

assign rstag_7to7_bb0__4_i_inputs_ready = local_bb0__4_i_valid_out_NO_SHIFT_REG;
assign rstag_7to7_bb0__4_i = (rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG ? rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG : local_bb0__4_i_NO_SHIFT_REG);
assign rstag_7to7_bb0__4_i_combined_valid = (rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG | rstag_7to7_bb0__4_i_inputs_ready);
assign rstag_7to7_bb0__4_i_stall_local = ((rstag_7to7_bb0__4_i_stall_in_0 & ~(rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG)) | (rstag_7to7_bb0__4_i_stall_in_1 & ~(rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG)));
assign rstag_7to7_bb0__4_i_valid_out_0 = (rstag_7to7_bb0__4_i_combined_valid & ~(rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG));
assign rstag_7to7_bb0__4_i_valid_out_1 = (rstag_7to7_bb0__4_i_combined_valid & ~(rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__4_i_stall_in = (|rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_7to7_bb0__4_i_stall_local)
			begin
				if (~(rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= rstag_7to7_bb0__4_i_inputs_ready;
				end
			end
			else
			begin
				rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_7to7_bb0__4_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_7to7_bb0__4_i_staging_reg_NO_SHIFT_REG <= local_bb0__4_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG <= (rstag_7to7_bb0__4_i_combined_valid & (rstag_7to7_bb0__4_i_consumed_0_NO_SHIFT_REG | ~(rstag_7to7_bb0__4_i_stall_in_0)) & rstag_7to7_bb0__4_i_stall_local);
			rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG <= (rstag_7to7_bb0__4_i_combined_valid & (rstag_7to7_bb0__4_i_consumed_1_NO_SHIFT_REG | ~(rstag_7to7_bb0__4_i_stall_in_1)) & rstag_7to7_bb0__4_i_stall_local);
		end
	end
end


// This section implements a staging register.
// 
wire rstag_7to7_bb0__8_i_valid_out_0;
wire rstag_7to7_bb0__8_i_stall_in_0;
wire rstag_7to7_bb0__8_i_valid_out_1;
wire rstag_7to7_bb0__8_i_stall_in_1;
wire rstag_7to7_bb0__8_i_inputs_ready;
wire rstag_7to7_bb0__8_i_stall_local;
 reg rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG;
wire rstag_7to7_bb0__8_i_combined_valid;
 reg rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG;
wire rstag_7to7_bb0__8_i;
 reg rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG;
 reg rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG;

assign rstag_7to7_bb0__8_i_inputs_ready = local_bb0__8_i_valid_out_NO_SHIFT_REG;
assign rstag_7to7_bb0__8_i = (rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG ? rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG : local_bb0__8_i_NO_SHIFT_REG);
assign rstag_7to7_bb0__8_i_combined_valid = (rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG | rstag_7to7_bb0__8_i_inputs_ready);
assign rstag_7to7_bb0__8_i_stall_local = ((rstag_7to7_bb0__8_i_stall_in_0 & ~(rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG)) | (rstag_7to7_bb0__8_i_stall_in_1 & ~(rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG)));
assign rstag_7to7_bb0__8_i_valid_out_0 = (rstag_7to7_bb0__8_i_combined_valid & ~(rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG));
assign rstag_7to7_bb0__8_i_valid_out_1 = (rstag_7to7_bb0__8_i_combined_valid & ~(rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__8_i_stall_in = (|rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_7to7_bb0__8_i_stall_local)
			begin
				if (~(rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= rstag_7to7_bb0__8_i_inputs_ready;
				end
			end
			else
			begin
				rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_7to7_bb0__8_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_7to7_bb0__8_i_staging_reg_NO_SHIFT_REG <= local_bb0__8_i_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i_combined_valid & (rstag_7to7_bb0__8_i_consumed_0_NO_SHIFT_REG | ~(rstag_7to7_bb0__8_i_stall_in_0)) & rstag_7to7_bb0__8_i_stall_local);
			rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i_combined_valid & (rstag_7to7_bb0__8_i_consumed_1_NO_SHIFT_REG | ~(rstag_7to7_bb0__8_i_stall_in_1)) & rstag_7to7_bb0__8_i_stall_local);
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0__17_i_stall_local;
wire [31:0] local_bb0__17_i;

assign local_bb0__17_i = (rstag_7to7_bb0__4_i ? 32'h0 : 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb0__5_i_valid_out;
wire local_bb0__5_i_stall_in;
wire local_bb0__5_i_inputs_ready;
wire local_bb0__5_i_stall_local;
wire [31:0] local_bb0__5_i;

assign local_bb0__5_i_inputs_ready = rstag_7to7_bb0__4_i_valid_out_1;
assign local_bb0__5_i[31:1] = 31'h0;
assign local_bb0__5_i[0] = rstag_7to7_bb0__4_i;
assign local_bb0__5_i_valid_out = local_bb0__5_i_inputs_ready;
assign local_bb0__5_i_stall_local = local_bb0__5_i_stall_in;
assign rstag_7to7_bb0__4_i_stall_in_1 = (|local_bb0__5_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0__18_i_valid_out;
wire local_bb0__18_i_stall_in;
wire local_bb0__18_i_inputs_ready;
wire local_bb0__18_i_stall_local;
wire [31:0] local_bb0__18_i;

assign local_bb0__18_i_inputs_ready = (rstag_7to7_bb0__4_i_valid_out_0 & rstag_7to7_bb0__8_i_valid_out_0);
assign local_bb0__18_i = (rstag_7to7_bb0__8_i ? 32'h1 : (local_bb0__17_i & 32'h100));
assign local_bb0__18_i_valid_out = local_bb0__18_i_inputs_ready;
assign local_bb0__18_i_stall_local = local_bb0__18_i_stall_in;
assign rstag_7to7_bb0__4_i_stall_in_0 = (local_bb0__18_i_stall_local | ~(local_bb0__18_i_inputs_ready));
assign rstag_7to7_bb0__8_i_stall_in_0 = (local_bb0__18_i_stall_local | ~(local_bb0__18_i_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb0__9_i_inputs_ready;
 reg local_bb0__9_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__9_i_valid_out_NO_SHIFT_REG;
wire local_bb0__9_i_stall_in;
wire local_bb0__9_i_output_regs_ready;
 reg [31:0] local_bb0__9_i_NO_SHIFT_REG;
wire local_bb0__9_i_causedstall;

assign local_bb0__9_i_inputs_ready = (local_bb0__5_i_valid_out & rstag_7to7_bb0__8_i_valid_out_1);
assign local_bb0__9_i_output_regs_ready = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__9_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__9_i_stall_in))));
assign local_bb0__5_i_stall_in = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__9_i_output_regs_ready) | ~(local_bb0__9_i_inputs_ready)));
assign rstag_7to7_bb0__8_i_stall_in_1 = (~(local_bb0__9_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__9_i_output_regs_ready) | ~(local_bb0__9_i_inputs_ready)));
assign local_bb0__9_i_causedstall = (local_bb0__9_i_inputs_ready && (~(local_bb0__9_i_output_regs_ready) && !(~(local_bb0__9_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__9_i_NO_SHIFT_REG <= 'x;
		local_bb0__9_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__9_i_NO_SHIFT_REG <= 'x;
			local_bb0__9_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__9_i_output_regs_ready)
			begin
				local_bb0__9_i_NO_SHIFT_REG <= (rstag_7to7_bb0__8_i ? 32'h0 : (local_bb0__5_i & 32'h1));
				local_bb0__9_i_valid_out_NO_SHIFT_REG <= local_bb0__9_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__9_i_stall_in))
				begin
					local_bb0__9_i_valid_out_NO_SHIFT_REG <= local_bb0__9_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__9_i_inputs_ready)
			begin
				local_bb0__9_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0__19_i_inputs_ready;
 reg local_bb0__19_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0__19_i_valid_out_NO_SHIFT_REG;
wire local_bb0__19_i_stall_in;
wire local_bb0__19_i_output_regs_ready;
 reg [31:0] local_bb0__19_i_NO_SHIFT_REG;
wire local_bb0__19_i_causedstall;

assign local_bb0__19_i_inputs_ready = (local_bb0__12_i_valid_out_1_NO_SHIFT_REG & local_bb0__18_i_valid_out);
assign local_bb0__19_i_output_regs_ready = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0__19_i_valid_out_NO_SHIFT_REG) | ~(local_bb0__19_i_stall_in))));
assign local_bb0__12_i_stall_in_1 = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__19_i_output_regs_ready) | ~(local_bb0__19_i_inputs_ready)));
assign local_bb0__18_i_stall_in = (~(local_bb0__19_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0__19_i_output_regs_ready) | ~(local_bb0__19_i_inputs_ready)));
assign local_bb0__19_i_causedstall = (local_bb0__19_i_inputs_ready && (~(local_bb0__19_i_output_regs_ready) && !(~(local_bb0__19_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__19_i_NO_SHIFT_REG <= 'x;
		local_bb0__19_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__19_i_NO_SHIFT_REG <= 'x;
			local_bb0__19_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__19_i_output_regs_ready)
			begin
				local_bb0__19_i_NO_SHIFT_REG <= ((local_bb0__12_i_NO_SHIFT_REG & 1'b0) ? 32'hFFFFFF00 : (local_bb0__18_i & 32'h101));
				local_bb0__19_i_valid_out_NO_SHIFT_REG <= local_bb0__19_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0__19_i_stall_in))
				begin
					local_bb0__19_i_valid_out_NO_SHIFT_REG <= local_bb0__19_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0__19_i_inputs_ready)
			begin
				local_bb0__19_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0__13_i_valid_out;
wire local_bb0__13_i_stall_in;
wire local_bb0__13_i_inputs_ready;
wire local_bb0__13_i_stall_local;
wire [31:0] local_bb0__13_i;

assign local_bb0__13_i_inputs_ready = (local_bb0__12_i_valid_out_0_NO_SHIFT_REG & local_bb0__9_i_valid_out_NO_SHIFT_REG);
assign local_bb0__13_i = ((local_bb0__12_i_NO_SHIFT_REG & 1'b0) ? 32'h0 : (local_bb0__9_i_NO_SHIFT_REG & 32'h1));
assign local_bb0__13_i_valid_out = local_bb0__13_i_inputs_ready;
assign local_bb0__13_i_stall_local = local_bb0__13_i_stall_in;
assign local_bb0__12_i_stall_in_0 = (local_bb0__13_i_stall_local | ~(local_bb0__13_i_inputs_ready));
assign local_bb0__9_i_stall_in = (local_bb0__13_i_stall_local | ~(local_bb0__13_i_inputs_ready));

// This section implements a staging register.
// 
wire rstag_8to8_bb0__19_i_valid_out_0;
wire rstag_8to8_bb0__19_i_stall_in_0;
wire rstag_8to8_bb0__19_i_valid_out_1;
wire rstag_8to8_bb0__19_i_stall_in_1;
wire rstag_8to8_bb0__19_i_inputs_ready;
wire rstag_8to8_bb0__19_i_stall_local;
 reg rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG;
wire rstag_8to8_bb0__19_i_combined_valid;
 reg [31:0] rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_8to8_bb0__19_i;
 reg rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG;
 reg rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG;

assign rstag_8to8_bb0__19_i_inputs_ready = local_bb0__19_i_valid_out_NO_SHIFT_REG;
assign rstag_8to8_bb0__19_i = (rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG ? rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG : (local_bb0__19_i_NO_SHIFT_REG & 32'hFFFFFF01));
assign rstag_8to8_bb0__19_i_combined_valid = (rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG | rstag_8to8_bb0__19_i_inputs_ready);
assign rstag_8to8_bb0__19_i_stall_local = ((rstag_8to8_bb0__19_i_stall_in_0 & ~(rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG)) | (rstag_8to8_bb0__19_i_stall_in_1 & ~(rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG)));
assign rstag_8to8_bb0__19_i_valid_out_0 = (rstag_8to8_bb0__19_i_combined_valid & ~(rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG));
assign rstag_8to8_bb0__19_i_valid_out_1 = (rstag_8to8_bb0__19_i_combined_valid & ~(rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG));
assign local_bb0__19_i_stall_in = (|rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_8to8_bb0__19_i_stall_local)
			begin
				if (~(rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG))
				begin
					rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= rstag_8to8_bb0__19_i_inputs_ready;
				end
			end
			else
			begin
				rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_8to8_bb0__19_i_staging_valid_NO_SHIFT_REG))
		begin
			rstag_8to8_bb0__19_i_staging_reg_NO_SHIFT_REG <= (local_bb0__19_i_NO_SHIFT_REG & 32'hFFFFFF01);
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= 1'b0;
			rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG <= (rstag_8to8_bb0__19_i_combined_valid & (rstag_8to8_bb0__19_i_consumed_0_NO_SHIFT_REG | ~(rstag_8to8_bb0__19_i_stall_in_0)) & rstag_8to8_bb0__19_i_stall_local);
			rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG <= (rstag_8to8_bb0__19_i_combined_valid & (rstag_8to8_bb0__19_i_consumed_1_NO_SHIFT_REG | ~(rstag_8to8_bb0__19_i_stall_in_1)) & rstag_8to8_bb0__19_i_stall_local);
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_fold_i_valid_out;
wire local_bb0_fold_i_stall_in;
wire local_bb0_fold_i_inputs_ready;
wire local_bb0_fold_i_stall_local;
wire [31:0] local_bb0_fold_i;

assign local_bb0_fold_i_inputs_ready = (local_bb0_shr_i_valid_out_1_NO_SHIFT_REG & rstag_8to8_bb0__19_i_valid_out_0);
assign local_bb0_fold_i = ((rstag_8to8_bb0__19_i & 32'hFFFFFF01) + (local_bb0_shr_i_NO_SHIFT_REG & 32'h1FF));
assign local_bb0_fold_i_valid_out = local_bb0_fold_i_inputs_ready;
assign local_bb0_fold_i_stall_local = local_bb0_fold_i_stall_in;
assign local_bb0_shr_i_stall_in_1 = (local_bb0_fold_i_stall_local | ~(local_bb0_fold_i_inputs_ready));
assign rstag_8to8_bb0__19_i_stall_in_0 = (local_bb0_fold_i_stall_local | ~(local_bb0_fold_i_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb0_add_i_inputs_ready;
 reg local_bb0_add_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_add_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_add_i_stall_in_0;
 reg local_bb0_add_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_add_i_stall_in_1;
wire local_bb0_add_i_output_regs_ready;
 reg [31:0] local_bb0_add_i_NO_SHIFT_REG;
wire local_bb0_add_i_causedstall;

assign local_bb0_add_i_inputs_ready = (rstag_8to8_bb0__19_i_valid_out_1 & rstag_4to4_bb0_and1_i_valid_out_0);
assign local_bb0_add_i_output_regs_ready = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_add_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_add_i_stall_in_0)) & (~(local_bb0_add_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_add_i_stall_in_1))));
assign rstag_8to8_bb0__19_i_stall_in_1 = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_add_i_output_regs_ready) | ~(local_bb0_add_i_inputs_ready)));
assign rstag_4to4_bb0_and1_i_stall_in_0 = (~(local_bb0_add_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_add_i_output_regs_ready) | ~(local_bb0_add_i_inputs_ready)));
assign local_bb0_add_i_causedstall = (local_bb0_add_i_inputs_ready && (~(local_bb0_add_i_output_regs_ready) && !(~(local_bb0_add_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add_i_NO_SHIFT_REG <= 'x;
		local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add_i_NO_SHIFT_REG <= 'x;
			local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add_i_output_regs_ready)
			begin
				local_bb0_add_i_NO_SHIFT_REG <= ((rstag_8to8_bb0__19_i & 32'hFFFFFF01) + (rstag_4to4_bb0_and1_i & 32'hFF));
				local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= local_bb0_add_i_inputs_ready;
				local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= local_bb0_add_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_add_i_stall_in_0))
				begin
					local_bb0_add_i_valid_out_0_NO_SHIFT_REG <= local_bb0_add_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_add_i_stall_in_1))
				begin
					local_bb0_add_i_valid_out_1_NO_SHIFT_REG <= local_bb0_add_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_add_i_inputs_ready)
			begin
				local_bb0_add_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_and32_i_inputs_ready;
 reg local_bb0_and32_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_and32_i_valid_out_NO_SHIFT_REG;
wire local_bb0_and32_i_stall_in;
wire local_bb0_and32_i_output_regs_ready;
 reg [31:0] local_bb0_and32_i_NO_SHIFT_REG;
wire local_bb0_and32_i_causedstall;

assign local_bb0_and32_i_inputs_ready = local_bb0_fold_i_valid_out;
assign local_bb0_and32_i_output_regs_ready = (~(local_bb0_and32_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_and32_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_and32_i_stall_in))));
assign local_bb0_fold_i_stall_in = (~(local_bb0_and32_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_and32_i_output_regs_ready) | ~(local_bb0_and32_i_inputs_ready)));
assign local_bb0_and32_i_causedstall = (local_bb0_and32_i_inputs_ready && (~(local_bb0_and32_i_output_regs_ready) && !(~(local_bb0_and32_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and32_i_NO_SHIFT_REG <= 'x;
		local_bb0_and32_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and32_i_NO_SHIFT_REG <= 'x;
			local_bb0_and32_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and32_i_output_regs_ready)
			begin
				local_bb0_and32_i_NO_SHIFT_REG <= (local_bb0_fold_i << 32'h17);
				local_bb0_and32_i_valid_out_NO_SHIFT_REG <= local_bb0_and32_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_and32_i_stall_in))
				begin
					local_bb0_and32_i_valid_out_NO_SHIFT_REG <= local_bb0_and32_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_and32_i_inputs_ready)
			begin
				local_bb0_and32_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_cmp20_i_stall_local;
wire local_bb0_cmp20_i;

assign local_bb0_cmp20_i = ($signed(local_bb0_add_i_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb0_cmp25_i_stall_local;
wire local_bb0_cmp25_i;

assign local_bb0_cmp25_i = ($signed(local_bb0_add_i_NO_SHIFT_REG) < $signed(32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_shl_i_stall_local;
wire [31:0] local_bb0_shl_i;

assign local_bb0_shl_i = ((local_bb0_and32_i_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb0_conv_i_valid_out;
wire local_bb0_conv_i_stall_in;
wire local_bb0_conv_i_inputs_ready;
wire local_bb0_conv_i_stall_local;
wire [31:0] local_bb0_conv_i;

assign local_bb0_conv_i_inputs_ready = local_bb0_add_i_valid_out_0_NO_SHIFT_REG;
assign local_bb0_conv_i[31:1] = 31'h0;
assign local_bb0_conv_i[0] = local_bb0_cmp20_i;
assign local_bb0_conv_i_valid_out = local_bb0_conv_i_inputs_ready;
assign local_bb0_conv_i_stall_local = local_bb0_conv_i_stall_in;
assign local_bb0_add_i_stall_in_0 = (|local_bb0_conv_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0_conv26_i_valid_out;
wire local_bb0_conv26_i_stall_in;
wire local_bb0_conv26_i_inputs_ready;
wire local_bb0_conv26_i_stall_local;
wire [31:0] local_bb0_conv26_i;

assign local_bb0_conv26_i_inputs_ready = local_bb0_add_i_valid_out_1_NO_SHIFT_REG;
assign local_bb0_conv26_i[31:1] = 31'h0;
assign local_bb0_conv26_i[0] = local_bb0_cmp25_i;
assign local_bb0_conv26_i_valid_out = local_bb0_conv26_i_inputs_ready;
assign local_bb0_conv26_i_stall_local = local_bb0_conv26_i_stall_in;
assign local_bb0_add_i_stall_in_1 = (|local_bb0_conv26_i_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb0_or34_i_stall_local;
wire [31:0] local_bb0_or34_i;

assign local_bb0_or34_i = ((local_bb0_shl_i & 32'h7F800000) | (local_bb0_and33_i_NO_SHIFT_REG & 32'h807FFFFF));

// This section implements a registered operation.
// 
wire local_bb0_or_i_inputs_ready;
 reg local_bb0_or_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_or_i_valid_out_0_NO_SHIFT_REG;
wire local_bb0_or_i_stall_in_0;
 reg local_bb0_or_i_valid_out_1_NO_SHIFT_REG;
wire local_bb0_or_i_stall_in_1;
wire local_bb0_or_i_output_regs_ready;
 reg [31:0] local_bb0_or_i_NO_SHIFT_REG;
wire local_bb0_or_i_causedstall;

assign local_bb0_or_i_inputs_ready = (local_bb0_conv_i_valid_out & local_bb0_conv22_i_valid_out_NO_SHIFT_REG);
assign local_bb0_or_i_output_regs_ready = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_or_i_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_or_i_stall_in_0)) & (~(local_bb0_or_i_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_or_i_stall_in_1))));
assign local_bb0_conv_i_stall_in = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or_i_output_regs_ready) | ~(local_bb0_or_i_inputs_ready)));
assign local_bb0_conv22_i_stall_in = (~(local_bb0_or_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or_i_output_regs_ready) | ~(local_bb0_or_i_inputs_ready)));
assign local_bb0_or_i_causedstall = (local_bb0_or_i_inputs_ready && (~(local_bb0_or_i_output_regs_ready) && !(~(local_bb0_or_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or_i_NO_SHIFT_REG <= 'x;
		local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or_i_NO_SHIFT_REG <= 'x;
			local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or_i_output_regs_ready)
			begin
				local_bb0_or_i_NO_SHIFT_REG <= ((local_bb0_conv_i & 32'h1) | (local_bb0_conv22_i_NO_SHIFT_REG & 32'h1));
				local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= local_bb0_or_i_inputs_ready;
				local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= local_bb0_or_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_or_i_stall_in_0))
				begin
					local_bb0_or_i_valid_out_0_NO_SHIFT_REG <= local_bb0_or_i_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_or_i_stall_in_1))
				begin
					local_bb0_or_i_valid_out_1_NO_SHIFT_REG <= local_bb0_or_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or_i_inputs_ready)
			begin
				local_bb0_or_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_or29_i_inputs_ready;
 reg local_bb0_or29_i_wii_reg_NO_SHIFT_REG;
 reg local_bb0_or29_i_valid_out_NO_SHIFT_REG;
wire local_bb0_or29_i_stall_in;
wire local_bb0_or29_i_output_regs_ready;
 reg [31:0] local_bb0_or29_i_NO_SHIFT_REG;
wire local_bb0_or29_i_causedstall;

assign local_bb0_or29_i_inputs_ready = (local_bb0_conv26_i_valid_out & local_bb0__13_i_valid_out);
assign local_bb0_or29_i_output_regs_ready = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_or29_i_valid_out_NO_SHIFT_REG) | ~(local_bb0_or29_i_stall_in))));
assign local_bb0_conv26_i_stall_in = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or29_i_output_regs_ready) | ~(local_bb0_or29_i_inputs_ready)));
assign local_bb0__13_i_stall_in = (~(local_bb0_or29_i_wii_reg_NO_SHIFT_REG) & (~(local_bb0_or29_i_output_regs_ready) | ~(local_bb0_or29_i_inputs_ready)));
assign local_bb0_or29_i_causedstall = (local_bb0_or29_i_inputs_ready && (~(local_bb0_or29_i_output_regs_ready) && !(~(local_bb0_or29_i_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or29_i_NO_SHIFT_REG <= 'x;
		local_bb0_or29_i_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or29_i_NO_SHIFT_REG <= 'x;
			local_bb0_or29_i_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or29_i_output_regs_ready)
			begin
				local_bb0_or29_i_NO_SHIFT_REG <= ((local_bb0_conv26_i & 32'h1) | (local_bb0__13_i & 32'h1));
				local_bb0_or29_i_valid_out_NO_SHIFT_REG <= local_bb0_or29_i_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_or29_i_stall_in))
				begin
					local_bb0_or29_i_valid_out_NO_SHIFT_REG <= local_bb0_or29_i_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_or29_i_inputs_ready)
			begin
				local_bb0_or29_i_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb0_or45_i_stall_local;
wire [31:0] local_bb0_or45_i;

assign local_bb0_or45_i = ((local_bb0_or_i_NO_SHIFT_REG & 32'h1) | (local_bb0_conv44_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_or39_i_stall_local;
wire [31:0] local_bb0_or39_i;

assign local_bb0_or39_i = ((local_bb0_or29_i_NO_SHIFT_REG & 32'h1) | (local_bb0_or_i_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb0_tobool46_i_stall_local;
wire local_bb0_tobool46_i;

assign local_bb0_tobool46_i = ((local_bb0_or45_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_tobool40_i_stall_local;
wire local_bb0_tobool40_i;

assign local_bb0_tobool40_i = ((local_bb0_or39_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_cond47_i_stall_local;
wire [31:0] local_bb0_cond47_i;

assign local_bb0_cond47_i = (local_bb0_tobool46_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb0_cond_i_stall_local;
wire [31:0] local_bb0_cond_i;

assign local_bb0_cond_i = (local_bb0_tobool40_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb0_or52_i_stall_local;
wire [31:0] local_bb0_or52_i;

assign local_bb0_or52_i = ((local_bb0_cond47_i & 32'h7F800000) | (local_bb0_cond50_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb0_and51_i_stall_local;
wire [31:0] local_bb0_and51_i;

assign local_bb0_and51_i = ((local_bb0_cond_i | 32'h80000000) & local_bb0_or34_i);

// This section implements an unregistered operation.
// 
wire local_bb0_or53_i_stall_local;
wire [31:0] local_bb0_or53_i;

assign local_bb0_or53_i = ((local_bb0_or52_i & 32'h7FC00000) | local_bb0_and51_i);

// This section implements an unregistered operation.
// 
wire local_bb0_var__u2_valid_out;
wire local_bb0_var__u2_stall_in;
wire local_bb0_var__u2_inputs_ready;
wire local_bb0_var__u2_stall_local;
wire [31:0] local_bb0_var__u2;

assign local_bb0_var__u2_inputs_ready = (local_bb0_and33_i_valid_out_NO_SHIFT_REG & local_bb0_and32_i_valid_out_NO_SHIFT_REG & local_bb0___i_valid_out_1_NO_SHIFT_REG & local_bb0___i_valid_out_0_NO_SHIFT_REG & local_bb0_or_i_valid_out_1_NO_SHIFT_REG & local_bb0_or29_i_valid_out_NO_SHIFT_REG & local_bb0_or_i_valid_out_0_NO_SHIFT_REG);
assign local_bb0_var__u2 = local_bb0_or53_i;
assign local_bb0_var__u2_valid_out = local_bb0_var__u2_inputs_ready;
assign local_bb0_var__u2_stall_local = local_bb0_var__u2_stall_in;
assign local_bb0_and33_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_and32_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0___i_stall_in_1 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0___i_stall_in_0 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or_i_stall_in_1 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or29_i_stall_in = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));
assign local_bb0_or_i_stall_in_0 = (local_bb0_var__u2_stall_local | ~(local_bb0_var__u2_inputs_ready));

// This section implements a staging register.
// 
wire rstag_10to10_bb0_var__u2_valid_out;
wire rstag_10to10_bb0_var__u2_stall_in;
wire rstag_10to10_bb0_var__u2_inputs_ready;
wire rstag_10to10_bb0_var__u2_stall_local;
 reg rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG;
wire rstag_10to10_bb0_var__u2_combined_valid;
 reg [31:0] rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_10to10_bb0_var__u2;

assign rstag_10to10_bb0_var__u2_inputs_ready = local_bb0_var__u2_valid_out;
assign rstag_10to10_bb0_var__u2 = (rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG ? rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG : local_bb0_var__u2);
assign rstag_10to10_bb0_var__u2_combined_valid = (rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG | rstag_10to10_bb0_var__u2_inputs_ready);
assign rstag_10to10_bb0_var__u2_valid_out = rstag_10to10_bb0_var__u2_combined_valid;
assign rstag_10to10_bb0_var__u2_stall_local = rstag_10to10_bb0_var__u2_stall_in;
assign local_bb0_var__u2_stall_in = (|rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (start)
		begin
			rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (rstag_10to10_bb0_var__u2_stall_local)
			begin
				if (~(rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG))
				begin
					rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= rstag_10to10_bb0_var__u2_inputs_ready;
				end
			end
			else
			begin
				rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
			end
		end
		if (~(rstag_10to10_bb0_var__u2_staging_valid_NO_SHIFT_REG))
		begin
			rstag_10to10_bb0_var__u2_staging_reg_NO_SHIFT_REG <= local_bb0_var__u2;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_mul48_inputs_ready;
 reg local_bb0_mul48_wii_reg_NO_SHIFT_REG;
 reg local_bb0_mul48_valid_out_NO_SHIFT_REG;
wire local_bb0_mul48_stall_in;
wire local_bb0_mul48_output_regs_ready;
wire [31:0] local_bb0_mul48;
 reg local_bb0_mul48_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb0_mul48_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb0_mul48_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb0_mul48_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb0_mul48_valid_pipe_4_NO_SHIFT_REG;
wire local_bb0_mul48_causedstall;

acl_fp_mul_ll_s5 fp_module_local_bb0_mul48 (
	.clock(clock),
	.dataa(rstag_10to10_bb0_var__u2),
	.datab(input_e_d),
	.enable(local_bb0_mul48_output_regs_ready),
	.result(local_bb0_mul48)
);


assign local_bb0_mul48_inputs_ready = (merge_node_valid_out_5_NO_SHIFT_REG & rstag_10to10_bb0_var__u2_valid_out);
assign local_bb0_mul48_output_regs_ready = (~(local_bb0_mul48_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_mul48_valid_out_NO_SHIFT_REG) | ~(local_bb0_mul48_stall_in))));
assign merge_node_stall_in_5 = (~(local_bb0_mul48_wii_reg_NO_SHIFT_REG) & (~(local_bb0_mul48_output_regs_ready) | ~(local_bb0_mul48_inputs_ready)));
assign rstag_10to10_bb0_var__u2_stall_in = (~(local_bb0_mul48_wii_reg_NO_SHIFT_REG) & (~(local_bb0_mul48_output_regs_ready) | ~(local_bb0_mul48_inputs_ready)));
assign local_bb0_mul48_causedstall = (local_bb0_mul48_inputs_ready && (~(local_bb0_mul48_output_regs_ready) && !(~(local_bb0_mul48_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul48_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul48_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul48_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul48_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb0_mul48_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul48_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul48_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul48_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul48_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
			local_bb0_mul48_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul48_output_regs_ready)
			begin
				local_bb0_mul48_valid_pipe_0_NO_SHIFT_REG <= local_bb0_mul48_inputs_ready;
				local_bb0_mul48_valid_pipe_1_NO_SHIFT_REG <= local_bb0_mul48_valid_pipe_0_NO_SHIFT_REG;
				local_bb0_mul48_valid_pipe_2_NO_SHIFT_REG <= local_bb0_mul48_valid_pipe_1_NO_SHIFT_REG;
				local_bb0_mul48_valid_pipe_3_NO_SHIFT_REG <= local_bb0_mul48_valid_pipe_2_NO_SHIFT_REG;
				local_bb0_mul48_valid_pipe_4_NO_SHIFT_REG <= local_bb0_mul48_valid_pipe_3_NO_SHIFT_REG;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul48_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul48_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul48_output_regs_ready)
			begin
				local_bb0_mul48_valid_out_NO_SHIFT_REG <= local_bb0_mul48_valid_pipe_4_NO_SHIFT_REG;
			end
			else
			begin
				if (~(local_bb0_mul48_stall_in))
				begin
					local_bb0_mul48_valid_out_NO_SHIFT_REG <= local_bb0_mul48_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_mul48_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_mul48_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_mul48_valid_pipe_4_NO_SHIFT_REG)
			begin
				local_bb0_mul48_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg lvb_bb0_cmp1526_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_sub24_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_sub27_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb0_mul48_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb0_var__reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb0_var__u0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb0_var__u0_valid_out_NO_SHIFT_REG & local_bb0_var__valid_out_NO_SHIFT_REG & local_bb0_mul48_valid_out_NO_SHIFT_REG & local_bb0_sub27_valid_out_NO_SHIFT_REG & local_bb0_sub24_valid_out_NO_SHIFT_REG & local_bb0_cmp1526_valid_out_NO_SHIFT_REG & merge_node_valid_out_7_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb0_var__u0_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_var__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_mul48_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_sub27_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_sub24_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_cmp1526_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign merge_node_stall_in_7 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb0_cmp1526 = lvb_bb0_cmp1526_reg_NO_SHIFT_REG;
assign lvb_bb0_sub24 = lvb_bb0_sub24_reg_NO_SHIFT_REG;
assign lvb_bb0_sub27 = lvb_bb0_sub27_reg_NO_SHIFT_REG;
assign lvb_bb0_mul48 = lvb_bb0_mul48_reg_NO_SHIFT_REG;
assign lvb_bb0_var_ = lvb_bb0_var__reg_NO_SHIFT_REG;
assign lvb_bb0_var__u0 = lvb_bb0_var__u0_reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb0_cmp1526_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_sub24_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_sub27_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_mul48_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_var__u0_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb0_cmp1526_reg_NO_SHIFT_REG <= local_bb0_cmp1526_NO_SHIFT_REG;
			lvb_bb0_sub24_reg_NO_SHIFT_REG <= local_bb0_sub24_NO_SHIFT_REG;
			lvb_bb0_sub27_reg_NO_SHIFT_REG <= local_bb0_sub27_NO_SHIFT_REG;
			lvb_bb0_mul48_reg_NO_SHIFT_REG <= local_bb0_mul48;
			lvb_bb0_var__reg_NO_SHIFT_REG <= local_bb0_var__NO_SHIFT_REG;
			lvb_bb0_var__u0_reg_NO_SHIFT_REG <= local_bb0_var__u0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_1
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_global_size_1,
		input [31:0] 		input_global_size_0,
		input 		input_wii_cmp1526,
		input [31:0] 		input_wii_sub24,
		input [31:0] 		input_wii_sub27,
		input [31:0] 		input_wii_mul48,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u3,
		input 		valid_in_0,
		output 		stall_out_0,
		input [31:0] 		input_pos_y_0_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [31:0] 		input_pos_y_0_1,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start,
		output [31:0] 		ffwd_0_0,
		output 		ffwd_1_0,
		output [31:0] 		ffwd_2_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pos_y_0_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_pos_y_0_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_pos_y_0_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_pos_y_0_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_pos_y_0_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_pos_y_0_0_staging_reg_NO_SHIFT_REG <= input_pos_y_0_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_pos_y_0_1_staging_reg_NO_SHIFT_REG <= input_pos_y_0_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_pos_y_0_NO_SHIFT_REG <= input_pos_y_0_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_pos_y_0_NO_SHIFT_REG <= input_pos_y_0_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_pos_y_0_NO_SHIFT_REG <= input_pos_y_0_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_pos_y_0_NO_SHIFT_REG <= input_pos_y_0_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1_cmp_valid_out;
wire local_bb1_cmp_stall_in;
wire local_bb1_cmp_inputs_ready;
wire local_bb1_cmp_stall_local;
wire local_bb1_cmp;

assign local_bb1_cmp_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb1_cmp = (local_lvm_pos_y_0_NO_SHIFT_REG < input_global_size_1);
assign local_bb1_cmp_valid_out = local_bb1_cmp_inputs_ready;
assign local_bb1_cmp_stall_local = local_bb1_cmp_stall_in;
assign merge_node_stall_in_0 = (|local_bb1_cmp_stall_local);

// This section implements a registered operation.
// 
wire local_bb1_mul_inputs_ready;
 reg local_bb1_mul_valid_out_NO_SHIFT_REG;
wire local_bb1_mul_stall_in;
wire local_bb1_mul_output_regs_ready;
wire [31:0] local_bb1_mul;
 reg local_bb1_mul_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb1_mul_valid_pipe_1_NO_SHIFT_REG;
wire local_bb1_mul_causedstall;

acl_int_mult int_module_local_bb1_mul (
	.clock(clock),
	.dataa(local_lvm_pos_y_0_NO_SHIFT_REG),
	.datab(input_global_size_0),
	.enable(local_bb1_mul_output_regs_ready),
	.result(local_bb1_mul)
);

defparam int_module_local_bb1_mul.INPUT1_WIDTH = 32;
defparam int_module_local_bb1_mul.INPUT2_WIDTH = 32;
defparam int_module_local_bb1_mul.OUTPUT_WIDTH = 32;
defparam int_module_local_bb1_mul.LATENCY = 3;
defparam int_module_local_bb1_mul.SIGNED = 0;

assign local_bb1_mul_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb1_mul_output_regs_ready = (&(~(local_bb1_mul_valid_out_NO_SHIFT_REG) | ~(local_bb1_mul_stall_in)));
assign merge_node_stall_in_1 = (~(local_bb1_mul_output_regs_ready) | ~(local_bb1_mul_inputs_ready));
assign local_bb1_mul_causedstall = (local_bb1_mul_inputs_ready && (~(local_bb1_mul_output_regs_ready) && !(~(local_bb1_mul_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb1_mul_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul_output_regs_ready)
		begin
			local_bb1_mul_valid_pipe_0_NO_SHIFT_REG <= local_bb1_mul_inputs_ready;
			local_bb1_mul_valid_pipe_1_NO_SHIFT_REG <= local_bb1_mul_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul_output_regs_ready)
		begin
			local_bb1_mul_valid_out_NO_SHIFT_REG <= local_bb1_mul_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb1_mul_stall_in))
			begin
				local_bb1_mul_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1__pos_y_0_valid_out;
wire local_bb1__pos_y_0_stall_in;
wire local_bb1__pos_y_0_inputs_ready;
wire local_bb1__pos_y_0_stall_local;
 reg [31:0] ffwd_0_0_reg_NO_SHIFT_REG;

assign local_bb1__pos_y_0_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign ffwd_0_0 = ffwd_0_0_reg_NO_SHIFT_REG;
assign local_bb1__pos_y_0_valid_out = local_bb1__pos_y_0_inputs_ready;
assign local_bb1__pos_y_0_stall_local = local_bb1__pos_y_0_stall_in;
assign merge_node_stall_in_2 = (|local_bb1__pos_y_0_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb1__pos_y_0_inputs_ready))
	begin
		ffwd_0_0_reg_NO_SHIFT_REG <= local_lvm_pos_y_0_NO_SHIFT_REG;
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb1_cmp_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb1_cmp_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb1_cmp_0_NO_SHIFT_REG;
 logic rnode_1to2_bb1_cmp_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb1_cmp_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_cmp_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_cmp_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb1_cmp_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb1_cmp_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb1_cmp_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb1_cmp_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb1_cmp_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb1_cmp_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb1_cmp),
	.data_out(rnode_1to2_bb1_cmp_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb1_cmp_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb1_cmp_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb1_cmp_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb1_cmp_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb1_cmp_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb1_cmp_valid_out;
assign local_bb1_cmp_stall_in = rnode_1to2_bb1_cmp_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb1_cmp_0_NO_SHIFT_REG = rnode_1to2_bb1_cmp_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb1_cmp_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb1_cmp_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb1_cmp_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb1_cmp_0_valid_out_reg_2_NO_SHIFT_REG;

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_4to4_bb1_mul_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb1_mul_0_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb1_mul_0_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb1_mul_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_4to4_bb1_mul_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to4_bb1_mul_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to4_bb1_mul_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_4to4_bb1_mul_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_4to4_bb1_mul_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb1_mul),
	.data_out(rnode_4to4_bb1_mul_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_4to4_bb1_mul_0_reg_4_fifo.DEPTH = 3;
defparam rnode_4to4_bb1_mul_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_4to4_bb1_mul_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to4_bb1_mul_0_reg_4_fifo.IMPL = "zl_reg";

assign rnode_4to4_bb1_mul_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb1_mul_valid_out_NO_SHIFT_REG;
assign local_bb1_mul_stall_in = rnode_4to4_bb1_mul_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb1_mul_0_NO_SHIFT_REG = rnode_4to4_bb1_mul_0_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb1_mul_0_stall_in_reg_4_NO_SHIFT_REG = rnode_4to4_bb1_mul_0_stall_in_NO_SHIFT_REG;
assign rnode_4to4_bb1_mul_0_valid_out_NO_SHIFT_REG = rnode_4to4_bb1_mul_0_valid_out_reg_4_NO_SHIFT_REG;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_bb1__pos_y_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to4_bb1__pos_y_0_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to4_bb1__pos_y_0_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to4_bb1__pos_y_0_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1__pos_y_0_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_bb1__pos_y_0_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_1to4_bb1__pos_y_0_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_bb1__pos_y_0_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_bb1__pos_y_0_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_bb1__pos_y_0_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_bb1__pos_y_0_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to4_bb1__pos_y_0_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_bb1__pos_y_0_0_reg_4_fifo.DATA_WIDTH = 0;
defparam rnode_1to4_bb1__pos_y_0_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_bb1__pos_y_0_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_bb1__pos_y_0_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb1__pos_y_0_valid_out;
assign local_bb1__pos_y_0_stall_in = rnode_1to4_bb1__pos_y_0_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_bb1__pos_y_0_0_stall_in_reg_4_NO_SHIFT_REG = rnode_1to4_bb1__pos_y_0_0_stall_in_NO_SHIFT_REG;
assign rnode_1to4_bb1__pos_y_0_0_valid_out_NO_SHIFT_REG = rnode_1to4_bb1__pos_y_0_0_valid_out_reg_4_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb1__cmp_valid_out;
wire local_bb1__cmp_stall_in;
wire local_bb1__cmp_inputs_ready;
wire local_bb1__cmp_stall_local;
 reg ffwd_1_0_reg_NO_SHIFT_REG;

assign local_bb1__cmp_inputs_ready = rnode_1to2_bb1_cmp_0_valid_out_NO_SHIFT_REG;
assign ffwd_1_0 = ffwd_1_0_reg_NO_SHIFT_REG;
assign local_bb1__cmp_valid_out = local_bb1__cmp_inputs_ready;
assign local_bb1__cmp_stall_local = local_bb1__cmp_stall_in;
assign rnode_1to2_bb1_cmp_0_stall_in_NO_SHIFT_REG = (|local_bb1__cmp_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb1__cmp_inputs_ready))
	begin
		ffwd_1_0_reg_NO_SHIFT_REG <= rnode_1to2_bb1_cmp_0_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb1__mul_valid_out;
wire local_bb1__mul_stall_in;
wire local_bb1__mul_inputs_ready;
wire local_bb1__mul_stall_local;
 reg [31:0] ffwd_2_0_reg_NO_SHIFT_REG;

assign local_bb1__mul_inputs_ready = rnode_4to4_bb1_mul_0_valid_out_NO_SHIFT_REG;
assign ffwd_2_0 = ffwd_2_0_reg_NO_SHIFT_REG;
assign local_bb1__mul_valid_out = local_bb1__mul_inputs_ready;
assign local_bb1__mul_stall_local = local_bb1__mul_stall_in;
assign rnode_4to4_bb1_mul_0_stall_in_NO_SHIFT_REG = (|local_bb1__mul_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb1__mul_inputs_ready))
	begin
		ffwd_2_0_reg_NO_SHIFT_REG <= rnode_4to4_bb1_mul_0_NO_SHIFT_REG;
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_2to4_bb1__cmp_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to4_bb1__cmp_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to4_bb1__cmp_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to4_bb1__cmp_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_2to4_bb1__cmp_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_2to4_bb1__cmp_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_2to4_bb1__cmp_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to4_bb1__cmp_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to4_bb1__cmp_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_2to4_bb1__cmp_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_2to4_bb1__cmp_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to4_bb1__cmp_0_reg_4_fifo.DEPTH = 3;
defparam rnode_2to4_bb1__cmp_0_reg_4_fifo.DATA_WIDTH = 0;
defparam rnode_2to4_bb1__cmp_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_2to4_bb1__cmp_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_2to4_bb1__cmp_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb1__cmp_valid_out;
assign local_bb1__cmp_stall_in = rnode_2to4_bb1__cmp_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_2to4_bb1__cmp_0_stall_in_reg_4_NO_SHIFT_REG = rnode_2to4_bb1__cmp_0_stall_in_NO_SHIFT_REG;
assign rnode_2to4_bb1__cmp_0_valid_out_NO_SHIFT_REG = rnode_2to4_bb1__cmp_0_valid_out_reg_4_NO_SHIFT_REG;

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;

assign branch_var__inputs_ready = (local_bb1__mul_valid_out & rnode_2to4_bb1__cmp_0_valid_out_NO_SHIFT_REG & rnode_1to4_bb1__pos_y_0_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb1__mul_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_2to4_bb1__cmp_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to4_bb1__pos_y_0_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_2
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_global_size_0,
		input [63:0] 		input_in,
		input 		input_wii_cmp1526,
		input [31:0] 		input_wii_sub24,
		input [31:0] 		input_wii_sub27,
		input [31:0] 		input_wii_mul48,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u4,
		input 		valid_in_0,
		output 		stall_out_0,
		input [63:0] 		input_indvars_iv39_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [63:0] 		input_indvars_iv39_1,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start,
		input [31:0] 		ffwd_2_0,
		output [63:0] 		ffwd_3_0,
		input 		ffwd_1_0,
		output [31:0] 		ffwd_4_0,
		output [63:0] 		ffwd_6_0,
		output 		ffwd_5_0,
		input [511:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [32:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [511:0] 		avm_local_bb2_ld__writedata,
		output [63:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		output 		local_bb2_ld__active,
		input 		clock2x,
		output [31:0] 		ffwd_7_0,
		output 		ffwd_8_0,
		output 		ffwd_9_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv39_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv39_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv39_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_indvars_iv39_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_indvars_iv39_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_indvars_iv39_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv39_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_indvars_iv39_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv39_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_indvars_iv39_NO_SHIFT_REG <= input_indvars_iv39_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_indvars_iv39_NO_SHIFT_REG <= input_indvars_iv39_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_indvars_iv39_NO_SHIFT_REG <= input_indvars_iv39_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_indvars_iv39_NO_SHIFT_REG <= input_indvars_iv39_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__stall_local;
wire [31:0] local_bb2_var_;

assign local_bb2_var_ = local_lvm_indvars_iv39_NO_SHIFT_REG[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_mul5_acl_ffwd_dest_i32_2_stall_local;
wire [31:0] local_bb2_mul5_acl_ffwd_dest_i32_2;

assign local_bb2_mul5_acl_ffwd_dest_i32_2 = ffwd_2_0;

// This section implements an unregistered operation.
// 
wire local_bb2__indvars_iv39_valid_out;
wire local_bb2__indvars_iv39_stall_in;
wire local_bb2__indvars_iv39_inputs_ready;
wire local_bb2__indvars_iv39_stall_local;
 reg [63:0] ffwd_3_0_reg_NO_SHIFT_REG;

assign local_bb2__indvars_iv39_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign ffwd_3_0 = ffwd_3_0_reg_NO_SHIFT_REG;
assign local_bb2__indvars_iv39_valid_out = local_bb2__indvars_iv39_inputs_ready;
assign local_bb2__indvars_iv39_stall_local = local_bb2__indvars_iv39_stall_in;
assign merge_node_stall_in_2 = (|local_bb2__indvars_iv39_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2__indvars_iv39_inputs_ready))
	begin
		ffwd_3_0_reg_NO_SHIFT_REG <= local_lvm_indvars_iv39_NO_SHIFT_REG;
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_fifo.DEPTH = 3;
defparam rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_reg_3_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_3_NO_SHIFT_REG;
assign merge_node_stall_in_3 = rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_in_reg_3_NO_SHIFT_REG = rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_in_NO_SHIFT_REG;
assign rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_valid_out_NO_SHIFT_REG = rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_valid_out_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_var__valid_out_1;
wire local_bb2_var__stall_in_1;
wire local_bb2_add_valid_out;
wire local_bb2_add_stall_in;
wire local_bb2_add_inputs_ready;
wire local_bb2_add_stall_local;
wire [31:0] local_bb2_add;
 reg local_bb2_var__consumed_1_NO_SHIFT_REG;
 reg local_bb2_add_consumed_0_NO_SHIFT_REG;

assign local_bb2_add_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign local_bb2_add = (local_bb2_var_ + local_bb2_mul5_acl_ffwd_dest_i32_2);
assign local_bb2_add_stall_local = ((local_bb2_var__stall_in_1 & ~(local_bb2_var__consumed_1_NO_SHIFT_REG)) | (local_bb2_add_stall_in & ~(local_bb2_add_consumed_0_NO_SHIFT_REG)));
assign local_bb2_var__valid_out_1 = (local_bb2_add_inputs_ready & ~(local_bb2_var__consumed_1_NO_SHIFT_REG));
assign local_bb2_add_valid_out = (local_bb2_add_inputs_ready & ~(local_bb2_add_consumed_0_NO_SHIFT_REG));
assign merge_node_stall_in_0 = (local_bb2_add_stall_local | ~(local_bb2_add_inputs_ready));
assign merge_node_stall_in_1 = (local_bb2_add_stall_local | ~(local_bb2_add_inputs_ready));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_var__consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_var__consumed_1_NO_SHIFT_REG <= (local_bb2_add_inputs_ready & (local_bb2_var__consumed_1_NO_SHIFT_REG | ~(local_bb2_var__stall_in_1)) & local_bb2_add_stall_local);
		local_bb2_add_consumed_0_NO_SHIFT_REG <= (local_bb2_add_inputs_ready & (local_bb2_add_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_stall_in)) & local_bb2_add_stall_local);
	end
end


// Register node:
//  * latency = 164
//  * capacity = 164
 logic rnode_1to165_bb2__indvars_iv39_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to165_bb2__indvars_iv39_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to165_bb2__indvars_iv39_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to165_bb2__indvars_iv39_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_1to165_bb2__indvars_iv39_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_1to165_bb2__indvars_iv39_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_1to165_bb2__indvars_iv39_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to165_bb2__indvars_iv39_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to165_bb2__indvars_iv39_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_1to165_bb2__indvars_iv39_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_1to165_bb2__indvars_iv39_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to165_bb2__indvars_iv39_0_reg_165_fifo.DEPTH = 165;
defparam rnode_1to165_bb2__indvars_iv39_0_reg_165_fifo.DATA_WIDTH = 0;
defparam rnode_1to165_bb2__indvars_iv39_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to165_bb2__indvars_iv39_0_reg_165_fifo.IMPL = "ram";

assign rnode_1to165_bb2__indvars_iv39_0_reg_165_inputs_ready_NO_SHIFT_REG = local_bb2__indvars_iv39_valid_out;
assign local_bb2__indvars_iv39_stall_in = rnode_1to165_bb2__indvars_iv39_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_1to165_bb2__indvars_iv39_0_stall_in_reg_165_NO_SHIFT_REG = rnode_1to165_bb2__indvars_iv39_0_stall_in_NO_SHIFT_REG;
assign rnode_1to165_bb2__indvars_iv39_0_valid_out_NO_SHIFT_REG = rnode_1to165_bb2__indvars_iv39_0_valid_out_reg_165_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp4_acl_ffwd_dest_i1_1_stall_local;
wire local_bb2_cmp4_acl_ffwd_dest_i1_1;

assign local_bb2_cmp4_acl_ffwd_dest_i1_1 = ffwd_1_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb2_var__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_var__0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_var__1_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_var__0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_var__0_stall_out_reg_2_NO_SHIFT_REG;
 reg rnode_1to2_bb2_var__0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to2_bb2_var__0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb2_var__0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb2_var__0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb2_var__0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb2_var__0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb2_var__0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb2_var_),
	.data_out(rnode_1to2_bb2_var__0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb2_var__0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb2_var__0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb2_var__0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb2_var__0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb2_var__0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb2_var__valid_out_1;
assign local_bb2_var__stall_in_1 = rnode_1to2_bb2_var__0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__0_stall_in_0_reg_2_NO_SHIFT_REG = ((rnode_1to2_bb2_var__0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__0_consumed_0_NO_SHIFT_REG)) | (rnode_1to2_bb2_var__0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to2_bb2_var__0_valid_out_0_NO_SHIFT_REG = (rnode_1to2_bb2_var__0_valid_out_0_reg_2_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__0_consumed_0_NO_SHIFT_REG));
assign rnode_1to2_bb2_var__0_valid_out_1_NO_SHIFT_REG = (rnode_1to2_bb2_var__0_valid_out_0_reg_2_NO_SHIFT_REG & ~(rnode_1to2_bb2_var__0_consumed_1_NO_SHIFT_REG));
assign rnode_1to2_bb2_var__0_NO_SHIFT_REG = rnode_1to2_bb2_var__0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_var__1_NO_SHIFT_REG = rnode_1to2_bb2_var__0_reg_2_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to2_bb2_var__0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to2_bb2_var__0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to2_bb2_var__0_consumed_0_NO_SHIFT_REG <= (rnode_1to2_bb2_var__0_valid_out_0_reg_2_NO_SHIFT_REG & (rnode_1to2_bb2_var__0_consumed_0_NO_SHIFT_REG | ~(rnode_1to2_bb2_var__0_stall_in_0_NO_SHIFT_REG)) & rnode_1to2_bb2_var__0_stall_in_0_reg_2_NO_SHIFT_REG);
		rnode_1to2_bb2_var__0_consumed_1_NO_SHIFT_REG <= (rnode_1to2_bb2_var__0_valid_out_0_reg_2_NO_SHIFT_REG & (rnode_1to2_bb2_var__0_consumed_1_NO_SHIFT_REG | ~(rnode_1to2_bb2_var__0_stall_in_1_NO_SHIFT_REG)) & rnode_1to2_bb2_var__0_stall_in_0_reg_2_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb2_add_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_add_0_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb2_add_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb2_add_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb2_add_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb2_add_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb2_add_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb2_add_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb2_add_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb2_add),
	.data_out(rnode_1to2_bb2_add_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb2_add_0_reg_2_fifo.DEPTH = 2;
defparam rnode_1to2_bb2_add_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb2_add_0_reg_2_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to2_bb2_add_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb2_add_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb2_add_valid_out;
assign local_bb2_add_stall_in = rnode_1to2_bb2_add_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_add_0_NO_SHIFT_REG = rnode_1to2_bb2_add_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb2_add_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb2_add_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb2_add_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb2_add_0_valid_out_reg_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp5_valid_out;
wire local_bb2_cmp5_stall_in;
wire local_bb2_cmp5_inputs_ready;
wire local_bb2_cmp5_stall_local;
wire local_bb2_cmp5;

assign local_bb2_cmp5_inputs_ready = rnode_1to2_bb2_var__0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_cmp5 = (rnode_1to2_bb2_var__0_NO_SHIFT_REG < input_global_size_0);
assign local_bb2_cmp5_valid_out = local_bb2_cmp5_inputs_ready;
assign local_bb2_cmp5_stall_local = local_bb2_cmp5_stall_in;
assign rnode_1to2_bb2_var__0_stall_in_0_NO_SHIFT_REG = (|local_bb2_cmp5_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb2___valid_out;
wire local_bb2___stall_in;
wire local_bb2___inputs_ready;
wire local_bb2___stall_local;
 reg [31:0] ffwd_4_0_reg_NO_SHIFT_REG;

assign local_bb2___inputs_ready = rnode_1to2_bb2_var__0_valid_out_1_NO_SHIFT_REG;
assign ffwd_4_0 = ffwd_4_0_reg_NO_SHIFT_REG;
assign local_bb2___valid_out = local_bb2___inputs_ready;
assign local_bb2___stall_local = local_bb2___stall_in;
assign rnode_1to2_bb2_var__0_stall_in_1_NO_SHIFT_REG = (|local_bb2___stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___inputs_ready))
	begin
		ffwd_4_0_reg_NO_SHIFT_REG <= rnode_1to2_bb2_var__1_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_idxprom_stall_local;
wire [63:0] local_bb2_idxprom;

assign local_bb2_idxprom[63:32] = 32'h0;
assign local_bb2_idxprom[31:0] = rnode_1to2_bb2_add_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb2_cmp5_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb2_cmp5_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb2_cmp5_0_NO_SHIFT_REG;
 logic rnode_2to3_bb2_cmp5_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb2_cmp5_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_cmp5_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_cmp5_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_cmp5_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb2_cmp5_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb2_cmp5_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb2_cmp5_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb2_cmp5_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb2_cmp5_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb2_cmp5),
	.data_out(rnode_2to3_bb2_cmp5_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb2_cmp5_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb2_cmp5_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb2_cmp5_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb2_cmp5_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_2to3_bb2_cmp5_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb2_cmp5_valid_out;
assign local_bb2_cmp5_stall_in = rnode_2to3_bb2_cmp5_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_cmp5_0_NO_SHIFT_REG = rnode_2to3_bb2_cmp5_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_cmp5_0_stall_in_reg_3_NO_SHIFT_REG = rnode_2to3_bb2_cmp5_0_stall_in_NO_SHIFT_REG;
assign rnode_2to3_bb2_cmp5_0_valid_out_NO_SHIFT_REG = rnode_2to3_bb2_cmp5_0_valid_out_reg_3_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx_stall_local;
wire [63:0] local_bb2_arrayidx;

assign local_bb2_arrayidx = ((input_in & 64'hFFFFFFFFFFFFFC00) + ((local_bb2_idxprom & 64'hFFFFFFFF) << 6'h2));

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx_valid_out;
wire local_bb2_arrayidx_stall_in;
wire local_bb2__idxprom_valid_out;
wire local_bb2__idxprom_stall_in;
wire local_bb2__idxprom_inputs_ready;
wire local_bb2__idxprom_stall_local;
 reg [63:0] ffwd_6_0_reg_NO_SHIFT_REG;
 reg local_bb2_arrayidx_consumed_0_NO_SHIFT_REG;
 reg local_bb2__idxprom_consumed_0_NO_SHIFT_REG;

assign local_bb2__idxprom_inputs_ready = rnode_1to2_bb2_add_0_valid_out_NO_SHIFT_REG;
assign ffwd_6_0 = ffwd_6_0_reg_NO_SHIFT_REG;
assign local_bb2__idxprom_stall_local = ((local_bb2_arrayidx_stall_in & ~(local_bb2_arrayidx_consumed_0_NO_SHIFT_REG)) | (local_bb2__idxprom_stall_in & ~(local_bb2__idxprom_consumed_0_NO_SHIFT_REG)));
assign local_bb2_arrayidx_valid_out = (local_bb2__idxprom_inputs_ready & ~(local_bb2_arrayidx_consumed_0_NO_SHIFT_REG));
assign local_bb2__idxprom_valid_out = (local_bb2__idxprom_inputs_ready & ~(local_bb2__idxprom_consumed_0_NO_SHIFT_REG));
assign rnode_1to2_bb2_add_0_stall_in_NO_SHIFT_REG = (|local_bb2__idxprom_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2__idxprom_inputs_ready))
	begin
		ffwd_6_0_reg_NO_SHIFT_REG <= (local_bb2_idxprom & 64'hFFFFFFFF);
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_arrayidx_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__idxprom_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_arrayidx_consumed_0_NO_SHIFT_REG <= (local_bb2__idxprom_inputs_ready & (local_bb2_arrayidx_consumed_0_NO_SHIFT_REG | ~(local_bb2_arrayidx_stall_in)) & local_bb2__idxprom_stall_local);
		local_bb2__idxprom_consumed_0_NO_SHIFT_REG <= (local_bb2__idxprom_inputs_ready & (local_bb2__idxprom_consumed_0_NO_SHIFT_REG | ~(local_bb2__idxprom_stall_in)) & local_bb2__idxprom_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__u5_stall_local;
wire local_bb2_var__u5;

assign local_bb2_var__u5 = (local_bb2_cmp4_acl_ffwd_dest_i1_1 & rnode_2to3_bb2_cmp5_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb2_arrayidx_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb2_arrayidx_0_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb2_arrayidx_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb2_arrayidx_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb2_arrayidx_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb2_arrayidx_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb2_arrayidx_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb2_arrayidx_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb2_arrayidx_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in((local_bb2_arrayidx & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_2to3_bb2_arrayidx_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.DEPTH = 2;
defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.DATA_WIDTH = 64;
defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_2to3_bb2_arrayidx_0_reg_3_fifo.IMPL = "ll_reg";

assign rnode_2to3_bb2_arrayidx_0_reg_3_inputs_ready_NO_SHIFT_REG = local_bb2_arrayidx_valid_out;
assign local_bb2_arrayidx_stall_in = rnode_2to3_bb2_arrayidx_0_stall_out_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx_0_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx_0_stall_in_reg_3_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx_0_stall_in_NO_SHIFT_REG;
assign rnode_2to3_bb2_arrayidx_0_valid_out_NO_SHIFT_REG = rnode_2to3_bb2_arrayidx_0_valid_out_reg_3_NO_SHIFT_REG;

// Register node:
//  * latency = 163
//  * capacity = 163
 logic rcnode_2to165_rc0_bb2___0_valid_out_NO_SHIFT_REG;
 logic rcnode_2to165_rc0_bb2___0_stall_in_NO_SHIFT_REG;
 logic rcnode_2to165_rc0_bb2___0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rcnode_2to165_rc0_bb2___0_valid_out_reg_165_NO_SHIFT_REG;
 logic rcnode_2to165_rc0_bb2___0_stall_in_reg_165_NO_SHIFT_REG;
 logic rcnode_2to165_rc0_bb2___0_stall_out_0_reg_165_IP_NO_SHIFT_REG;
 logic rcnode_2to165_rc0_bb2___0_stall_out_0_reg_165_NO_SHIFT_REG;

acl_data_fifo rcnode_2to165_rc0_bb2___0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_2to165_rc0_bb2___0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_2to165_rc0_bb2___0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rcnode_2to165_rc0_bb2___0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rcnode_2to165_rc0_bb2___0_stall_out_0_reg_165_IP_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rcnode_2to165_rc0_bb2___0_reg_165_fifo.DEPTH = 164;
defparam rcnode_2to165_rc0_bb2___0_reg_165_fifo.DATA_WIDTH = 0;
defparam rcnode_2to165_rc0_bb2___0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_2to165_rc0_bb2___0_reg_165_fifo.IMPL = "ram";

assign rcnode_2to165_rc0_bb2___0_reg_165_inputs_ready_NO_SHIFT_REG = (local_bb2___valid_out & local_bb2__idxprom_valid_out);
assign rcnode_2to165_rc0_bb2___0_stall_out_0_reg_165_NO_SHIFT_REG = (~(rcnode_2to165_rc0_bb2___0_reg_165_inputs_ready_NO_SHIFT_REG) | rcnode_2to165_rc0_bb2___0_stall_out_0_reg_165_IP_NO_SHIFT_REG);
assign local_bb2___stall_in = rcnode_2to165_rc0_bb2___0_stall_out_0_reg_165_NO_SHIFT_REG;
assign local_bb2__idxprom_stall_in = rcnode_2to165_rc0_bb2___0_stall_out_0_reg_165_NO_SHIFT_REG;
assign rcnode_2to165_rc0_bb2___0_stall_in_reg_165_NO_SHIFT_REG = rcnode_2to165_rc0_bb2___0_stall_in_NO_SHIFT_REG;
assign rcnode_2to165_rc0_bb2___0_valid_out_NO_SHIFT_REG = rcnode_2to165_rc0_bb2___0_valid_out_reg_165_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__phi_decision_xor_stall_local;
wire local_bb2__phi_decision_xor;

assign local_bb2__phi_decision_xor = (local_bb2_var__u5 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__phi_decision_xor_valid_out;
wire local_bb2__phi_decision_xor_stall_in;
wire local_bb2___u6_valid_out;
wire local_bb2___u6_stall_in;
wire local_bb2___u6_inputs_ready;
wire local_bb2___u6_stall_local;
 reg ffwd_5_0_reg_NO_SHIFT_REG;
 reg local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG;
 reg local_bb2___u6_consumed_0_NO_SHIFT_REG;

assign local_bb2___u6_inputs_ready = (rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb2_cmp5_0_valid_out_NO_SHIFT_REG);
assign ffwd_5_0 = ffwd_5_0_reg_NO_SHIFT_REG;
assign local_bb2___u6_stall_local = ((local_bb2__phi_decision_xor_stall_in & ~(local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG)) | (local_bb2___u6_stall_in & ~(local_bb2___u6_consumed_0_NO_SHIFT_REG)));
assign local_bb2__phi_decision_xor_valid_out = (local_bb2___u6_inputs_ready & ~(local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG));
assign local_bb2___u6_valid_out = (local_bb2___u6_inputs_ready & ~(local_bb2___u6_consumed_0_NO_SHIFT_REG));
assign rnode_1to3_bb2_cmp4_acl_ffwd_dest_i1_1_0_stall_in_NO_SHIFT_REG = (local_bb2___u6_stall_local | ~(local_bb2___u6_inputs_ready));
assign rnode_2to3_bb2_cmp5_0_stall_in_NO_SHIFT_REG = (local_bb2___u6_stall_local | ~(local_bb2___u6_inputs_ready));

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___u6_inputs_ready))
	begin
		ffwd_5_0_reg_NO_SHIFT_REG <= local_bb2_var__u5;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2___u6_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= (local_bb2___u6_inputs_ready & (local_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG | ~(local_bb2__phi_decision_xor_stall_in)) & local_bb2___u6_stall_local);
		local_bb2___u6_consumed_0_NO_SHIFT_REG <= (local_bb2___u6_inputs_ready & (local_bb2___u6_consumed_0_NO_SHIFT_REG | ~(local_bb2___u6_stall_in)) & local_bb2___u6_stall_local);
	end
end


// This section implements a staging register.
// 
wire rstag_3to3_bb2__phi_decision_xor_valid_out_0;
wire rstag_3to3_bb2__phi_decision_xor_stall_in_0;
wire rstag_3to3_bb2__phi_decision_xor_valid_out_1;
wire rstag_3to3_bb2__phi_decision_xor_stall_in_1;
wire rstag_3to3_bb2__phi_decision_xor_inputs_ready;
wire rstag_3to3_bb2__phi_decision_xor_stall_local;
 reg rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG;
wire rstag_3to3_bb2__phi_decision_xor_combined_valid;
 reg rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG;
wire rstag_3to3_bb2__phi_decision_xor;
 reg rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG;
 reg rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG;

assign rstag_3to3_bb2__phi_decision_xor_inputs_ready = local_bb2__phi_decision_xor_valid_out;
assign rstag_3to3_bb2__phi_decision_xor = (rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG ? rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG : local_bb2__phi_decision_xor);
assign rstag_3to3_bb2__phi_decision_xor_combined_valid = (rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG | rstag_3to3_bb2__phi_decision_xor_inputs_ready);
assign rstag_3to3_bb2__phi_decision_xor_stall_local = ((rstag_3to3_bb2__phi_decision_xor_stall_in_0 & ~(rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG)) | (rstag_3to3_bb2__phi_decision_xor_stall_in_1 & ~(rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG)));
assign rstag_3to3_bb2__phi_decision_xor_valid_out_0 = (rstag_3to3_bb2__phi_decision_xor_combined_valid & ~(rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG));
assign rstag_3to3_bb2__phi_decision_xor_valid_out_1 = (rstag_3to3_bb2__phi_decision_xor_combined_valid & ~(rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG));
assign local_bb2__phi_decision_xor_stall_in = (|rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_3to3_bb2__phi_decision_xor_stall_local)
		begin
			if (~(rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG))
			begin
				rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG <= rstag_3to3_bb2__phi_decision_xor_inputs_ready;
			end
		end
		else
		begin
			rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_3to3_bb2__phi_decision_xor_staging_valid_NO_SHIFT_REG))
		begin
			rstag_3to3_bb2__phi_decision_xor_staging_reg_NO_SHIFT_REG <= local_bb2__phi_decision_xor;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG <= (rstag_3to3_bb2__phi_decision_xor_combined_valid & (rstag_3to3_bb2__phi_decision_xor_consumed_0_NO_SHIFT_REG | ~(rstag_3to3_bb2__phi_decision_xor_stall_in_0)) & rstag_3to3_bb2__phi_decision_xor_stall_local);
		rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG <= (rstag_3to3_bb2__phi_decision_xor_combined_valid & (rstag_3to3_bb2__phi_decision_xor_consumed_1_NO_SHIFT_REG | ~(rstag_3to3_bb2__phi_decision_xor_stall_in_1)) & rstag_3to3_bb2__phi_decision_xor_stall_local);
	end
end


// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_3to165_bb2___u6_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u6_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u6_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u6_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u6_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2___u6_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_3to165_bb2___u6_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to165_bb2___u6_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to165_bb2___u6_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_3to165_bb2___u6_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_3to165_bb2___u6_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to165_bb2___u6_0_reg_165_fifo.DEPTH = 163;
defparam rnode_3to165_bb2___u6_0_reg_165_fifo.DATA_WIDTH = 0;
defparam rnode_3to165_bb2___u6_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_3to165_bb2___u6_0_reg_165_fifo.IMPL = "ram";

assign rnode_3to165_bb2___u6_0_reg_165_inputs_ready_NO_SHIFT_REG = local_bb2___u6_valid_out;
assign local_bb2___u6_stall_in = rnode_3to165_bb2___u6_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_3to165_bb2___u6_0_stall_in_reg_165_NO_SHIFT_REG = rnode_3to165_bb2___u6_0_stall_in_NO_SHIFT_REG;
assign rnode_3to165_bb2___u6_0_valid_out_NO_SHIFT_REG = rnode_3to165_bb2___u6_0_valid_out_reg_165_NO_SHIFT_REG;

// Register node:
//  * latency = 162
//  * capacity = 162
 logic rnode_3to165_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_3to165_bb2__phi_decision_xor_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to165_bb2__phi_decision_xor_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to165_bb2__phi_decision_xor_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_3to165_bb2__phi_decision_xor_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_3to165_bb2__phi_decision_xor_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(rstag_3to3_bb2__phi_decision_xor),
	.data_out(rnode_3to165_bb2__phi_decision_xor_0_reg_165_NO_SHIFT_REG)
);

defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.DEPTH = 163;
defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.DATA_WIDTH = 1;
defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_3to165_bb2__phi_decision_xor_0_reg_165_fifo.IMPL = "ram";

assign rnode_3to165_bb2__phi_decision_xor_0_reg_165_inputs_ready_NO_SHIFT_REG = rstag_3to3_bb2__phi_decision_xor_valid_out_0;
assign rstag_3to3_bb2__phi_decision_xor_stall_in_0 = rnode_3to165_bb2__phi_decision_xor_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_reg_165_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_stall_in_reg_165_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_valid_out_reg_165_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb2_ld__inputs_ready;
 reg local_bb2_ld__valid_out_NO_SHIFT_REG;
wire local_bb2_ld__stall_in;
wire local_bb2_ld__output_regs_ready;
wire local_bb2_ld__fu_stall_out;
wire local_bb2_ld__fu_valid_out;
wire [31:0] local_bb2_ld__lsu_dataout;
 reg [31:0] local_bb2_ld__NO_SHIFT_REG;
wire local_bb2_ld__causedstall;

lsu_top lsu_local_bb2_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld__fu_stall_out),
	.i_valid(local_bb2_ld__inputs_ready),
	.i_address((rnode_2to3_bb2_arrayidx_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_3to3_bb2__phi_decision_xor),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld__output_regs_ready)),
	.o_valid(local_bb2_ld__fu_valid_out),
	.o_readdata(local_bb2_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld__active),
	.avm_address(avm_local_bb2_ld__address),
	.avm_read(avm_local_bb2_ld__read),
	.avm_readdata(avm_local_bb2_ld__readdata),
	.avm_write(avm_local_bb2_ld__write),
	.avm_writeack(avm_local_bb2_ld__writeack),
	.avm_burstcount(avm_local_bb2_ld__burstcount),
	.avm_writedata(avm_local_bb2_ld__writedata),
	.avm_byteenable(avm_local_bb2_ld__byteenable),
	.avm_waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld_.AWIDTH = 33;
defparam lsu_local_bb2_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb2_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb2_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb2_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld_.READ = 1;
defparam lsu_local_bb2_ld_.ATOMIC = 0;
defparam lsu_local_bb2_ld_.WIDTH = 32;
defparam lsu_local_bb2_ld_.MWIDTH = 512;
defparam lsu_local_bb2_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld_.MEMORY_SIDE_MEM_LATENCY = 115;
defparam lsu_local_bb2_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb2_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld_.USECACHING = 0;
defparam lsu_local_bb2_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld_.ADDRSPACE = 1;
defparam lsu_local_bb2_ld_.STYLE = "BURST-COALESCED";

assign local_bb2_ld__inputs_ready = (rnode_2to3_bb2_arrayidx_0_valid_out_NO_SHIFT_REG & rstag_3to3_bb2__phi_decision_xor_valid_out_1);
assign local_bb2_ld__output_regs_ready = (&(~(local_bb2_ld__valid_out_NO_SHIFT_REG) | ~(local_bb2_ld__stall_in)));
assign rnode_2to3_bb2_arrayidx_0_stall_in_NO_SHIFT_REG = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign rstag_3to3_bb2__phi_decision_xor_stall_in_1 = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign local_bb2_ld__causedstall = (local_bb2_ld__inputs_ready && (local_bb2_ld__fu_stall_out && !(~(local_bb2_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld__NO_SHIFT_REG <= 'x;
		local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld__output_regs_ready)
		begin
			local_bb2_ld__NO_SHIFT_REG <= local_bb2_ld__lsu_dataout;
			local_bb2_ld__valid_out_NO_SHIFT_REG <= local_bb2_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld__stall_in))
			begin
				local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_165to166_rc0_bb2__indvars_iv39_0_valid_out_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_in_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv39_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_IP_NO_SHIFT_REG;
 logic rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_NO_SHIFT_REG;

acl_data_fifo rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rcnode_165to166_rc0_bb2__indvars_iv39_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_IP_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_fifo.DEPTH = 1;
defparam rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_fifo.DATA_WIDTH = 0;
defparam rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_fifo.IMPL = "ll_reg";

assign rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_inputs_ready_NO_SHIFT_REG = (rnode_1to165_bb2__indvars_iv39_0_valid_out_NO_SHIFT_REG & rnode_3to165_bb2___u6_0_valid_out_NO_SHIFT_REG & rcnode_2to165_rc0_bb2___0_valid_out_NO_SHIFT_REG);
assign rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_NO_SHIFT_REG = (~(rcnode_165to166_rc0_bb2__indvars_iv39_0_reg_166_inputs_ready_NO_SHIFT_REG) | rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_IP_NO_SHIFT_REG);
assign rnode_1to165_bb2__indvars_iv39_0_stall_in_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rnode_3to165_bb2___u6_0_stall_in_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_2to165_rc0_bb2___0_stall_in_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_out_0_reg_166_NO_SHIFT_REG;
assign rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_in_reg_166_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_in_NO_SHIFT_REG;
assign rcnode_165to166_rc0_bb2__indvars_iv39_0_valid_out_NO_SHIFT_REG = rcnode_165to166_rc0_bb2__indvars_iv39_0_valid_out_reg_166_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_reg_166_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rnode_165to166_bb2__phi_decision_xor_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_165to166_bb2__phi_decision_xor_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_165to166_bb2__phi_decision_xor_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_165to166_bb2__phi_decision_xor_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_165to166_bb2__phi_decision_xor_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(rnode_3to165_bb2__phi_decision_xor_0_NO_SHIFT_REG),
	.data_out(rnode_165to166_bb2__phi_decision_xor_0_reg_166_NO_SHIFT_REG)
);

defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.DEPTH = 1;
defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.DATA_WIDTH = 1;
defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_165to166_bb2__phi_decision_xor_0_reg_166_fifo.IMPL = "ll_reg";

assign rnode_165to166_bb2__phi_decision_xor_0_reg_166_inputs_ready_NO_SHIFT_REG = rnode_3to165_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG;
assign rnode_3to165_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_165to166_bb2__phi_decision_xor_0_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_reg_166_NO_SHIFT_REG;
assign rnode_165to166_bb2__phi_decision_xor_0_stall_in_reg_166_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG;
assign rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG = rnode_165to166_bb2__phi_decision_xor_0_valid_out_reg_166_NO_SHIFT_REG;

// This section implements a staging register.
// 
wire rstag_163to163_bb2_ld__valid_out_0;
wire rstag_163to163_bb2_ld__stall_in_0;
wire rstag_163to163_bb2_ld__valid_out_1;
wire rstag_163to163_bb2_ld__stall_in_1;
wire rstag_163to163_bb2_ld__inputs_ready;
wire rstag_163to163_bb2_ld__stall_local;
 reg rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG;
wire rstag_163to163_bb2_ld__combined_valid;
 reg [31:0] rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_163to163_bb2_ld_;
 reg rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG;
 reg rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG;

assign rstag_163to163_bb2_ld__inputs_ready = local_bb2_ld__valid_out_NO_SHIFT_REG;
assign rstag_163to163_bb2_ld_ = (rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG ? rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG : local_bb2_ld__NO_SHIFT_REG);
assign rstag_163to163_bb2_ld__combined_valid = (rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG | rstag_163to163_bb2_ld__inputs_ready);
assign rstag_163to163_bb2_ld__stall_local = ((rstag_163to163_bb2_ld__stall_in_0 & ~(rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG)) | (rstag_163to163_bb2_ld__stall_in_1 & ~(rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG)));
assign rstag_163to163_bb2_ld__valid_out_0 = (rstag_163to163_bb2_ld__combined_valid & ~(rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG));
assign rstag_163to163_bb2_ld__valid_out_1 = (rstag_163to163_bb2_ld__combined_valid & ~(rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG));
assign local_bb2_ld__stall_in = (|rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_163to163_bb2_ld__stall_local)
		begin
			if (~(rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG <= rstag_163to163_bb2_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_163to163_bb2_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_163to163_bb2_ld__staging_reg_NO_SHIFT_REG <= local_bb2_ld__NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG <= (rstag_163to163_bb2_ld__combined_valid & (rstag_163to163_bb2_ld__consumed_0_NO_SHIFT_REG | ~(rstag_163to163_bb2_ld__stall_in_0)) & rstag_163to163_bb2_ld__stall_local);
		rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG <= (rstag_163to163_bb2_ld__combined_valid & (rstag_163to163_bb2_ld__consumed_1_NO_SHIFT_REG | ~(rstag_163to163_bb2_ld__stall_in_1)) & rstag_163to163_bb2_ld__stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2___u7_valid_out;
wire local_bb2___u7_stall_in;
wire local_bb2___u7_inputs_ready;
wire local_bb2___u7_stall_local;
 reg [31:0] ffwd_7_0_reg_NO_SHIFT_REG;

assign local_bb2___u7_inputs_ready = rstag_163to163_bb2_ld__valid_out_0;
assign ffwd_7_0 = ffwd_7_0_reg_NO_SHIFT_REG;
assign local_bb2___u7_valid_out = local_bb2___u7_inputs_ready;
assign local_bb2___u7_stall_local = local_bb2___u7_stall_in;
assign rstag_163to163_bb2_ld__stall_in_0 = (|local_bb2___u7_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___u7_inputs_ready))
	begin
		ffwd_7_0_reg_NO_SHIFT_REG <= rstag_163to163_bb2_ld_;
	end
end


// This section implements a registered operation.
// 
wire local_bb2_cmp8_inputs_ready;
 reg local_bb2_cmp8_valid_out_NO_SHIFT_REG;
wire local_bb2_cmp8_stall_in;
wire local_bb2_cmp8_output_regs_ready;
wire local_bb2_cmp8;
 reg local_bb2_cmp8_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_cmp8_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_cmp8_causedstall;

acl_fp_cmp fp_module_local_bb2_cmp8 (
	.clock(clock),
	.dataa(rstag_163to163_bb2_ld_),
	.datab(32'h0),
	.enable(local_bb2_cmp8_output_regs_ready),
	.result(local_bb2_cmp8)
);

defparam fp_module_local_bb2_cmp8.COMPARISON_MODE = 0;

assign local_bb2_cmp8_inputs_ready = rstag_163to163_bb2_ld__valid_out_1;
assign local_bb2_cmp8_output_regs_ready = (&(~(local_bb2_cmp8_valid_out_NO_SHIFT_REG) | ~(local_bb2_cmp8_stall_in)));
assign rstag_163to163_bb2_ld__stall_in_1 = (~(local_bb2_cmp8_output_regs_ready) | ~(local_bb2_cmp8_inputs_ready));
assign local_bb2_cmp8_causedstall = (local_bb2_cmp8_inputs_ready && (~(local_bb2_cmp8_output_regs_ready) && !(~(local_bb2_cmp8_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp8_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp8_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_cmp8_output_regs_ready)
		begin
			local_bb2_cmp8_valid_pipe_0_NO_SHIFT_REG <= local_bb2_cmp8_inputs_ready;
			local_bb2_cmp8_valid_pipe_1_NO_SHIFT_REG <= local_bb2_cmp8_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp8_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_cmp8_output_regs_ready)
		begin
			local_bb2_cmp8_valid_out_NO_SHIFT_REG <= local_bb2_cmp8_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb2_cmp8_stall_in))
			begin
				local_bb2_cmp8_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_163to166_bb2___u7_0_valid_out_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u7_0_stall_in_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u7_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u7_0_valid_out_reg_166_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u7_0_stall_in_reg_166_NO_SHIFT_REG;
 logic rnode_163to166_bb2___u7_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_163to166_bb2___u7_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_163to166_bb2___u7_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_163to166_bb2___u7_0_stall_in_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_163to166_bb2___u7_0_valid_out_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_163to166_bb2___u7_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_163to166_bb2___u7_0_reg_166_fifo.DEPTH = 4;
defparam rnode_163to166_bb2___u7_0_reg_166_fifo.DATA_WIDTH = 0;
defparam rnode_163to166_bb2___u7_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_163to166_bb2___u7_0_reg_166_fifo.IMPL = "ll_reg";

assign rnode_163to166_bb2___u7_0_reg_166_inputs_ready_NO_SHIFT_REG = local_bb2___u7_valid_out;
assign local_bb2___u7_stall_in = rnode_163to166_bb2___u7_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_163to166_bb2___u7_0_stall_in_reg_166_NO_SHIFT_REG = rnode_163to166_bb2___u7_0_stall_in_NO_SHIFT_REG;
assign rnode_163to166_bb2___u7_0_valid_out_NO_SHIFT_REG = rnode_163to166_bb2___u7_0_valid_out_reg_166_NO_SHIFT_REG;

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_166to166_bb2_cmp8_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_1_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_reg_166_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_reg_166_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_valid_out_0_reg_166_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_stall_in_0_reg_166_NO_SHIFT_REG;
 logic rnode_166to166_bb2_cmp8_0_stall_out_reg_166_NO_SHIFT_REG;

acl_data_fifo rnode_166to166_bb2_cmp8_0_reg_166_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to166_bb2_cmp8_0_reg_166_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to166_bb2_cmp8_0_stall_in_0_reg_166_NO_SHIFT_REG),
	.valid_out(rnode_166to166_bb2_cmp8_0_valid_out_0_reg_166_NO_SHIFT_REG),
	.stall_out(rnode_166to166_bb2_cmp8_0_stall_out_reg_166_NO_SHIFT_REG),
	.data_in(local_bb2_cmp8),
	.data_out(rnode_166to166_bb2_cmp8_0_reg_166_NO_SHIFT_REG)
);

defparam rnode_166to166_bb2_cmp8_0_reg_166_fifo.DEPTH = 3;
defparam rnode_166to166_bb2_cmp8_0_reg_166_fifo.DATA_WIDTH = 1;
defparam rnode_166to166_bb2_cmp8_0_reg_166_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_166to166_bb2_cmp8_0_reg_166_fifo.IMPL = "zl_reg";

assign rnode_166to166_bb2_cmp8_0_reg_166_inputs_ready_NO_SHIFT_REG = local_bb2_cmp8_valid_out_NO_SHIFT_REG;
assign local_bb2_cmp8_stall_in = rnode_166to166_bb2_cmp8_0_stall_out_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp8_0_stall_in_0_reg_166_NO_SHIFT_REG = (rnode_166to166_bb2_cmp8_0_stall_in_0_NO_SHIFT_REG | rnode_166to166_bb2_cmp8_0_stall_in_1_NO_SHIFT_REG);
assign rnode_166to166_bb2_cmp8_0_valid_out_0_NO_SHIFT_REG = rnode_166to166_bb2_cmp8_0_valid_out_0_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp8_0_valid_out_1_NO_SHIFT_REG = rnode_166to166_bb2_cmp8_0_valid_out_0_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp8_0_NO_SHIFT_REG = rnode_166to166_bb2_cmp8_0_reg_166_NO_SHIFT_REG;
assign rnode_166to166_bb2_cmp8_1_NO_SHIFT_REG = rnode_166to166_bb2_cmp8_0_reg_166_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__cmp8_stall_local;
 reg ffwd_8_0_reg_NO_SHIFT_REG;
wire local_bb2__cmp8_inputs_ready;

assign ffwd_8_0 = ffwd_8_0_reg_NO_SHIFT_REG;

always @(posedge clock)
begin
	if ((1'b1 & local_bb2__cmp8_inputs_ready))
	begin
		ffwd_8_0_reg_NO_SHIFT_REG <= rnode_166to166_bb2_cmp8_0_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_var__u8_stall_local;
wire local_bb2_var__u8;

assign local_bb2_var__u8 = (rnode_166to166_bb2_cmp8_1_NO_SHIFT_REG | rnode_165to166_bb2__phi_decision_xor_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u9_stall_local;
wire local_bb2_var__u9;

assign local_bb2_var__u9 = (local_bb2_var__u8 | input_wii_cmp1526);

// This section implements an unregistered operation.
// 
wire local_bb2___u10_valid_out;
wire local_bb2___u10_stall_in;
wire local_bb2__cmp8_valid_out;
wire local_bb2__cmp8_stall_in;
wire local_bb2___u10_inputs_ready;
wire local_bb2___u10_stall_local;
 reg ffwd_9_0_reg_NO_SHIFT_REG;

assign local_bb2___u10_inputs_ready = (rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG & rnode_166to166_bb2_cmp8_0_valid_out_1_NO_SHIFT_REG & rnode_166to166_bb2_cmp8_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__cmp8_inputs_ready = (rnode_165to166_bb2__phi_decision_xor_0_valid_out_NO_SHIFT_REG & rnode_166to166_bb2_cmp8_0_valid_out_1_NO_SHIFT_REG & rnode_166to166_bb2_cmp8_0_valid_out_0_NO_SHIFT_REG);
assign ffwd_9_0 = ffwd_9_0_reg_NO_SHIFT_REG;
assign local_bb2___u10_stall_local = (local_bb2___u10_stall_in | local_bb2__cmp8_stall_in);
assign local_bb2___u10_valid_out = local_bb2___u10_inputs_ready;
assign local_bb2__cmp8_valid_out = local_bb2___u10_inputs_ready;
assign rnode_165to166_bb2__phi_decision_xor_0_stall_in_NO_SHIFT_REG = (local_bb2___u10_stall_local | ~(local_bb2___u10_inputs_ready));
assign rnode_166to166_bb2_cmp8_0_stall_in_1_NO_SHIFT_REG = (local_bb2___u10_stall_local | ~(local_bb2___u10_inputs_ready));
assign rnode_166to166_bb2_cmp8_0_stall_in_0_NO_SHIFT_REG = (local_bb2___u10_stall_local | ~(local_bb2___u10_inputs_ready));

always @(posedge clock)
begin
	if ((1'b1 & local_bb2___u10_inputs_ready))
	begin
		ffwd_9_0_reg_NO_SHIFT_REG <= local_bb2_var__u9;
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;

assign branch_var__inputs_ready = (local_bb2___u10_valid_out & local_bb2__cmp8_valid_out & rnode_163to166_bb2___u7_0_valid_out_NO_SHIFT_REG & rcnode_165to166_rc0_bb2__indvars_iv39_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb2___u10_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb2__cmp8_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_163to166_bb2___u7_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_165to166_rc0_bb2__indvars_iv39_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_3
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_r,
		input 		input_wii_cmp1526,
		input [31:0] 		input_wii_sub24,
		input [31:0] 		input_wii_sub27,
		input [31:0] 		input_wii_mul48,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u11,
		input 		valid_in_0,
		output 		stall_out_0,
		input 		input_forked_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input 		input_forked_1,
		output 		valid_out,
		input 		stall_in,
		output [31:0] 		lvb_bb3_c0_exe1,
		output [31:0] 		lvb_bb3_c0_exe2,
		output 		lvb_bb3_c0_exe3,
		output 		lvb_bb3_c0_exe4,
		output [31:0] 		lvb_bb3_t_228_pop5_,
		output [31:0] 		lvb_bb3_sum_227_pop6_,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		feedback_valid_in_5,
		output 		feedback_stall_out_5,
		input [31:0] 		feedback_data_in_5,
		input 		feedback_valid_in_6,
		output 		feedback_stall_out_6,
		input [31:0] 		feedback_data_in_6,
		input 		feedback_valid_in_4,
		output 		feedback_stall_out_4,
		input [63:0] 		feedback_data_in_4,
		input 		ffwd_9_0,
		output 		feedback_stall_out_2,
		input 		feedback_valid_in_3,
		output 		feedback_stall_out_3,
		input 		feedback_data_in_3,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		input [31:0] 		ffwd_4_0,
		output 		feedback_valid_out_3,
		input 		feedback_stall_in_3,
		output 		feedback_data_out_3,
		output 		feedback_valid_out_4,
		input 		feedback_stall_in_4,
		output [63:0] 		feedback_data_out_4
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg input_forked_0_staging_reg_NO_SHIFT_REG;
 reg local_lvm_forked_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg input_forked_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_forked_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_forked_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_forked_0_staging_reg_NO_SHIFT_REG <= input_forked_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_forked_1_staging_reg_NO_SHIFT_REG <= input_forked_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_forked_NO_SHIFT_REG <= input_forked_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_eni1_stall_local;
wire [15:0] local_bb3_c0_eni1;

assign local_bb3_c0_eni1[7:0] = 8'bx;
assign local_bb3_c0_eni1[8] = local_lvm_forked_NO_SHIFT_REG;
assign local_bb3_c0_eni1[15:9] = 7'bx;

// Register node:
//  * latency = 8
//  * capacity = 8
 logic rnode_1to9_forked_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to9_forked_1_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_reg_9_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG;
 logic rnode_1to9_forked_0_stall_out_reg_9_NO_SHIFT_REG;
 reg rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG;
 reg rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_1to9_forked_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to9_forked_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_1to9_forked_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(local_lvm_forked_NO_SHIFT_REG),
	.data_out(rnode_1to9_forked_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_1to9_forked_0_reg_9_fifo.DEPTH = 9;
defparam rnode_1to9_forked_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_1to9_forked_0_reg_9_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to9_forked_0_reg_9_fifo.IMPL = "ram_plus_reg";

assign rnode_1to9_forked_0_reg_9_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign merge_node_stall_in_1 = rnode_1to9_forked_0_stall_out_reg_9_NO_SHIFT_REG;
assign rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG = ((rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG)) | (rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG)));
assign rnode_1to9_forked_0_valid_out_0_NO_SHIFT_REG = (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG));
assign rnode_1to9_forked_0_valid_out_1_NO_SHIFT_REG = (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & ~(rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG));
assign rnode_1to9_forked_0_NO_SHIFT_REG = rnode_1to9_forked_0_reg_9_NO_SHIFT_REG;
assign rnode_1to9_forked_1_NO_SHIFT_REG = rnode_1to9_forked_0_reg_9_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG <= (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & (rnode_1to9_forked_0_consumed_0_NO_SHIFT_REG | ~(rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG)) & rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG);
		rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG <= (rnode_1to9_forked_0_valid_out_0_reg_9_NO_SHIFT_REG & (rnode_1to9_forked_0_consumed_1_NO_SHIFT_REG | ~(rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG)) & rnode_1to9_forked_0_stall_in_0_reg_9_NO_SHIFT_REG);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_valid_out_1;
wire local_bb3_c0_ene1_stall_in_1;
wire SFC_1_VALID_1_1_0_valid_out_0;
wire SFC_1_VALID_1_1_0_stall_in_0;
wire local_bb3_indvars_iv35_pop4__valid_out;
wire local_bb3_indvars_iv35_pop4__stall_in;
wire local_bb3_c0_enter_c0_eni1_inputs_ready;
wire local_bb3_c0_enter_c0_eni1_stall_local;
wire local_bb3_c0_enter_c0_eni1_input_accepted;
wire [15:0] local_bb3_c0_enter_c0_eni1;
wire local_bb3_c0_exit_c0_exi4_entry_stall;
wire local_bb3_c0_enter_c0_eni1_valid_bit;
wire local_bb3_c0_exit_c0_exi4_output_regs_ready;
wire local_bb3_c0_exit_c0_exi4_valid_in;
wire local_bb3_c0_exit_c0_exi4_phases;
wire local_bb3_c0_enter_c0_eni1_inc_pipelined_thread;
wire local_bb3_c0_enter_c0_eni1_dec_pipelined_thread;
wire local_bb3_c0_enter_c0_eni1_fu_stall_out;

assign local_bb3_c0_enter_c0_eni1_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb3_c0_enter_c0_eni1 = local_bb3_c0_eni1;
assign local_bb3_c0_enter_c0_eni1_input_accepted = (local_bb3_c0_enter_c0_eni1_inputs_ready && !(local_bb3_c0_exit_c0_exi4_entry_stall));
assign local_bb3_c0_enter_c0_eni1_valid_bit = local_bb3_c0_enter_c0_eni1_input_accepted;
assign local_bb3_c0_enter_c0_eni1_inc_pipelined_thread = 1'b1;
assign local_bb3_c0_enter_c0_eni1_dec_pipelined_thread = ~(1'b0);
assign local_bb3_c0_enter_c0_eni1_fu_stall_out = (~(local_bb3_c0_enter_c0_eni1_inputs_ready) | local_bb3_c0_exit_c0_exi4_entry_stall);
assign local_bb3_c0_enter_c0_eni1_stall_local = (local_bb3_c0_ene1_stall_in_1 | SFC_1_VALID_1_1_0_stall_in_0 | local_bb3_indvars_iv35_pop4__stall_in);
assign local_bb3_c0_ene1_valid_out_1 = local_bb3_c0_enter_c0_eni1_inputs_ready;
assign SFC_1_VALID_1_1_0_valid_out_0 = local_bb3_c0_enter_c0_eni1_inputs_ready;
assign local_bb3_indvars_iv35_pop4__valid_out = local_bb3_c0_enter_c0_eni1_inputs_ready;
assign merge_node_stall_in_0 = (|local_bb3_c0_enter_c0_eni1_fu_stall_out);

// This section implements a registered operation.
// 
wire local_bb3_t_228_pop5__inputs_ready;
 reg local_bb3_t_228_pop5__valid_out_NO_SHIFT_REG;
wire local_bb3_t_228_pop5__stall_in;
wire local_bb3_t_228_pop5__output_regs_ready;
wire [31:0] local_bb3_t_228_pop5__result;
wire local_bb3_t_228_pop5__fu_valid_out;
wire local_bb3_t_228_pop5__fu_stall_out;
 reg [31:0] local_bb3_t_228_pop5__NO_SHIFT_REG;
wire local_bb3_t_228_pop5__causedstall;

acl_pop local_bb3_t_228_pop5__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to9_forked_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(32'h0),
	.stall_out(local_bb3_t_228_pop5__fu_stall_out),
	.valid_in(local_bb3_t_228_pop5__inputs_ready),
	.valid_out(local_bb3_t_228_pop5__fu_valid_out),
	.stall_in(~(local_bb3_t_228_pop5__output_regs_ready)),
	.data_out(local_bb3_t_228_pop5__result),
	.feedback_in(feedback_data_in_5),
	.feedback_valid_in(feedback_valid_in_5),
	.feedback_stall_out(feedback_stall_out_5)
);

defparam local_bb3_t_228_pop5__feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_t_228_pop5__feedback.DATA_WIDTH = 32;
defparam local_bb3_t_228_pop5__feedback.STYLE = "REGULAR";

assign local_bb3_t_228_pop5__inputs_ready = rnode_1to9_forked_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_t_228_pop5__output_regs_ready = (&(~(local_bb3_t_228_pop5__valid_out_NO_SHIFT_REG) | ~(local_bb3_t_228_pop5__stall_in)));
assign rnode_1to9_forked_0_stall_in_0_NO_SHIFT_REG = (local_bb3_t_228_pop5__fu_stall_out | ~(local_bb3_t_228_pop5__inputs_ready));
assign local_bb3_t_228_pop5__causedstall = (local_bb3_t_228_pop5__inputs_ready && (local_bb3_t_228_pop5__fu_stall_out && !(~(local_bb3_t_228_pop5__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_t_228_pop5__NO_SHIFT_REG <= 'x;
		local_bb3_t_228_pop5__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_t_228_pop5__output_regs_ready)
		begin
			local_bb3_t_228_pop5__NO_SHIFT_REG <= local_bb3_t_228_pop5__result;
			local_bb3_t_228_pop5__valid_out_NO_SHIFT_REG <= local_bb3_t_228_pop5__fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_t_228_pop5__stall_in))
			begin
				local_bb3_t_228_pop5__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_sum_227_pop6__inputs_ready;
 reg local_bb3_sum_227_pop6__valid_out_NO_SHIFT_REG;
wire local_bb3_sum_227_pop6__stall_in;
wire local_bb3_sum_227_pop6__output_regs_ready;
wire [31:0] local_bb3_sum_227_pop6__result;
wire local_bb3_sum_227_pop6__fu_valid_out;
wire local_bb3_sum_227_pop6__fu_stall_out;
 reg [31:0] local_bb3_sum_227_pop6__NO_SHIFT_REG;
wire local_bb3_sum_227_pop6__causedstall;

acl_pop local_bb3_sum_227_pop6__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to9_forked_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(32'h0),
	.stall_out(local_bb3_sum_227_pop6__fu_stall_out),
	.valid_in(local_bb3_sum_227_pop6__inputs_ready),
	.valid_out(local_bb3_sum_227_pop6__fu_valid_out),
	.stall_in(~(local_bb3_sum_227_pop6__output_regs_ready)),
	.data_out(local_bb3_sum_227_pop6__result),
	.feedback_in(feedback_data_in_6),
	.feedback_valid_in(feedback_valid_in_6),
	.feedback_stall_out(feedback_stall_out_6)
);

defparam local_bb3_sum_227_pop6__feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_sum_227_pop6__feedback.DATA_WIDTH = 32;
defparam local_bb3_sum_227_pop6__feedback.STYLE = "REGULAR";

assign local_bb3_sum_227_pop6__inputs_ready = rnode_1to9_forked_0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_sum_227_pop6__output_regs_ready = (&(~(local_bb3_sum_227_pop6__valid_out_NO_SHIFT_REG) | ~(local_bb3_sum_227_pop6__stall_in)));
assign rnode_1to9_forked_0_stall_in_1_NO_SHIFT_REG = (local_bb3_sum_227_pop6__fu_stall_out | ~(local_bb3_sum_227_pop6__inputs_ready));
assign local_bb3_sum_227_pop6__causedstall = (local_bb3_sum_227_pop6__inputs_ready && (local_bb3_sum_227_pop6__fu_stall_out && !(~(local_bb3_sum_227_pop6__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_sum_227_pop6__NO_SHIFT_REG <= 'x;
		local_bb3_sum_227_pop6__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_sum_227_pop6__output_regs_ready)
		begin
			local_bb3_sum_227_pop6__NO_SHIFT_REG <= local_bb3_sum_227_pop6__result;
			local_bb3_sum_227_pop6__valid_out_NO_SHIFT_REG <= local_bb3_sum_227_pop6__fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_sum_227_pop6__stall_in))
			begin
				local_bb3_sum_227_pop6__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_ene1_stall_local;
wire local_bb3_c0_ene1;

assign local_bb3_c0_ene1 = local_bb3_c0_enter_c0_eni1[8];

// This section implements an unregistered operation.
// 
wire SFC_1_VALID_1_1_0_stall_local;
wire SFC_1_VALID_1_1_0;

assign SFC_1_VALID_1_1_0 = local_bb3_c0_enter_c0_eni1_valid_bit;

// This section implements an unregistered operation.
// 
wire local_bb3_indvars_iv35_pop4__stall_local;
wire [63:0] local_bb3_indvars_iv35_pop4_;
wire local_bb3_indvars_iv35_pop4__fu_valid_out;
wire local_bb3_indvars_iv35_pop4__fu_stall_out;

acl_pop local_bb3_indvars_iv35_pop4__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_c0_ene1),
	.predicate(1'b0),
	.data_in(input_wii_var_),
	.stall_out(local_bb3_indvars_iv35_pop4__fu_stall_out),
	.valid_in(SFC_1_VALID_1_1_0),
	.valid_out(local_bb3_indvars_iv35_pop4__fu_valid_out),
	.stall_in(local_bb3_indvars_iv35_pop4__stall_local),
	.data_out(local_bb3_indvars_iv35_pop4_),
	.feedback_in(feedback_data_in_4),
	.feedback_valid_in(feedback_valid_in_4),
	.feedback_stall_out(feedback_stall_out_4)
);

defparam local_bb3_indvars_iv35_pop4__feedback.COALESCE_DISTANCE = 1;
defparam local_bb3_indvars_iv35_pop4__feedback.DATA_WIDTH = 64;
defparam local_bb3_indvars_iv35_pop4__feedback.STYLE = "REGULAR";

assign local_bb3_indvars_iv35_pop4__stall_local = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_c0_ene1_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_c0_ene1_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_c0_ene1_0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_c0_ene1_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_c0_ene1),
	.data_out(rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_c0_ene1_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb3_c0_ene1_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_c0_ene1_stall_in_1 = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_0_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_1_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_c0_ene1_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_2_NO_SHIFT_REG = rnode_1to2_bb3_c0_ene1_0_reg_2_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_1_VALID_1_2_0_inputs_ready;
 reg SFC_1_VALID_1_2_0_valid_out_0_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_0;
 reg SFC_1_VALID_1_2_0_valid_out_1_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_1;
 reg SFC_1_VALID_1_2_0_valid_out_2_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_2;
 reg SFC_1_VALID_1_2_0_valid_out_3_NO_SHIFT_REG;
wire SFC_1_VALID_1_2_0_stall_in_3;
wire SFC_1_VALID_1_2_0_output_regs_ready;
 reg SFC_1_VALID_1_2_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_1_2_0_causedstall;

assign SFC_1_VALID_1_2_0_inputs_ready = 1'b1;
assign SFC_1_VALID_1_2_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_1_1_0_stall_in_0 = 1'b0;
assign SFC_1_VALID_1_2_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_1_2_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_1_2_0_output_regs_ready)
		begin
			SFC_1_VALID_1_2_0_NO_SHIFT_REG <= SFC_1_VALID_1_1_0;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb3_indvars_iv35_pop4__0_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb3_indvars_iv35_pop4__1_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_2_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb3_indvars_iv35_pop4__2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb3_indvars_iv35_pop4__0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_0_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_0_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb3_indvars_iv35_pop4__0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb3_indvars_iv35_pop4_),
	.data_out(rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_fifo.DATA_WIDTH = 64;
defparam rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_indvars_iv35_pop4__stall_in = 1'b0;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_0_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_NO_SHIFT_REG = rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_indvars_iv35_pop4__1_NO_SHIFT_REG = rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_indvars_iv35_pop4__2_NO_SHIFT_REG = rnode_1to2_bb3_indvars_iv35_pop4__0_reg_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__acl_ffwd_dest_i1_9_stall_local;
wire local_bb3__acl_ffwd_dest_i1_9;

assign local_bb3__acl_ffwd_dest_i1_9 = ffwd_9_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_c0_ene1_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_c0_ene1_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_c0_ene1_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_c0_ene1_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_c0_ene1_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb3_c0_ene1_2_NO_SHIFT_REG),
	.data_out(rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_c0_ene1_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_c0_ene1_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_NO_SHIFT_REG = rnode_2to3_bb3_c0_ene1_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_1_VALID_2_3_0_inputs_ready;
 reg SFC_1_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_2_3_0_stall_in;
wire SFC_1_VALID_2_3_0_output_regs_ready;
 reg SFC_1_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_2_3_0_causedstall;

assign SFC_1_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_1_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_1_2_0_stall_in_0 = 1'b0;
assign SFC_1_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_2_3_0_output_regs_ready)
		begin
			SFC_1_VALID_2_3_0_NO_SHIFT_REG <= SFC_1_VALID_1_2_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_keep_going14_acl_pipeline_1_inputs_ready;
 reg local_bb3_keep_going14_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb3_keep_going14_acl_pipeline_1_stall_in;
wire local_bb3_keep_going14_acl_pipeline_1_output_regs_ready;
wire local_bb3_keep_going14_acl_pipeline_1_keep_going;
wire local_bb3_keep_going14_acl_pipeline_1_fu_valid_out;
wire local_bb3_keep_going14_acl_pipeline_1_fu_stall_out;
 reg local_bb3_keep_going14_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb3_keep_going14_acl_pipeline_1_feedback_pipelined;
wire local_bb3_keep_going14_acl_pipeline_1_causedstall;

acl_pipeline local_bb3_keep_going14_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb3_keep_going14_acl_pipeline_1_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_keep_going14_acl_pipeline_1_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_keep_going14_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_2),
	.not_exitcond_in(feedback_data_in_3),
	.not_exitcond_valid_in(feedback_valid_in_3),
	.not_exitcond_stall_out(feedback_stall_out_3),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb3_keep_going14_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb3_keep_going14_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb3_keep_going14_acl_pipeline_1_inputs_ready = 1'b1;
assign local_bb3_keep_going14_acl_pipeline_1_output_regs_ready = 1'b1;
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign SFC_1_VALID_1_2_0_stall_in_1 = 1'b0;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb3_keep_going14_acl_pipeline_1_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_keep_going14_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb3_keep_going14_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_keep_going14_acl_pipeline_1_output_regs_ready)
		begin
			local_bb3_keep_going14_acl_pipeline_1_NO_SHIFT_REG <= local_bb3_keep_going14_acl_pipeline_1_keep_going;
			local_bb3_keep_going14_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_keep_going14_acl_pipeline_1_stall_in))
			begin
				local_bb3_keep_going14_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_var__valid_out;
wire local_bb3_var__stall_in;
wire local_bb3_var__inputs_ready;
wire local_bb3_var__stall_local;
wire [31:0] local_bb3_var_;

assign local_bb3_var__inputs_ready = rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_var_ = rnode_1to2_bb3_indvars_iv35_pop4__0_NO_SHIFT_REG[31:0];
assign local_bb3_var__valid_out = 1'b1;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u12_valid_out;
wire local_bb3_var__u12_stall_in;
wire local_bb3_var__u12_inputs_ready;
wire local_bb3_var__u12_stall_local;
wire [63:0] local_bb3_var__u12;

assign local_bb3_var__u12_inputs_ready = rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_1_NO_SHIFT_REG;
assign local_bb3_var__u12 = (rnode_1to2_bb3_indvars_iv35_pop4__1_NO_SHIFT_REG + input_wii_var__u11);
assign local_bb3_var__u12_valid_out = 1'b1;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb3_indvars_iv_next36_stall_local;
wire [63:0] local_bb3_indvars_iv_next36;

assign local_bb3_indvars_iv_next36 = (rnode_1to2_bb3_indvars_iv35_pop4__2_NO_SHIFT_REG + 64'h1);

// This section implements an unregistered operation.
// 
wire local_bb3__acl_ffwd_dest_i32_4_stall_local;
wire [31:0] local_bb3__acl_ffwd_dest_i32_4;

assign local_bb3__acl_ffwd_dest_i32_4 = ffwd_4_0;

// This section implements a registered operation.
// 
wire SFC_1_VALID_3_4_0_inputs_ready;
 reg SFC_1_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_3_4_0_stall_in;
wire SFC_1_VALID_3_4_0_output_regs_ready;
 reg SFC_1_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_3_4_0_causedstall;

assign SFC_1_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_1_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_2_3_0_stall_in = 1'b0;
assign SFC_1_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_3_4_0_output_regs_ready)
		begin
			SFC_1_VALID_3_4_0_NO_SHIFT_REG <= SFC_1_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_keep_going14_acl_pipeline_1_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_keep_going14_acl_pipeline_1_stall_in = 1'b0;
assign rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_NO_SHIFT_REG = rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to3_bb3_var__0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to3_bb3_var__0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_var__0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_var__0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_var__0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_var__0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_var__0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_var_),
	.data_out(rnode_2to3_bb3_var__0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_var__0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_var__0_reg_3_fifo.DATA_WIDTH = 32;
defparam rnode_2to3_bb3_var__0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_var__0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_var__0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__stall_in = 1'b0;
assign rnode_2to3_bb3_var__0_NO_SHIFT_REG = rnode_2to3_bb3_var__0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_var__0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_var__0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_var__u12_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u12_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb3_var__u12_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u12_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_2to3_bb3_var__u12_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u12_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u12_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u12_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_var__u12_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_var__u12_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_var__u12_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_var__u12_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_var__u12_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_var__u12),
	.data_out(rnode_2to3_bb3_var__u12_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_var__u12_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_var__u12_0_reg_3_fifo.DATA_WIDTH = 64;
defparam rnode_2to3_bb3_var__u12_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_var__u12_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_var__u12_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u12_stall_in = 1'b0;
assign rnode_2to3_bb3_var__u12_0_NO_SHIFT_REG = rnode_2to3_bb3_var__u12_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_var__u12_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_var__u12_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u13_stall_local;
wire [31:0] local_bb3_var__u13;

assign local_bb3_var__u13 = local_bb3_indvars_iv_next36[31:0];

// This section implements a registered operation.
// 
wire SFC_1_VALID_4_5_0_inputs_ready;
 reg SFC_1_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_1_VALID_4_5_0_stall_in;
wire SFC_1_VALID_4_5_0_output_regs_ready;
 reg SFC_1_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_1_VALID_4_5_0_causedstall;

assign SFC_1_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_1_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_1_VALID_3_4_0_stall_in = 1'b0;
assign SFC_1_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_1_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_1_VALID_4_5_0_output_regs_ready)
		begin
			SFC_1_VALID_4_5_0_NO_SHIFT_REG <= SFC_1_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_add23_valid_out;
wire local_bb3_add23_stall_in;
wire local_bb3_add23_inputs_ready;
wire local_bb3_add23_stall_local;
wire [31:0] local_bb3_add23;

assign local_bb3_add23_inputs_ready = (rnode_2to3_bb3_c0_ene1_0_valid_out_NO_SHIFT_REG & rnode_2to3_bb3_var__0_valid_out_NO_SHIFT_REG);
assign local_bb3_add23 = (rnode_2to3_bb3_var__0_NO_SHIFT_REG + local_bb3__acl_ffwd_dest_i32_4);
assign local_bb3_add23_valid_out = 1'b1;
assign rnode_2to3_bb3_c0_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_var__0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb3_arrayidx41_inputs_ready;
 reg local_bb3_arrayidx41_valid_out_NO_SHIFT_REG;
wire local_bb3_arrayidx41_stall_in;
wire local_bb3_arrayidx41_output_regs_ready;
 reg [63:0] local_bb3_arrayidx41_NO_SHIFT_REG;
wire [63:0] local_bb3_arrayidx41_op_wire;
wire local_bb3_arrayidx41_causedstall;

assign local_bb3_arrayidx41_inputs_ready = 1'b1;
assign local_bb3_arrayidx41_output_regs_ready = 1'b1;
assign local_bb3_arrayidx41_op_wire = (64'h0 + (rnode_2to3_bb3_var__u12_0_NO_SHIFT_REG << 6'h2));
assign rnode_2to3_bb3_var__u12_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb3_arrayidx41_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_arrayidx41_NO_SHIFT_REG <= 'x;
		local_bb3_arrayidx41_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_arrayidx41_output_regs_ready)
		begin
			local_bb3_arrayidx41_NO_SHIFT_REG <= local_bb3_arrayidx41_op_wire;
			local_bb3_arrayidx41_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_arrayidx41_stall_in))
			begin
				local_bb3_arrayidx41_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_cmp15_stall_local;
wire local_bb3_cmp15;

assign local_bb3_cmp15 = ($signed(local_bb3_var__u13) > $signed(input_r));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_add23_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add23_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_add23_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add23_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add23_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_add23_1_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add23_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb3_add23_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add23_0_valid_out_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add23_0_stall_in_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_add23_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_add23_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_add23_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_add23_0_stall_in_0_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_add23_0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_add23_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_add23),
	.data_out(rnode_3to4_bb3_add23_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_add23_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_add23_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb3_add23_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_add23_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_add23_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_add23_stall_in = 1'b0;
assign rnode_3to4_bb3_add23_0_stall_in_0_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_add23_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_add23_0_NO_SHIFT_REG = rnode_3to4_bb3_add23_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_add23_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_add23_1_NO_SHIFT_REG = rnode_3to4_bb3_add23_0_reg_4_NO_SHIFT_REG;

// This section implements a registered operation.
// 
// Filescope constant lowered to ROM: gaussian.ROM41
wire local_bb3_gaussian_ROM41_arrayidx41_inputs_ready;
 reg local_bb3_gaussian_ROM41_arrayidx41_valid_out_NO_SHIFT_REG;
wire local_bb3_gaussian_ROM41_arrayidx41_stall_in;
wire local_bb3_gaussian_ROM41_arrayidx41_output_regs_ready;
 reg [31:0] local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG;
wire [63:0] local_bb3_gaussian_ROM41_arrayidx41$addr$ps;
wire local_bb3_gaussian_ROM41_arrayidx41_causedstall;

assign local_bb3_gaussian_ROM41_arrayidx41_inputs_ready = 1'b1;
assign local_bb3_gaussian_ROM41_arrayidx41_output_regs_ready = 1'b1;
assign local_bb3_gaussian_ROM41_arrayidx41$addr$ps = (local_bb3_arrayidx41_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign local_bb3_arrayidx41_stall_in = 1'b0;
assign local_bb3_gaussian_ROM41_arrayidx41_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (local_bb3_gaussian_ROM41_arrayidx41_output_regs_ready)
		begin
			case (local_bb3_gaussian_ROM41_arrayidx41$addr$ps[4:2])
				3'h0:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h3F61EB85;
				end

				3'h1:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h3F781D7E;
				end

				3'h2:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h3F800000;
				end

				3'h3:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h3F781D7E;
				end

				3'h4:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h3F61EB85;
				end

				3'h5:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h3F413A93;
				end

				3'h6:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h0;
				end

				3'h7:
				begin
					local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG <= 32'h0;
				end

				default:
				begin
				end

			endcase
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_gaussian_ROM41_arrayidx41_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_gaussian_ROM41_arrayidx41_output_regs_ready)
		begin
			local_bb3_gaussian_ROM41_arrayidx41_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_gaussian_ROM41_arrayidx41_stall_in))
			begin
				local_bb3_gaussian_ROM41_arrayidx41_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_var__u14_stall_local;
wire local_bb3_var__u14;

assign local_bb3_var__u14 = (local_bb3__acl_ffwd_dest_i1_9 | local_bb3_cmp15);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp1_i_valid_out;
wire local_bb3_cmp1_i_stall_in;
wire local_bb3_cmp1_i_inputs_ready;
wire local_bb3_cmp1_i_stall_local;
wire local_bb3_cmp1_i;

assign local_bb3_cmp1_i_inputs_ready = rnode_3to4_bb3_add23_0_valid_out_0_NO_SHIFT_REG;
assign local_bb3_cmp1_i = (rnode_3to4_bb3_add23_0_NO_SHIFT_REG > input_wii_sub24);
assign local_bb3_cmp1_i_valid_out = 1'b1;
assign rnode_3to4_bb3_add23_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_add23_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add23_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_add23_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add23_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_add23_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add23_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add23_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add23_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_add23_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_add23_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_add23_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_add23_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_add23_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_add23_1_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_add23_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_add23_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_add23_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3_add23_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_add23_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_add23_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_add23_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_add23_0_NO_SHIFT_REG = rnode_4to5_bb3_add23_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_add23_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_add23_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u14_valid_out_1;
wire local_bb3_var__u14_stall_in_1;
wire local_bb3_notexit16_valid_out_0;
wire local_bb3_notexit16_stall_in_0;
wire local_bb3_notexit16_valid_out_1;
wire local_bb3_notexit16_stall_in_1;
wire local_bb3_indvars_iv_next36_valid_out_1;
wire local_bb3_indvars_iv_next36_stall_in_1;
wire local_bb3_notexit16_inputs_ready;
wire local_bb3_notexit16_stall_local;
wire local_bb3_notexit16;

assign local_bb3_notexit16_inputs_ready = (rnode_1to2_bb3_c0_ene1_0_valid_out_1_NO_SHIFT_REG & rnode_1to2_bb3_indvars_iv35_pop4__0_valid_out_2_NO_SHIFT_REG);
assign local_bb3_notexit16 = (local_bb3_var__u14 ^ 1'b1);
assign local_bb3_var__u14_valid_out_1 = 1'b1;
assign local_bb3_notexit16_valid_out_0 = 1'b1;
assign local_bb3_notexit16_valid_out_1 = 1'b1;
assign local_bb3_indvars_iv_next36_valid_out_1 = 1'b1;
assign rnode_1to2_bb3_c0_ene1_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb3_indvars_iv35_pop4__0_stall_in_2_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_cmp1_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_cmp1_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_cmp1_i_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_cmp1_i_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_cmp1_i_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_cmp1_i_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_cmp1_i_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_cmp1_i_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_cmp1_i_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_cmp1_i_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_cmp1_i_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_cmp1_i_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_cmp1_i_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_cmp1_i),
	.data_out(rnode_4to5_bb3_cmp1_i_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_cmp1_i_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_cmp1_i_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_cmp1_i_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_cmp1_i_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_cmp1_i_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_cmp1_i_stall_in = 1'b0;
assign rnode_4to5_bb3_cmp1_i_0_NO_SHIFT_REG = rnode_4to5_bb3_cmp1_i_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_cmp1_i_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_cmp1_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb3_var__u14_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u14_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u14_0_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u14_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u14_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u14_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u14_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb3_var__u14_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb3_var__u14_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb3_var__u14_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb3_var__u14_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb3_var__u14_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb3_var__u14_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb3_var__u14),
	.data_out(rnode_2to3_bb3_var__u14_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb3_var__u14_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb3_var__u14_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb3_var__u14_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb3_var__u14_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb3_var__u14_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_var__u14_stall_in_1 = 1'b0;
assign rnode_2to3_bb3_var__u14_0_NO_SHIFT_REG = rnode_2to3_bb3_var__u14_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb3_var__u14_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb3_var__u14_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb3_notexitcond15_notexit16_inputs_ready;
 reg local_bb3_notexitcond15_notexit16_valid_out_NO_SHIFT_REG;
wire local_bb3_notexitcond15_notexit16_stall_in;
wire local_bb3_notexitcond15_notexit16_output_regs_ready;
wire local_bb3_notexitcond15_notexit16_result;
wire local_bb3_notexitcond15_notexit16_fu_valid_out;
wire local_bb3_notexitcond15_notexit16_fu_stall_out;
 reg local_bb3_notexitcond15_notexit16_NO_SHIFT_REG;
wire local_bb3_notexitcond15_notexit16_causedstall;

acl_push local_bb3_notexitcond15_notexit16_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(local_bb3_notexit16),
	.stall_out(local_bb3_notexitcond15_notexit16_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_notexitcond15_notexit16_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_notexitcond15_notexit16_result),
	.feedback_out(feedback_data_out_3),
	.feedback_valid_out(feedback_valid_out_3),
	.feedback_stall_in(feedback_stall_in_3)
);

defparam local_bb3_notexitcond15_notexit16_feedback.STALLFREE = 1;
defparam local_bb3_notexitcond15_notexit16_feedback.DATA_WIDTH = 1;
defparam local_bb3_notexitcond15_notexit16_feedback.FIFO_DEPTH = 1;
defparam local_bb3_notexitcond15_notexit16_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb3_notexitcond15_notexit16_feedback.STYLE = "REGULAR";

assign local_bb3_notexitcond15_notexit16_inputs_ready = 1'b1;
assign local_bb3_notexitcond15_notexit16_output_regs_ready = 1'b1;
assign local_bb3_notexit16_stall_in_0 = 1'b0;
assign SFC_1_VALID_1_2_0_stall_in_2 = 1'b0;
assign local_bb3_notexitcond15_notexit16_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_notexitcond15_notexit16_NO_SHIFT_REG <= 'x;
		local_bb3_notexitcond15_notexit16_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_notexitcond15_notexit16_output_regs_ready)
		begin
			local_bb3_notexitcond15_notexit16_NO_SHIFT_REG <= local_bb3_notexitcond15_notexit16_result;
			local_bb3_notexitcond15_notexit16_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_notexitcond15_notexit16_stall_in))
			begin
				local_bb3_notexitcond15_notexit16_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_indvars_iv35_push4_indvars_iv_next36_inputs_ready;
 reg local_bb3_indvars_iv35_push4_indvars_iv_next36_valid_out_NO_SHIFT_REG;
wire local_bb3_indvars_iv35_push4_indvars_iv_next36_stall_in;
wire local_bb3_indvars_iv35_push4_indvars_iv_next36_output_regs_ready;
wire [63:0] local_bb3_indvars_iv35_push4_indvars_iv_next36_result;
wire local_bb3_indvars_iv35_push4_indvars_iv_next36_fu_valid_out;
wire local_bb3_indvars_iv35_push4_indvars_iv_next36_fu_stall_out;
 reg [63:0] local_bb3_indvars_iv35_push4_indvars_iv_next36_NO_SHIFT_REG;
wire local_bb3_indvars_iv35_push4_indvars_iv_next36_causedstall;

acl_push local_bb3_indvars_iv35_push4_indvars_iv_next36_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb3_notexit16),
	.predicate(1'b0),
	.data_in(local_bb3_indvars_iv_next36),
	.stall_out(local_bb3_indvars_iv35_push4_indvars_iv_next36_fu_stall_out),
	.valid_in(SFC_1_VALID_1_2_0_NO_SHIFT_REG),
	.valid_out(local_bb3_indvars_iv35_push4_indvars_iv_next36_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb3_indvars_iv35_push4_indvars_iv_next36_result),
	.feedback_out(feedback_data_out_4),
	.feedback_valid_out(feedback_valid_out_4),
	.feedback_stall_in(feedback_stall_in_4)
);

defparam local_bb3_indvars_iv35_push4_indvars_iv_next36_feedback.STALLFREE = 1;
defparam local_bb3_indvars_iv35_push4_indvars_iv_next36_feedback.DATA_WIDTH = 64;
defparam local_bb3_indvars_iv35_push4_indvars_iv_next36_feedback.FIFO_DEPTH = 2;
defparam local_bb3_indvars_iv35_push4_indvars_iv_next36_feedback.MIN_FIFO_LATENCY = 1;
defparam local_bb3_indvars_iv35_push4_indvars_iv_next36_feedback.STYLE = "REGULAR";

assign local_bb3_indvars_iv35_push4_indvars_iv_next36_inputs_ready = 1'b1;
assign local_bb3_indvars_iv35_push4_indvars_iv_next36_output_regs_ready = 1'b1;
assign local_bb3_indvars_iv_next36_stall_in_1 = 1'b0;
assign local_bb3_notexit16_stall_in_1 = 1'b0;
assign SFC_1_VALID_1_2_0_stall_in_3 = 1'b0;
assign local_bb3_indvars_iv35_push4_indvars_iv_next36_causedstall = (SFC_1_VALID_1_2_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_indvars_iv35_push4_indvars_iv_next36_NO_SHIFT_REG <= 'x;
		local_bb3_indvars_iv35_push4_indvars_iv_next36_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_indvars_iv35_push4_indvars_iv_next36_output_regs_ready)
		begin
			local_bb3_indvars_iv35_push4_indvars_iv_next36_NO_SHIFT_REG <= local_bb3_indvars_iv35_push4_indvars_iv_next36_result;
			local_bb3_indvars_iv35_push4_indvars_iv_next36_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb3_indvars_iv35_push4_indvars_iv_next36_stall_in))
			begin
				local_bb3_indvars_iv35_push4_indvars_iv_next36_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_sub24_add23_stall_local;
wire [31:0] local_bb3_sub24_add23;

assign local_bb3_sub24_add23 = (rnode_4to5_bb3_cmp1_i_0_NO_SHIFT_REG ? input_wii_sub24 : rnode_4to5_bb3_add23_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb3_var__u14_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u14_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u14_0_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u14_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u14_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u14_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u14_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb3_var__u14_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb3_var__u14_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb3_var__u14_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb3_var__u14_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb3_var__u14_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb3_var__u14_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(rnode_2to3_bb3_var__u14_0_NO_SHIFT_REG),
	.data_out(rnode_3to4_bb3_var__u14_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb3_var__u14_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb3_var__u14_0_reg_4_fifo.DATA_WIDTH = 1;
defparam rnode_3to4_bb3_var__u14_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb3_var__u14_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb3_var__u14_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb3_var__u14_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_var__u14_0_NO_SHIFT_REG = rnode_3to4_bb3_var__u14_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb3_var__u14_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb3_var__u14_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_notexitcond15_notexit16_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb3_notexitcond15_notexit16_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb3_notexitcond15_notexit16_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb3_notexitcond15_notexit16_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_notexitcond15_notexit16_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_notexitcond15_notexit16_stall_in = 1'b0;
assign rnode_3to5_bb3_notexitcond15_notexit16_0_NO_SHIFT_REG = rnode_3to5_bb3_notexitcond15_notexit16_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb3_notexitcond15_notexit16_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_notexitcond15_notexit16_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_indvars_iv35_push4_indvars_iv_next36_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_fifo.DATA_WIDTH = 64;
defparam rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb3_indvars_iv35_push4_indvars_iv_next36_stall_in = 1'b0;
assign rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_NO_SHIFT_REG = rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi1_stall_local;
wire [127:0] local_bb3_c0_exi1;

assign local_bb3_c0_exi1[31:0] = 32'bx;
assign local_bb3_c0_exi1[63:32] = local_bb3_sub24_add23;
assign local_bb3_c0_exi1[127:64] = 64'bx;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_var__u14_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u14_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u14_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u14_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u14_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u14_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u14_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_var__u14_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_var__u14_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_var__u14_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_var__u14_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_var__u14_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_var__u14_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_3to4_bb3_var__u14_0_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb3_var__u14_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_var__u14_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb3_var__u14_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb3_var__u14_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb3_var__u14_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb3_var__u14_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to4_bb3_var__u14_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_var__u14_0_NO_SHIFT_REG = rnode_4to5_bb3_var__u14_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_var__u14_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_var__u14_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi2_stall_local;
wire [127:0] local_bb3_c0_exi2;

assign local_bb3_c0_exi2[63:0] = local_bb3_c0_exi1[63:0];
assign local_bb3_c0_exi2[95:64] = local_bb3_gaussian_ROM41_arrayidx41_NO_SHIFT_REG;
assign local_bb3_c0_exi2[127:96] = local_bb3_c0_exi1[127:96];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi3_stall_local;
wire [127:0] local_bb3_c0_exi3;

assign local_bb3_c0_exi3[95:0] = local_bb3_c0_exi2[95:0];
assign local_bb3_c0_exi3[96] = rnode_4to5_bb3_var__u14_0_NO_SHIFT_REG;
assign local_bb3_c0_exi3[127:97] = local_bb3_c0_exi2[127:97];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exi4_valid_out;
wire local_bb3_c0_exi4_stall_in;
wire local_bb3_c0_exi4_inputs_ready;
wire local_bb3_c0_exi4_stall_local;
wire [127:0] local_bb3_c0_exi4;

assign local_bb3_c0_exi4_inputs_ready = (rnode_3to5_bb3_notexitcond15_notexit16_0_valid_out_NO_SHIFT_REG & local_bb3_gaussian_ROM41_arrayidx41_valid_out_NO_SHIFT_REG & rnode_4to5_bb3_var__u14_0_valid_out_NO_SHIFT_REG & rnode_4to5_bb3_cmp1_i_0_valid_out_NO_SHIFT_REG & rnode_4to5_bb3_add23_0_valid_out_NO_SHIFT_REG);
assign local_bb3_c0_exi4[103:0] = local_bb3_c0_exi3[103:0];
assign local_bb3_c0_exi4[104] = rnode_3to5_bb3_notexitcond15_notexit16_0_NO_SHIFT_REG;
assign local_bb3_c0_exi4[127:105] = local_bb3_c0_exi3[127:105];
assign local_bb3_c0_exi4_valid_out = 1'b1;
assign rnode_3to5_bb3_notexitcond15_notexit16_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb3_gaussian_ROM41_arrayidx41_stall_in = 1'b0;
assign rnode_4to5_bb3_var__u14_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_cmp1_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb3_add23_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb3_c0_exit_c0_exi4_inputs_ready;
 reg local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_0;
 reg local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_1;
 reg local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_2;
 reg local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG;
wire local_bb3_c0_exit_c0_exi4_stall_in_3;
 reg [127:0] local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG;
wire [127:0] local_bb3_c0_exit_c0_exi4_in;
wire local_bb3_c0_exit_c0_exi4_valid;
wire local_bb3_c0_exit_c0_exi4_causedstall;

acl_stall_free_sink local_bb3_c0_exit_c0_exi4_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb3_c0_exi4),
	.data_out(local_bb3_c0_exit_c0_exi4_in),
	.input_accepted(local_bb3_c0_enter_c0_eni1_input_accepted),
	.valid_out(local_bb3_c0_exit_c0_exi4_valid),
	.stall_in(~(local_bb3_c0_exit_c0_exi4_output_regs_ready)),
	.stall_entry(local_bb3_c0_exit_c0_exi4_entry_stall),
	.valid_in(local_bb3_c0_exit_c0_exi4_valid_in),
	.IIphases(local_bb3_c0_exit_c0_exi4_phases),
	.inc_pipelined_thread(local_bb3_c0_enter_c0_eni1_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb3_c0_enter_c0_eni1_dec_pipelined_thread)
);

defparam local_bb3_c0_exit_c0_exi4_instance.DATA_WIDTH = 128;
defparam local_bb3_c0_exit_c0_exi4_instance.PIPELINE_DEPTH = 9;
defparam local_bb3_c0_exit_c0_exi4_instance.SHARINGII = 1;
defparam local_bb3_c0_exit_c0_exi4_instance.SCHEDULEII = 1;
defparam local_bb3_c0_exit_c0_exi4_instance.ALWAYS_THROTTLE = 0;

assign local_bb3_c0_exit_c0_exi4_inputs_ready = 1'b1;
assign local_bb3_c0_exit_c0_exi4_output_regs_ready = ((~(local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_0)) & (~(local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_1)) & (~(local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_2)) & (~(local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG) | ~(local_bb3_c0_exit_c0_exi4_stall_in_3)));
assign local_bb3_c0_exit_c0_exi4_valid_in = SFC_1_VALID_4_5_0_NO_SHIFT_REG;
assign local_bb3_c0_exi4_stall_in = 1'b0;
assign SFC_1_VALID_4_5_0_stall_in = 1'b0;
assign rnode_3to5_bb3_keep_going14_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb3_indvars_iv35_push4_indvars_iv_next36_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb3_c0_exit_c0_exi4_causedstall = (1'b1 && (1'b0 && !(~(local_bb3_c0_exit_c0_exi4_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG <= 'x;
		local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_c0_exit_c0_exi4_output_regs_ready)
		begin
			local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_in;
			local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
			local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
			local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
			local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG <= local_bb3_c0_exit_c0_exi4_valid;
		end
		else
		begin
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_0))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_1))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_2))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb3_c0_exit_c0_exi4_stall_in_3))
			begin
				local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe1_stall_local;
wire [31:0] local_bb3_c0_exe1;

assign local_bb3_c0_exe1 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe2_stall_local;
wire [31:0] local_bb3_c0_exe2;

assign local_bb3_c0_exe2 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[95:64];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe3_stall_local;
wire local_bb3_c0_exe3;

assign local_bb3_c0_exe3 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[96];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe4_valid_out;
wire local_bb3_c0_exe4_stall_in;
wire local_bb3_c0_exe3_valid_out;
wire local_bb3_c0_exe3_stall_in;
wire local_bb3_c0_exe2_valid_out;
wire local_bb3_c0_exe2_stall_in;
wire local_bb3_c0_exe1_valid_out;
wire local_bb3_c0_exe1_stall_in;
wire local_bb3_c0_exe4_inputs_ready;
wire local_bb3_c0_exe4_stall_local;
wire local_bb3_c0_exe4;

assign local_bb3_c0_exe4_inputs_ready = (local_bb3_c0_exit_c0_exi4_valid_out_3_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG & local_bb3_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG);
assign local_bb3_c0_exe4 = local_bb3_c0_exit_c0_exi4_NO_SHIFT_REG[104];
assign local_bb3_c0_exe4_stall_local = (local_bb3_c0_exe4_stall_in | local_bb3_c0_exe3_stall_in | local_bb3_c0_exe2_stall_in | local_bb3_c0_exe1_stall_in);
assign local_bb3_c0_exe4_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exe3_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exe2_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exe1_valid_out = local_bb3_c0_exe4_inputs_ready;
assign local_bb3_c0_exit_c0_exi4_stall_in_3 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));
assign local_bb3_c0_exit_c0_exi4_stall_in_2 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));
assign local_bb3_c0_exit_c0_exi4_stall_in_1 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));
assign local_bb3_c0_exit_c0_exi4_stall_in_0 = (local_bb3_c0_exe4_stall_local | ~(local_bb3_c0_exe4_inputs_ready));

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [31:0] lvb_bb3_c0_exe1_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_c0_exe2_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe3_reg_NO_SHIFT_REG;
 reg lvb_bb3_c0_exe4_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_t_228_pop5__reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb3_sum_227_pop6__reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb3_sum_227_pop6__valid_out_NO_SHIFT_REG & local_bb3_t_228_pop5__valid_out_NO_SHIFT_REG & local_bb3_c0_exe4_valid_out & local_bb3_c0_exe3_valid_out & local_bb3_c0_exe2_valid_out & local_bb3_c0_exe1_valid_out);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb3_sum_227_pop6__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_t_228_pop5__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe4_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe3_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb3_c0_exe1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb3_c0_exe1 = lvb_bb3_c0_exe1_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe2 = lvb_bb3_c0_exe2_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe3 = lvb_bb3_c0_exe3_reg_NO_SHIFT_REG;
assign lvb_bb3_c0_exe4 = lvb_bb3_c0_exe4_reg_NO_SHIFT_REG;
assign lvb_bb3_t_228_pop5_ = lvb_bb3_t_228_pop5__reg_NO_SHIFT_REG;
assign lvb_bb3_sum_227_pop6_ = lvb_bb3_sum_227_pop6__reg_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb3_c0_exe1_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe2_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe3_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_c0_exe4_reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_t_228_pop5__reg_NO_SHIFT_REG <= 'x;
		lvb_bb3_sum_227_pop6__reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb3_c0_exe1_reg_NO_SHIFT_REG <= local_bb3_c0_exe1;
			lvb_bb3_c0_exe2_reg_NO_SHIFT_REG <= local_bb3_c0_exe2;
			lvb_bb3_c0_exe3_reg_NO_SHIFT_REG <= local_bb3_c0_exe3;
			lvb_bb3_c0_exe4_reg_NO_SHIFT_REG <= local_bb3_c0_exe4;
			lvb_bb3_t_228_pop5__reg_NO_SHIFT_REG <= local_bb3_t_228_pop5__NO_SHIFT_REG;
			lvb_bb3_sum_227_pop6__reg_NO_SHIFT_REG <= local_bb3_sum_227_pop6__NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_4
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_global_size_0,
		input [63:0] 		input_in,
		input [31:0] 		input_r,
		input 		input_wii_cmp1526,
		input [31:0] 		input_wii_sub24,
		input [31:0] 		input_wii_sub27,
		input [31:0] 		input_wii_mul48,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u15,
		input 		valid_in_0,
		output 		stall_out_0,
		input [31:0] 		input_t_322_0,
		input [31:0] 		input_sum_321_0,
		input 		input_forked17_0,
		input [31:0] 		input_sub24_add2318_0,
		input [31:0] 		input_gaussian_ROM4119_0,
		input 		input_var__u16_0,
		input 		input_notexitcond1520_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [31:0] 		input_t_322_1,
		input [31:0] 		input_sum_321_1,
		input 		input_forked17_1,
		input [31:0] 		input_sub24_add2318_1,
		input [31:0] 		input_gaussian_ROM4119_1,
		input 		input_var__u16_1,
		input 		input_notexitcond1520_1,
		output 		valid_out_0,
		input 		stall_in_0,
		output [191:0] 		lvb_bb4_c0_exit28_c0_exi6_0,
		output 		lvb_bb4_c0_exe6_0,
		output [95:0] 		lvb_bb4_c1_exit_c1_exi2_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [191:0] 		lvb_bb4_c0_exit28_c0_exi6_1,
		output 		lvb_bb4_c0_exe6_1,
		output [95:0] 		lvb_bb4_c1_exit_c1_exi2_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		ffwd_9_0,
		input [31:0] 		ffwd_0_0,
		input 		feedback_valid_in_7,
		output 		feedback_stall_out_7,
		input [63:0] 		feedback_data_in_7,
		input 		feedback_valid_in_11,
		output 		feedback_stall_out_11,
		input [31:0] 		feedback_data_in_11,
		output 		feedback_stall_out_0,
		input 		feedback_valid_in_1,
		output 		feedback_stall_out_1,
		input 		feedback_data_in_1,
		output 		acl_pipelined_valid,
		input 		acl_pipelined_stall,
		output 		acl_pipelined_exiting_valid,
		output 		acl_pipelined_exiting_stall,
		input 		feedback_valid_in_10,
		output 		feedback_stall_out_10,
		input [31:0] 		feedback_data_in_10,
		input 		feedback_valid_in_12,
		output 		feedback_stall_out_12,
		input 		feedback_data_in_12,
		input 		feedback_valid_in_13,
		output 		feedback_stall_out_13,
		input 		feedback_data_in_13,
		output 		feedback_valid_out_7,
		input 		feedback_stall_in_7,
		output [63:0] 		feedback_data_out_7,
		output 		feedback_valid_out_1,
		input 		feedback_stall_in_1,
		output 		feedback_data_out_1,
		output 		feedback_valid_out_10,
		input 		feedback_stall_in_10,
		output [31:0] 		feedback_data_out_10,
		output 		feedback_valid_out_12,
		input 		feedback_stall_in_12,
		output 		feedback_data_out_12,
		output 		feedback_valid_out_13,
		input 		feedback_stall_in_13,
		output 		feedback_data_out_13,
		output 		feedback_valid_out_11,
		input 		feedback_stall_in_11,
		output [31:0] 		feedback_data_out_11,
		input [511:0] 		avm_local_bb4_ld__readdata,
		input 		avm_local_bb4_ld__readdatavalid,
		input 		avm_local_bb4_ld__waitrequest,
		output [32:0] 		avm_local_bb4_ld__address,
		output 		avm_local_bb4_ld__read,
		output 		avm_local_bb4_ld__write,
		input 		avm_local_bb4_ld__writeack,
		output [511:0] 		avm_local_bb4_ld__writedata,
		output [63:0] 		avm_local_bb4_ld__byteenable,
		output [4:0] 		avm_local_bb4_ld__burstcount,
		output 		local_bb4_ld__active,
		input 		clock2x,
		input [31:0] 		ffwd_7_0,
		input 		feedback_valid_in_9,
		output 		feedback_stall_out_9,
		input [31:0] 		feedback_data_in_9,
		input 		feedback_valid_in_8,
		output 		feedback_stall_out_8,
		input [31:0] 		feedback_data_in_8,
		output 		feedback_valid_out_9,
		input 		feedback_stall_in_9,
		output [31:0] 		feedback_data_out_9,
		output [31:0] 		ffwd_10_0,
		output 		feedback_valid_out_8,
		input 		feedback_stall_in_8,
		output [31:0] 		feedback_data_out_8,
		output [31:0] 		ffwd_11_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_322_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_321_0_staging_reg_NO_SHIFT_REG;
 reg input_forked17_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sub24_add2318_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_gaussian_ROM4119_0_staging_reg_NO_SHIFT_REG;
 reg input_var__u16_0_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1520_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_t_322_NO_SHIFT_REG;
 reg [31:0] local_lvm_sum_321_NO_SHIFT_REG;
 reg local_lvm_forked17_NO_SHIFT_REG;
 reg [31:0] local_lvm_sub24_add2318_NO_SHIFT_REG;
 reg [31:0] local_lvm_gaussian_ROM4119_NO_SHIFT_REG;
 reg local_lvm_var__u16_NO_SHIFT_REG;
 reg local_lvm_notexitcond1520_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_t_322_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sum_321_1_staging_reg_NO_SHIFT_REG;
 reg input_forked17_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_sub24_add2318_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_gaussian_ROM4119_1_staging_reg_NO_SHIFT_REG;
 reg input_var__u16_1_staging_reg_NO_SHIFT_REG;
 reg input_notexitcond1520_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_t_322_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_321_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_forked17_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_sub24_add2318_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_gaussian_ROM4119_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u16_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1520_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_t_322_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_sum_321_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_forked17_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_sub24_add2318_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_gaussian_ROM4119_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_var__u16_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_notexitcond1520_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_t_322_0_staging_reg_NO_SHIFT_REG <= input_t_322_0;
				input_sum_321_0_staging_reg_NO_SHIFT_REG <= input_sum_321_0;
				input_forked17_0_staging_reg_NO_SHIFT_REG <= input_forked17_0;
				input_sub24_add2318_0_staging_reg_NO_SHIFT_REG <= input_sub24_add2318_0;
				input_gaussian_ROM4119_0_staging_reg_NO_SHIFT_REG <= input_gaussian_ROM4119_0;
				input_var__u16_0_staging_reg_NO_SHIFT_REG <= input_var__u16_0;
				input_notexitcond1520_0_staging_reg_NO_SHIFT_REG <= input_notexitcond1520_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_t_322_1_staging_reg_NO_SHIFT_REG <= input_t_322_1;
				input_sum_321_1_staging_reg_NO_SHIFT_REG <= input_sum_321_1;
				input_forked17_1_staging_reg_NO_SHIFT_REG <= input_forked17_1;
				input_sub24_add2318_1_staging_reg_NO_SHIFT_REG <= input_sub24_add2318_1;
				input_gaussian_ROM4119_1_staging_reg_NO_SHIFT_REG <= input_gaussian_ROM4119_1;
				input_var__u16_1_staging_reg_NO_SHIFT_REG <= input_var__u16_1;
				input_notexitcond1520_1_staging_reg_NO_SHIFT_REG <= input_notexitcond1520_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_t_322_NO_SHIFT_REG <= input_t_322_0_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_321_NO_SHIFT_REG <= input_sum_321_0_staging_reg_NO_SHIFT_REG;
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_0_staging_reg_NO_SHIFT_REG;
					local_lvm_sub24_add2318_NO_SHIFT_REG <= input_sub24_add2318_0_staging_reg_NO_SHIFT_REG;
					local_lvm_gaussian_ROM4119_NO_SHIFT_REG <= input_gaussian_ROM4119_0_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_0_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1520_NO_SHIFT_REG <= input_notexitcond1520_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_t_322_NO_SHIFT_REG <= input_t_322_0;
					local_lvm_sum_321_NO_SHIFT_REG <= input_sum_321_0;
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_0;
					local_lvm_sub24_add2318_NO_SHIFT_REG <= input_sub24_add2318_0;
					local_lvm_gaussian_ROM4119_NO_SHIFT_REG <= input_gaussian_ROM4119_0;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_0;
					local_lvm_notexitcond1520_NO_SHIFT_REG <= input_notexitcond1520_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_t_322_NO_SHIFT_REG <= input_t_322_1_staging_reg_NO_SHIFT_REG;
					local_lvm_sum_321_NO_SHIFT_REG <= input_sum_321_1_staging_reg_NO_SHIFT_REG;
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_1_staging_reg_NO_SHIFT_REG;
					local_lvm_sub24_add2318_NO_SHIFT_REG <= input_sub24_add2318_1_staging_reg_NO_SHIFT_REG;
					local_lvm_gaussian_ROM4119_NO_SHIFT_REG <= input_gaussian_ROM4119_1_staging_reg_NO_SHIFT_REG;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_1_staging_reg_NO_SHIFT_REG;
					local_lvm_notexitcond1520_NO_SHIFT_REG <= input_notexitcond1520_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_t_322_NO_SHIFT_REG <= input_t_322_1;
					local_lvm_sum_321_NO_SHIFT_REG <= input_sum_321_1;
					local_lvm_forked17_NO_SHIFT_REG <= input_forked17_1;
					local_lvm_sub24_add2318_NO_SHIFT_REG <= input_sub24_add2318_1;
					local_lvm_gaussian_ROM4119_NO_SHIFT_REG <= input_gaussian_ROM4119_1;
					local_lvm_var__u16_NO_SHIFT_REG <= input_var__u16_1;
					local_lvm_notexitcond1520_NO_SHIFT_REG <= input_notexitcond1520_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni121_stall_local;
wire [127:0] local_bb4_c0_eni121;

assign local_bb4_c0_eni121[7:0] = 8'bx;
assign local_bb4_c0_eni121[8] = local_lvm_forked17_NO_SHIFT_REG;
assign local_bb4_c0_eni121[127:9] = 119'bx;

// Register node:
//  * latency = 14
//  * capacity = 14
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_out_reg_15_NO_SHIFT_REG;
wire [64:0] rci_rcnode_1to175_rc6_t_322_0_reg_1;

acl_data_fifo rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_fifo.DEPTH = 15;
defparam rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_fifo.IMPL = "ram";

assign rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_reg_15_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign merge_node_stall_in_5 = rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_out_reg_15_NO_SHIFT_REG;
assign rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_in_reg_15_NO_SHIFT_REG = rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG;
assign rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG = rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_valid_out_reg_15_NO_SHIFT_REG;
assign rci_rcnode_1to175_rc6_t_322_0_reg_1[31:0] = local_lvm_t_322_NO_SHIFT_REG;
assign rci_rcnode_1to175_rc6_t_322_0_reg_1[32] = local_lvm_forked17_NO_SHIFT_REG;
assign rci_rcnode_1to175_rc6_t_322_0_reg_1[64:33] = local_lvm_sum_321_NO_SHIFT_REG;

// Register node:
//  * latency = 174
//  * capacity = 174
 logic rcnode_1to175_rc6_t_322_0_valid_out_NO_SHIFT_REG;
 logic rcnode_1to175_rc6_t_322_0_stall_in_NO_SHIFT_REG;
 logic [64:0] rcnode_1to175_rc6_t_322_0_NO_SHIFT_REG;
 logic rcnode_1to175_rc6_t_322_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [64:0] rcnode_1to175_rc6_t_322_0_reg_175_NO_SHIFT_REG;
 logic rcnode_1to175_rc6_t_322_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rcnode_1to175_rc6_t_322_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rcnode_1to175_rc6_t_322_0_stall_out_reg_175_IP_NO_SHIFT_REG;
 logic rcnode_1to175_rc6_t_322_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rcnode_1to175_rc6_t_322_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_1to175_rc6_t_322_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_1to175_rc6_t_322_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rcnode_1to175_rc6_t_322_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rcnode_1to175_rc6_t_322_0_stall_out_reg_175_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_1to175_rc6_t_322_0_reg_1),
	.data_out(rcnode_1to175_rc6_t_322_0_reg_175_NO_SHIFT_REG)
);

defparam rcnode_1to175_rc6_t_322_0_reg_175_fifo.DEPTH = 175;
defparam rcnode_1to175_rc6_t_322_0_reg_175_fifo.DATA_WIDTH = 65;
defparam rcnode_1to175_rc6_t_322_0_reg_175_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_1to175_rc6_t_322_0_reg_175_fifo.IMPL = "ram";

assign rcnode_1to175_rc6_t_322_0_reg_175_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_6_NO_SHIFT_REG;
assign rcnode_1to175_rc6_t_322_0_stall_out_reg_175_NO_SHIFT_REG = (~(rcnode_1to175_rc6_t_322_0_reg_175_inputs_ready_NO_SHIFT_REG) | rcnode_1to175_rc6_t_322_0_stall_out_reg_175_IP_NO_SHIFT_REG);
assign merge_node_stall_in_6 = rcnode_1to175_rc6_t_322_0_stall_out_reg_175_NO_SHIFT_REG;
assign rcnode_1to175_rc6_t_322_0_NO_SHIFT_REG = rcnode_1to175_rc6_t_322_0_reg_175_NO_SHIFT_REG;
assign rcnode_1to175_rc6_t_322_0_stall_in_reg_175_NO_SHIFT_REG = rcnode_1to175_rc6_t_322_0_stall_in_NO_SHIFT_REG;
assign rcnode_1to175_rc6_t_322_0_valid_out_NO_SHIFT_REG = rcnode_1to175_rc6_t_322_0_valid_out_reg_175_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni2_stall_local;
wire [127:0] local_bb4_c0_eni2;

assign local_bb4_c0_eni2[31:0] = local_bb4_c0_eni121[31:0];
assign local_bb4_c0_eni2[63:32] = local_lvm_sub24_add2318_NO_SHIFT_REG;
assign local_bb4_c0_eni2[127:64] = local_bb4_c0_eni121[127:64];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_out_reg_16_NO_SHIFT_REG;
wire [64:0] rci_rcnode_175to176_rc0_t_322_0_reg_175;

acl_data_fifo rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_fifo.DEPTH = 2;
defparam rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_fifo.IMPL = "ll_reg";

assign rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_reg_16_inputs_ready_NO_SHIFT_REG = rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG;
assign rnode_1to15_bb4__acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG = rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_out_reg_16_NO_SHIFT_REG;
assign rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_in_reg_16_NO_SHIFT_REG = rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG;
assign rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG = rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_valid_out_reg_16_NO_SHIFT_REG;
assign rci_rcnode_175to176_rc0_t_322_0_reg_175[31:0] = rcnode_1to175_rc6_t_322_0_NO_SHIFT_REG[31:0];
assign rci_rcnode_175to176_rc0_t_322_0_reg_175[32] = rcnode_1to175_rc6_t_322_0_NO_SHIFT_REG[32];
assign rci_rcnode_175to176_rc0_t_322_0_reg_175[64:33] = rcnode_1to175_rc6_t_322_0_NO_SHIFT_REG[64:33];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_175to176_rc0_t_322_0_valid_out_0_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_stall_in_0_NO_SHIFT_REG;
 logic [64:0] rcnode_175to176_rc0_t_322_0_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_valid_out_1_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_stall_in_1_NO_SHIFT_REG;
 logic [64:0] rcnode_175to176_rc0_t_322_1_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_valid_out_2_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_stall_in_2_NO_SHIFT_REG;
 logic [64:0] rcnode_175to176_rc0_t_322_2_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_valid_out_3_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_stall_in_3_NO_SHIFT_REG;
 logic [64:0] rcnode_175to176_rc0_t_322_3_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [64:0] rcnode_175to176_rc0_t_322_0_reg_176_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_stall_out_reg_176_IP_NO_SHIFT_REG;
 logic rcnode_175to176_rc0_t_322_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rcnode_175to176_rc0_t_322_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_175to176_rc0_t_322_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_175to176_rc0_t_322_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rcnode_175to176_rc0_t_322_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rcnode_175to176_rc0_t_322_0_stall_out_reg_176_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_175to176_rc0_t_322_0_reg_175),
	.data_out(rcnode_175to176_rc0_t_322_0_reg_176_NO_SHIFT_REG)
);

defparam rcnode_175to176_rc0_t_322_0_reg_176_fifo.DEPTH = 1;
defparam rcnode_175to176_rc0_t_322_0_reg_176_fifo.DATA_WIDTH = 65;
defparam rcnode_175to176_rc0_t_322_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_175to176_rc0_t_322_0_reg_176_fifo.IMPL = "ll_reg";

assign rcnode_175to176_rc0_t_322_0_reg_176_inputs_ready_NO_SHIFT_REG = rcnode_1to175_rc6_t_322_0_valid_out_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_0_stall_out_reg_176_NO_SHIFT_REG = (~(rcnode_175to176_rc0_t_322_0_reg_176_inputs_ready_NO_SHIFT_REG) | rcnode_175to176_rc0_t_322_0_stall_out_reg_176_IP_NO_SHIFT_REG);
assign rcnode_1to175_rc6_t_322_0_stall_in_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_stall_out_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_0_stall_in_0_reg_176_NO_SHIFT_REG = (rcnode_175to176_rc0_t_322_0_stall_in_0_NO_SHIFT_REG | rcnode_175to176_rc0_t_322_0_stall_in_1_NO_SHIFT_REG | rcnode_175to176_rc0_t_322_0_stall_in_2_NO_SHIFT_REG | rcnode_175to176_rc0_t_322_0_stall_in_3_NO_SHIFT_REG);
assign rcnode_175to176_rc0_t_322_0_valid_out_0_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_0_valid_out_1_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_0_valid_out_2_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_0_valid_out_3_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_0_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_1_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_2_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_reg_176_NO_SHIFT_REG;
assign rcnode_175to176_rc0_t_322_3_NO_SHIFT_REG = rcnode_175to176_rc0_t_322_0_reg_176_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni3_stall_local;
wire [127:0] local_bb4_c0_eni3;

assign local_bb4_c0_eni3[63:0] = local_bb4_c0_eni2[63:0];
assign local_bb4_c0_eni3[95:64] = local_lvm_gaussian_ROM4119_NO_SHIFT_REG;
assign local_bb4_c0_eni3[127:96] = local_bb4_c0_eni2[127:96];

// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_i1_9_valid_out;
wire local_bb4__acl_ffwd_dest_i1_9_stall_in;
wire local_bb4__acl_ffwd_dest_i1_9_inputs_ready;
wire local_bb4__acl_ffwd_dest_i1_9_stall_local;
wire local_bb4__acl_ffwd_dest_i1_9;

assign local_bb4__acl_ffwd_dest_i1_9_inputs_ready = rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_valid_out_NO_SHIFT_REG;
assign local_bb4__acl_ffwd_dest_i1_9 = ffwd_9_0;
assign local_bb4__acl_ffwd_dest_i1_9_valid_out = local_bb4__acl_ffwd_dest_i1_9_inputs_ready;
assign local_bb4__acl_ffwd_dest_i1_9_stall_local = local_bb4__acl_ffwd_dest_i1_9_stall_in;
assign rnode_15to16_bb4__acl_ffwd_dest_i1_9_0_stall_in_NO_SHIFT_REG = (|local_bb4__acl_ffwd_dest_i1_9_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni4_stall_local;
wire [127:0] local_bb4_c0_eni4;

assign local_bb4_c0_eni4[95:0] = local_bb4_c0_eni3[95:0];
assign local_bb4_c0_eni4[96] = local_lvm_var__u16_NO_SHIFT_REG;
assign local_bb4_c0_eni4[127:97] = local_bb4_c0_eni3[127:97];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_eni5_stall_local;
wire [127:0] local_bb4_c0_eni5;

assign local_bb4_c0_eni5[103:0] = local_bb4_c0_eni4[103:0];
assign local_bb4_c0_eni5[104] = local_lvm_notexitcond1520_NO_SHIFT_REG;
assign local_bb4_c0_eni5[127:105] = local_bb4_c0_eni4[127:105];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene123_valid_out;
wire local_bb4_c0_ene123_stall_in;
wire local_bb4_c0_ene2_valid_out;
wire local_bb4_c0_ene2_stall_in;
wire local_bb4_c0_ene3_valid_out;
wire local_bb4_c0_ene3_stall_in;
wire local_bb4_c0_ene4_valid_out;
wire local_bb4_c0_ene4_stall_in;
wire local_bb4_c0_ene5_valid_out;
wire local_bb4_c0_ene5_stall_in;
wire SFC_2_VALID_1_1_0_valid_out;
wire SFC_2_VALID_1_1_0_stall_in;
wire local_bb4_c0_enter22_c0_eni5_inputs_ready;
wire local_bb4_c0_enter22_c0_eni5_stall_local;
wire local_bb4_c0_enter22_c0_eni5_input_accepted;
wire [127:0] local_bb4_c0_enter22_c0_eni5;
wire local_bb4_c0_exit28_c0_exi6_entry_stall;
wire local_bb4_c0_enter22_c0_eni5_valid_bit;
wire local_bb4_c0_exit28_c0_exi6_output_regs_ready;
wire local_bb4_c0_exit28_c0_exi6_valid_in;
wire local_bb4_c0_exit28_c0_exi6_phases;
wire local_bb4_c0_enter22_c0_eni5_inc_pipelined_thread;
wire local_bb4_c0_enter22_c0_eni5_dec_pipelined_thread;
wire local_bb4_c0_enter22_c0_eni5_fu_stall_out;

assign local_bb4_c0_enter22_c0_eni5_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_3_NO_SHIFT_REG & merge_node_valid_out_4_NO_SHIFT_REG);
assign local_bb4_c0_enter22_c0_eni5 = local_bb4_c0_eni5;
assign local_bb4_c0_enter22_c0_eni5_input_accepted = (local_bb4_c0_enter22_c0_eni5_inputs_ready && !(local_bb4_c0_exit28_c0_exi6_entry_stall));
assign local_bb4_c0_enter22_c0_eni5_valid_bit = local_bb4_c0_enter22_c0_eni5_input_accepted;
assign local_bb4_c0_enter22_c0_eni5_inc_pipelined_thread = 1'b1;
assign local_bb4_c0_enter22_c0_eni5_dec_pipelined_thread = ~(1'b0);
assign local_bb4_c0_enter22_c0_eni5_fu_stall_out = (~(local_bb4_c0_enter22_c0_eni5_inputs_ready) | local_bb4_c0_exit28_c0_exi6_entry_stall);
assign local_bb4_c0_enter22_c0_eni5_stall_local = (local_bb4_c0_ene123_stall_in | local_bb4_c0_ene2_stall_in | local_bb4_c0_ene3_stall_in | local_bb4_c0_ene4_stall_in | local_bb4_c0_ene5_stall_in | SFC_2_VALID_1_1_0_stall_in);
assign local_bb4_c0_ene123_valid_out = local_bb4_c0_enter22_c0_eni5_inputs_ready;
assign local_bb4_c0_ene2_valid_out = local_bb4_c0_enter22_c0_eni5_inputs_ready;
assign local_bb4_c0_ene3_valid_out = local_bb4_c0_enter22_c0_eni5_inputs_ready;
assign local_bb4_c0_ene4_valid_out = local_bb4_c0_enter22_c0_eni5_inputs_ready;
assign local_bb4_c0_ene5_valid_out = local_bb4_c0_enter22_c0_eni5_inputs_ready;
assign SFC_2_VALID_1_1_0_valid_out = local_bb4_c0_enter22_c0_eni5_inputs_ready;
assign merge_node_stall_in_0 = (local_bb4_c0_enter22_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter22_c0_eni5_inputs_ready));
assign merge_node_stall_in_1 = (local_bb4_c0_enter22_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter22_c0_eni5_inputs_ready));
assign merge_node_stall_in_2 = (local_bb4_c0_enter22_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter22_c0_eni5_inputs_ready));
assign merge_node_stall_in_3 = (local_bb4_c0_enter22_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter22_c0_eni5_inputs_ready));
assign merge_node_stall_in_4 = (local_bb4_c0_enter22_c0_eni5_fu_stall_out | ~(local_bb4_c0_enter22_c0_eni5_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene123_stall_local;
wire local_bb4_c0_ene123;

assign local_bb4_c0_ene123 = local_bb4_c0_enter22_c0_eni5[8];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene2_stall_local;
wire [31:0] local_bb4_c0_ene2;

assign local_bb4_c0_ene2 = local_bb4_c0_enter22_c0_eni5[63:32];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene3_stall_local;
wire [31:0] local_bb4_c0_ene3;

assign local_bb4_c0_ene3 = local_bb4_c0_enter22_c0_eni5[95:64];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene4_stall_local;
wire local_bb4_c0_ene4;

assign local_bb4_c0_ene4 = local_bb4_c0_enter22_c0_eni5[96];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_ene5_stall_local;
wire local_bb4_c0_ene5;

assign local_bb4_c0_ene5 = local_bb4_c0_enter22_c0_eni5[104];

// This section implements an unregistered operation.
// 
wire SFC_2_VALID_1_1_0_stall_local;
wire SFC_2_VALID_1_1_0;

assign SFC_2_VALID_1_1_0 = local_bb4_c0_enter22_c0_eni5_valid_bit;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_1to3_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_1_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_2_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_valid_out_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_stall_in_0_reg_3_NO_SHIFT_REG;
 logic rnode_1to3_bb4_c0_ene123_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_1to3_bb4_c0_ene123_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to3_bb4_c0_ene123_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to3_bb4_c0_ene123_0_stall_in_0_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_1to3_bb4_c0_ene123_0_valid_out_0_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_1to3_bb4_c0_ene123_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene123),
	.data_out(rnode_1to3_bb4_c0_ene123_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_1to3_bb4_c0_ene123_0_reg_3_fifo.DEPTH = 2;
defparam rnode_1to3_bb4_c0_ene123_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_1to3_bb4_c0_ene123_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to3_bb4_c0_ene123_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_1to3_bb4_c0_ene123_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene123_stall_in = 1'b0;
assign rnode_1to3_bb4_c0_ene123_0_stall_in_0_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_1to3_bb4_c0_ene123_0_NO_SHIFT_REG = rnode_1to3_bb4_c0_ene123_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_1to3_bb4_c0_ene123_1_NO_SHIFT_REG = rnode_1to3_bb4_c0_ene123_0_reg_3_NO_SHIFT_REG;
assign rnode_1to3_bb4_c0_ene123_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_1to3_bb4_c0_ene123_2_NO_SHIFT_REG = rnode_1to3_bb4_c0_ene123_0_reg_3_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene2_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene2_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene2_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene2_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene2_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene2_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene2_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene2),
	.data_out(rnode_1to2_bb4_c0_ene2_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene2_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene2_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene2_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene2_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene2_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene2_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to2_bb4_c0_ene3_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene3_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene3_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene3_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene3_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene3_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene3_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene3),
	.data_out(rnode_1to2_bb4_c0_ene3_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.DATA_WIDTH = 32;
defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene3_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene3_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene3_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene3_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene3_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene3_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene4_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene4_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene4_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene4_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene4_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene4_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene4),
	.data_out(rnode_1to2_bb4_c0_ene4_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene4_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene4_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene4_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene4_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene4_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene4_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb4_c0_ene5_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb4_c0_ene5_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb4_c0_ene5_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb4_c0_ene5_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb4_c0_ene5_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb4_c0_ene5_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb4_c0_ene5),
	.data_out(rnode_1to2_bb4_c0_ene5_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb4_c0_ene5_0_reg_2_fifo.IMPL = "shift_reg";

assign rnode_1to2_bb4_c0_ene5_0_reg_2_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c0_ene5_stall_in = 1'b0;
assign rnode_1to2_bb4_c0_ene5_0_NO_SHIFT_REG = rnode_1to2_bb4_c0_ene5_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb4_c0_ene5_0_stall_in_reg_2_NO_SHIFT_REG = 1'b0;
assign rnode_1to2_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_1_2_0_inputs_ready;
 reg SFC_2_VALID_1_2_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_1_2_0_stall_in;
wire SFC_2_VALID_1_2_0_output_regs_ready;
 reg SFC_2_VALID_1_2_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_1_2_0_causedstall;

assign SFC_2_VALID_1_2_0_inputs_ready = 1'b1;
assign SFC_2_VALID_1_2_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_1_1_0_stall_in = 1'b0;
assign SFC_2_VALID_1_2_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_1_2_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_1_2_0_output_regs_ready)
		begin
			SFC_2_VALID_1_2_0_NO_SHIFT_REG <= SFC_2_VALID_1_1_0;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_pos_y_02_acl_ffwd_dest_i32_0_stall_local;
wire [31:0] local_bb4_pos_y_02_acl_ffwd_dest_i32_0;

assign local_bb4_pos_y_02_acl_ffwd_dest_i32_0 = ffwd_0_0;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_1_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_valid_out_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_stall_in_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_c0_ene123_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb4_c0_ene123_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb4_c0_ene123_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb4_c0_ene123_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb4_c0_ene123_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb4_c0_ene123_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_1to3_bb4_c0_ene123_2_NO_SHIFT_REG),
	.data_out(rnode_3to5_bb4_c0_ene123_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb4_c0_ene123_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb4_c0_ene123_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_3to5_bb4_c0_ene123_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb4_c0_ene123_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb4_c0_ene123_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to3_bb4_c0_ene123_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb4_c0_ene123_0_stall_in_0_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_3to5_bb4_c0_ene123_0_NO_SHIFT_REG = rnode_3to5_bb4_c0_ene123_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_3to5_bb4_c0_ene123_1_NO_SHIFT_REG = rnode_3to5_bb4_c0_ene123_0_reg_5_NO_SHIFT_REG;

// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_2to8_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to8_bb4_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to8_bb4_c0_ene2_0_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_2to8_bb4_c0_ene2_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_2to8_bb4_c0_ene2_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to8_bb4_c0_ene2_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to8_bb4_c0_ene2_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_2to8_bb4_c0_ene2_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_2to8_bb4_c0_ene2_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_2to8_bb4_c0_ene2_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.DEPTH = 6;
defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to8_bb4_c0_ene2_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_2to8_bb4_c0_ene2_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene2_0_NO_SHIFT_REG = rnode_2to8_bb4_c0_ene2_0_reg_8_NO_SHIFT_REG;
assign rnode_2to8_bb4_c0_ene2_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_2to8_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_2to5_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to5_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_2to5_bb4_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_2to5_bb4_c0_ene3_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_2to5_bb4_c0_ene3_0_reg_5_NO_SHIFT_REG;
 logic rnode_2to5_bb4_c0_ene3_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_2to5_bb4_c0_ene3_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_2to5_bb4_c0_ene3_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_2to5_bb4_c0_ene3_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to5_bb4_c0_ene3_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to5_bb4_c0_ene3_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_2to5_bb4_c0_ene3_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_2to5_bb4_c0_ene3_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_2to5_bb4_c0_ene3_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_2to5_bb4_c0_ene3_0_reg_5_fifo.DEPTH = 3;
defparam rnode_2to5_bb4_c0_ene3_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_2to5_bb4_c0_ene3_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to5_bb4_c0_ene3_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_2to5_bb4_c0_ene3_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to5_bb4_c0_ene3_0_NO_SHIFT_REG = rnode_2to5_bb4_c0_ene3_0_reg_5_NO_SHIFT_REG;
assign rnode_2to5_bb4_c0_ene3_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_2to5_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene4_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene4_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene4_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene4_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene4_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene4_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene4_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene4_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene4_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene4_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene4_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene4_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 7
//  * capacity = 7
 logic rnode_2to9_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_2to9_bb4_c0_ene5_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_2to9_bb4_c0_ene5_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to9_bb4_c0_ene5_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to9_bb4_c0_ene5_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_2to9_bb4_c0_ene5_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_2to9_bb4_c0_ene5_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_1to2_bb4_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_2to9_bb4_c0_ene5_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.DEPTH = 7;
defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to9_bb4_c0_ene5_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_2to9_bb4_c0_ene5_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_1to2_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene5_0_NO_SHIFT_REG = rnode_2to9_bb4_c0_ene5_0_reg_9_NO_SHIFT_REG;
assign rnode_2to9_bb4_c0_ene5_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_2to9_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_2_3_0_inputs_ready;
 reg SFC_2_VALID_2_3_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_2_3_0_stall_in_0;
 reg SFC_2_VALID_2_3_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_2_3_0_stall_in_1;
wire SFC_2_VALID_2_3_0_output_regs_ready;
 reg SFC_2_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_2_3_0_causedstall;

assign SFC_2_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_1_2_0_stall_in = 1'b0;
assign SFC_2_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_2_3_0_output_regs_ready)
		begin
			SFC_2_VALID_2_3_0_NO_SHIFT_REG <= SFC_2_VALID_1_2_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_i1_9_u17_stall_local;
wire local_bb4__acl_ffwd_dest_i1_9_u17;

assign local_bb4__acl_ffwd_dest_i1_9_u17 = ffwd_9_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_1_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_valid_out_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_stall_in_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene123_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb4_c0_ene123_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb4_c0_ene123_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb4_c0_ene123_0_stall_in_0_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb4_c0_ene123_0_valid_out_0_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb4_c0_ene123_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_3to5_bb4_c0_ene123_1_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb4_c0_ene123_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb4_c0_ene123_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb4_c0_ene123_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb4_c0_ene123_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb4_c0_ene123_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb4_c0_ene123_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to5_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_c0_ene123_0_stall_in_0_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_5to6_bb4_c0_ene123_0_NO_SHIFT_REG = rnode_5to6_bb4_c0_ene123_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_5to6_bb4_c0_ene123_1_NO_SHIFT_REG = rnode_5to6_bb4_c0_ene123_0_reg_6_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_c0_ene2_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene2_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_c0_ene2_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_c0_ene2_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_c0_ene2_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_c0_ene2_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_c0_ene2_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_2to8_bb4_c0_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_c0_ene2_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_c0_ene2_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_c0_ene2_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to8_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene2_0_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene2_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_c0_ene2_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb4_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene3_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb4_c0_ene3_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene3_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene3_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_c0_ene3_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb4_c0_ene3_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb4_c0_ene3_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb4_c0_ene3_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb4_c0_ene3_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb4_c0_ene3_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_2to5_bb4_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb4_c0_ene3_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb4_c0_ene3_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb4_c0_ene3_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb4_c0_ene3_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb4_c0_ene3_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb4_c0_ene3_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to5_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_c0_ene3_0_NO_SHIFT_REG = rnode_5to6_bb4_c0_ene3_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb4_c0_ene3_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene4_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene4_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene4_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene4_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene4_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene4_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene4_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene4_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene4_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene4_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene4_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene4_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene5_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene5_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene5_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene5_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene5_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene5_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_2to9_bb4_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene5_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene5_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene5_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to9_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene5_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene5_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene5_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_3_4_0_inputs_ready;
 reg SFC_2_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_3_4_0_stall_in;
wire SFC_2_VALID_3_4_0_output_regs_ready;
 reg SFC_2_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_3_4_0_causedstall;

assign SFC_2_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_2_3_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_3_4_0_output_regs_ready)
		begin
			SFC_2_VALID_3_4_0_NO_SHIFT_REG <= SFC_2_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_indvars_iv_pop7__stall_local;
wire [63:0] local_bb4_indvars_iv_pop7_;
wire local_bb4_indvars_iv_pop7__fu_valid_out;
wire local_bb4_indvars_iv_pop7__fu_stall_out;

acl_pop local_bb4_indvars_iv_pop7__feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_1to3_bb4_c0_ene123_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(input_wii_var_),
	.stall_out(local_bb4_indvars_iv_pop7__fu_stall_out),
	.valid_in(SFC_2_VALID_2_3_0_NO_SHIFT_REG),
	.valid_out(local_bb4_indvars_iv_pop7__fu_valid_out),
	.stall_in(local_bb4_indvars_iv_pop7__stall_local),
	.data_out(local_bb4_indvars_iv_pop7_),
	.feedback_in(feedback_data_in_7),
	.feedback_valid_in(feedback_valid_in_7),
	.feedback_stall_out(feedback_stall_out_7)
);

defparam local_bb4_indvars_iv_pop7__feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_indvars_iv_pop7__feedback.DATA_WIDTH = 64;
defparam local_bb4_indvars_iv_pop7__feedback.STYLE = "REGULAR";

assign local_bb4_indvars_iv_pop7__stall_local = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_c0_ene123_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene123_0_stall_in_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene123_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene123_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene123_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene123_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene123_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_c0_ene123_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_c0_ene123_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_c0_ene123_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_c0_ene123_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_c0_ene123_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_c0_ene123_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(rnode_5to6_bb4_c0_ene123_1_NO_SHIFT_REG),
	.data_out(rnode_6to7_bb4_c0_ene123_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_c0_ene123_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_c0_ene123_0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_6to7_bb4_c0_ene123_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_c0_ene123_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_c0_ene123_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_5to6_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene123_0_NO_SHIFT_REG = rnode_6to7_bb4_c0_ene123_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_c0_ene123_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_c0_ene123_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_4_5_0_inputs_ready;
 reg SFC_2_VALID_4_5_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_4_5_0_stall_in_0;
 reg SFC_2_VALID_4_5_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_4_5_0_stall_in_1;
wire SFC_2_VALID_4_5_0_output_regs_ready;
 reg SFC_2_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_4_5_0_causedstall;

assign SFC_2_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_3_4_0_stall_in = 1'b0;
assign SFC_2_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_4_5_0_output_regs_ready)
		begin
			SFC_2_VALID_4_5_0_NO_SHIFT_REG <= SFC_2_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__stall_local;
wire [31:0] local_bb4_var_;

assign local_bb4_var_ = local_bb4_indvars_iv_pop7_[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u18_stall_local;
wire [63:0] local_bb4_var__u18;

assign local_bb4_var__u18 = (local_bb4_indvars_iv_pop7_ + input_wii_var__u15);

// This section implements an unregistered operation.
// 
wire local_bb4_indvars_iv_next_stall_local;
wire [63:0] local_bb4_indvars_iv_next;

assign local_bb4_indvars_iv_next = (local_bb4_indvars_iv_pop7_ + 64'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_c0_ene123_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb4_c0_ene123_0_stall_in_NO_SHIFT_REG;
 logic rnode_7to8_bb4_c0_ene123_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_c0_ene123_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic rnode_7to8_bb4_c0_ene123_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_c0_ene123_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_c0_ene123_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_c0_ene123_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_c0_ene123_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_c0_ene123_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_c0_ene123_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_c0_ene123_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_c0_ene123_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_c0_ene123_0_NO_SHIFT_REG),
	.data_out(rnode_7to8_bb4_c0_ene123_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_c0_ene123_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_c0_ene123_0_reg_8_fifo.DATA_WIDTH = 1;
defparam rnode_7to8_bb4_c0_ene123_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_c0_ene123_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_c0_ene123_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_c0_ene123_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_c0_ene123_0_NO_SHIFT_REG = rnode_7to8_bb4_c0_ene123_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_c0_ene123_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_c0_ene123_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_5_6_0_inputs_ready;
 reg SFC_2_VALID_5_6_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_5_6_0_stall_in_0;
 reg SFC_2_VALID_5_6_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_5_6_0_stall_in_1;
wire SFC_2_VALID_5_6_0_output_regs_ready;
 reg SFC_2_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_5_6_0_causedstall;

assign SFC_2_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_4_5_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_5_6_0_output_regs_ready)
		begin
			SFC_2_VALID_5_6_0_NO_SHIFT_REG <= SFC_2_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_add26_stall_local;
wire [31:0] local_bb4_add26;

assign local_bb4_add26 = (local_bb4_var_ + local_bb4_pos_y_02_acl_ffwd_dest_i32_0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u18_valid_out;
wire local_bb4_var__u18_stall_in;
wire local_bb4_indvars_iv_next_valid_out_1;
wire local_bb4_indvars_iv_next_stall_in_1;
wire local_bb4_add26_valid_out;
wire local_bb4_add26_stall_in;
wire local_bb4_var__u19_valid_out;
wire local_bb4_var__u19_stall_in;
wire local_bb4_var__u19_inputs_ready;
wire local_bb4_var__u19_stall_local;
wire [31:0] local_bb4_var__u19;

assign local_bb4_var__u19_inputs_ready = (SFC_2_VALID_2_3_0_valid_out_1_NO_SHIFT_REG & rnode_1to3_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG & rnode_1to3_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_var__u19 = local_bb4_indvars_iv_next[31:0];
assign local_bb4_var__u18_valid_out = 1'b1;
assign local_bb4_indvars_iv_next_valid_out_1 = 1'b1;
assign local_bb4_add26_valid_out = 1'b1;
assign local_bb4_var__u19_valid_out = 1'b1;
assign SFC_2_VALID_2_3_0_stall_in_1 = 1'b0;
assign rnode_1to3_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_1to3_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_2_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_valid_out_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_stall_in_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_c0_ene123_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_c0_ene123_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_c0_ene123_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_c0_ene123_0_stall_in_0_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_c0_ene123_0_valid_out_0_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_c0_ene123_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_7to8_bb4_c0_ene123_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_c0_ene123_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_c0_ene123_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_c0_ene123_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_c0_ene123_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_c0_ene123_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_c0_ene123_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_c0_ene123_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene123_0_stall_in_0_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_c0_ene123_0_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene123_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_c0_ene123_1_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene123_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_c0_ene123_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_c0_ene123_2_NO_SHIFT_REG = rnode_8to9_bb4_c0_ene123_0_reg_9_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_2_VALID_6_7_0_inputs_ready;
 reg SFC_2_VALID_6_7_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_6_7_0_stall_in;
wire SFC_2_VALID_6_7_0_output_regs_ready;
 reg SFC_2_VALID_6_7_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_6_7_0_causedstall;

assign SFC_2_VALID_6_7_0_inputs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_5_6_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_6_7_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_6_7_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_6_7_0_output_regs_ready)
		begin
			SFC_2_VALID_6_7_0_NO_SHIFT_REG <= SFC_2_VALID_5_6_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_gaussian_ROM4119_pop11_c0_ene3_stall_local;
wire [31:0] local_bb4_gaussian_ROM4119_pop11_c0_ene3;
wire local_bb4_gaussian_ROM4119_pop11_c0_ene3_fu_valid_out;
wire local_bb4_gaussian_ROM4119_pop11_c0_ene3_fu_stall_out;

acl_pop local_bb4_gaussian_ROM4119_pop11_c0_ene3_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_5to6_bb4_c0_ene123_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_5to6_bb4_c0_ene3_0_NO_SHIFT_REG),
	.stall_out(local_bb4_gaussian_ROM4119_pop11_c0_ene3_fu_stall_out),
	.valid_in(SFC_2_VALID_5_6_0_NO_SHIFT_REG),
	.valid_out(local_bb4_gaussian_ROM4119_pop11_c0_ene3_fu_valid_out),
	.stall_in(local_bb4_gaussian_ROM4119_pop11_c0_ene3_stall_local),
	.data_out(local_bb4_gaussian_ROM4119_pop11_c0_ene3),
	.feedback_in(feedback_data_in_11),
	.feedback_valid_in(feedback_valid_in_11),
	.feedback_stall_out(feedback_stall_out_11)
);

defparam local_bb4_gaussian_ROM4119_pop11_c0_ene3_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_gaussian_ROM4119_pop11_c0_ene3_feedback.DATA_WIDTH = 32;
defparam local_bb4_gaussian_ROM4119_pop11_c0_ene3_feedback.STYLE = "REGULAR";

assign local_bb4_gaussian_ROM4119_pop11_c0_ene3_stall_local = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb4_var__u18_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u18_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_3to4_bb4_var__u18_0_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u18_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_3to4_bb4_var__u18_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u18_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u18_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u18_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb4_var__u18_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb4_var__u18_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb4_var__u18_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb4_var__u18_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb4_var__u18_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb4_var__u18),
	.data_out(rnode_3to4_bb4_var__u18_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb4_var__u18_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb4_var__u18_0_reg_4_fifo.DATA_WIDTH = 64;
defparam rnode_3to4_bb4_var__u18_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb4_var__u18_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb4_var__u18_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u18_stall_in = 1'b0;
assign rnode_3to4_bb4_var__u18_0_NO_SHIFT_REG = rnode_3to4_bb4_var__u18_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb4_var__u18_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb4_var__u18_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb4_indvars_iv_next_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to5_bb4_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_3to5_bb4_indvars_iv_next_0_NO_SHIFT_REG;
 logic rnode_3to5_bb4_indvars_iv_next_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_3to5_bb4_indvars_iv_next_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_indvars_iv_next_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_indvars_iv_next_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_indvars_iv_next_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb4_indvars_iv_next_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb4_indvars_iv_next_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb4_indvars_iv_next_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb4_indvars_iv_next_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb4_indvars_iv_next_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb4_indvars_iv_next),
	.data_out(rnode_3to5_bb4_indvars_iv_next_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb4_indvars_iv_next_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb4_indvars_iv_next_0_reg_5_fifo.DATA_WIDTH = 64;
defparam rnode_3to5_bb4_indvars_iv_next_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb4_indvars_iv_next_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb4_indvars_iv_next_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_indvars_iv_next_stall_in_1 = 1'b0;
assign rnode_3to5_bb4_indvars_iv_next_0_NO_SHIFT_REG = rnode_3to5_bb4_indvars_iv_next_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb4_indvars_iv_next_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb4_indvars_iv_next_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_3to5_bb4_add26_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_3to5_bb4_add26_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_3to5_bb4_add26_0_NO_SHIFT_REG;
 logic rnode_3to5_bb4_add26_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_3to5_bb4_add26_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_3to5_bb4_add26_1_NO_SHIFT_REG;
 logic rnode_3to5_bb4_add26_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to5_bb4_add26_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_add26_0_valid_out_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_add26_0_stall_in_0_reg_5_NO_SHIFT_REG;
 logic rnode_3to5_bb4_add26_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_3to5_bb4_add26_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to5_bb4_add26_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to5_bb4_add26_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_3to5_bb4_add26_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_3to5_bb4_add26_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb4_add26),
	.data_out(rnode_3to5_bb4_add26_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_3to5_bb4_add26_0_reg_5_fifo.DEPTH = 2;
defparam rnode_3to5_bb4_add26_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_3to5_bb4_add26_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to5_bb4_add26_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_3to5_bb4_add26_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add26_stall_in = 1'b0;
assign rnode_3to5_bb4_add26_0_stall_in_0_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_3to5_bb4_add26_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_3to5_bb4_add26_0_NO_SHIFT_REG = rnode_3to5_bb4_add26_0_reg_5_NO_SHIFT_REG;
assign rnode_3to5_bb4_add26_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_3to5_bb4_add26_1_NO_SHIFT_REG = rnode_3to5_bb4_add26_0_reg_5_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_3to4_bb4_var__u19_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u19_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb4_var__u19_0_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u19_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_3to4_bb4_var__u19_0_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u19_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u19_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_3to4_bb4_var__u19_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_3to4_bb4_var__u19_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to4_bb4_var__u19_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to4_bb4_var__u19_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_3to4_bb4_var__u19_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_3to4_bb4_var__u19_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb4_var__u19),
	.data_out(rnode_3to4_bb4_var__u19_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_3to4_bb4_var__u19_0_reg_4_fifo.DEPTH = 1;
defparam rnode_3to4_bb4_var__u19_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_3to4_bb4_var__u19_0_reg_4_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to4_bb4_var__u19_0_reg_4_fifo.IMPL = "shift_reg";

assign rnode_3to4_bb4_var__u19_0_reg_4_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u19_stall_in = 1'b0;
assign rnode_3to4_bb4_var__u19_0_NO_SHIFT_REG = rnode_3to4_bb4_var__u19_0_reg_4_NO_SHIFT_REG;
assign rnode_3to4_bb4_var__u19_0_stall_in_reg_4_NO_SHIFT_REG = 1'b0;
assign rnode_3to4_bb4_var__u19_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_valid_out_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_stall_in_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_c0_ene123_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_c0_ene123_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_c0_ene123_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_c0_ene123_0_stall_in_0_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_c0_ene123_0_valid_out_0_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_c0_ene123_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_8to9_bb4_c0_ene123_2_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_c0_ene123_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_c0_ene123_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_c0_ene123_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_9to10_bb4_c0_ene123_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_c0_ene123_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_c0_ene123_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_c0_ene123_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene123_0_stall_in_0_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene123_0_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene123_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4_c0_ene123_1_NO_SHIFT_REG = rnode_9to10_bb4_c0_ene123_0_reg_10_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_2_VALID_7_8_0_inputs_ready;
 reg SFC_2_VALID_7_8_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_7_8_0_stall_in;
wire SFC_2_VALID_7_8_0_output_regs_ready;
 reg SFC_2_VALID_7_8_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_7_8_0_causedstall;

assign SFC_2_VALID_7_8_0_inputs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_6_7_0_stall_in = 1'b0;
assign SFC_2_VALID_7_8_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_7_8_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_7_8_0_output_regs_ready)
		begin
			SFC_2_VALID_7_8_0_NO_SHIFT_REG <= SFC_2_VALID_6_7_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u20_stall_local;
wire [31:0] local_bb4_var__u20;

assign local_bb4_var__u20 = local_bb4_gaussian_ROM4119_pop11_c0_ene3;

// This section implements a registered operation.
// 
wire local_bb4_arrayidx44_inputs_ready;
 reg local_bb4_arrayidx44_valid_out_NO_SHIFT_REG;
wire local_bb4_arrayidx44_stall_in;
wire local_bb4_arrayidx44_output_regs_ready;
 reg [63:0] local_bb4_arrayidx44_NO_SHIFT_REG;
wire [63:0] local_bb4_arrayidx44_op_wire;
wire local_bb4_arrayidx44_causedstall;

assign local_bb4_arrayidx44_inputs_ready = 1'b1;
assign local_bb4_arrayidx44_output_regs_ready = 1'b1;
assign local_bb4_arrayidx44_op_wire = (64'h0 + (rnode_3to4_bb4_var__u18_0_NO_SHIFT_REG << 6'h2));
assign rnode_3to4_bb4_var__u18_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_arrayidx44_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_arrayidx44_NO_SHIFT_REG <= 'x;
		local_bb4_arrayidx44_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_arrayidx44_output_regs_ready)
		begin
			local_bb4_arrayidx44_NO_SHIFT_REG <= local_bb4_arrayidx44_op_wire;
			local_bb4_arrayidx44_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_arrayidx44_stall_in))
			begin
				local_bb4_arrayidx44_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_cmp1_i5_valid_out;
wire local_bb4_cmp1_i5_stall_in;
wire local_bb4_cmp1_i5_inputs_ready;
wire local_bb4_cmp1_i5_stall_local;
wire local_bb4_cmp1_i5;

assign local_bb4_cmp1_i5_inputs_ready = rnode_3to5_bb4_add26_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_cmp1_i5 = (rnode_3to5_bb4_add26_0_NO_SHIFT_REG > input_wii_sub27);
assign local_bb4_cmp1_i5_valid_out = 1'b1;
assign rnode_3to5_bb4_add26_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb4_add26_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb4_add26_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb4_add26_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_add26_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_5to6_bb4_add26_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_add26_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_add26_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_add26_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb4_add26_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb4_add26_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb4_add26_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb4_add26_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb4_add26_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(rnode_3to5_bb4_add26_1_NO_SHIFT_REG),
	.data_out(rnode_5to6_bb4_add26_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb4_add26_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb4_add26_0_reg_6_fifo.DATA_WIDTH = 32;
defparam rnode_5to6_bb4_add26_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb4_add26_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb4_add26_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to5_bb4_add26_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_add26_0_NO_SHIFT_REG = rnode_5to6_bb4_add26_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb4_add26_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_add26_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp20_valid_out;
wire local_bb4_cmp20_stall_in;
wire local_bb4_cmp20_inputs_ready;
wire local_bb4_cmp20_stall_local;
wire local_bb4_cmp20;

assign local_bb4_cmp20_inputs_ready = rnode_3to4_bb4_var__u19_0_valid_out_NO_SHIFT_REG;
assign local_bb4_cmp20 = ($signed(rnode_3to4_bb4_var__u19_0_NO_SHIFT_REG) > $signed(input_r));
assign local_bb4_cmp20_valid_out = 1'b1;
assign rnode_3to4_bb4_var__u19_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_2_VALID_8_9_0_inputs_ready;
 reg SFC_2_VALID_8_9_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_0;
 reg SFC_2_VALID_8_9_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_1;
 reg SFC_2_VALID_8_9_0_valid_out_2_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_2;
 reg SFC_2_VALID_8_9_0_valid_out_3_NO_SHIFT_REG;
wire SFC_2_VALID_8_9_0_stall_in_3;
wire SFC_2_VALID_8_9_0_output_regs_ready;
 reg SFC_2_VALID_8_9_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_8_9_0_causedstall;

assign SFC_2_VALID_8_9_0_inputs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_7_8_0_stall_in = 1'b0;
assign SFC_2_VALID_8_9_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_8_9_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_8_9_0_output_regs_ready)
		begin
			SFC_2_VALID_8_9_0_NO_SHIFT_REG <= SFC_2_VALID_7_8_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr_i410_stall_local;
wire [31:0] local_bb4_shr_i410;

assign local_bb4_shr_i410 = (local_bb4_var__u20 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and5_i416_stall_local;
wire [31:0] local_bb4_and5_i416;

assign local_bb4_and5_i416 = (local_bb4_var__u20 & 32'h7FFFFF);

// This section implements a registered operation.
// 
// Filescope constant lowered to ROM: gaussian.ROM
wire local_bb4_gaussian_ROM_arrayidx44_inputs_ready;
 reg local_bb4_gaussian_ROM_arrayidx44_valid_out_NO_SHIFT_REG;
wire local_bb4_gaussian_ROM_arrayidx44_stall_in;
wire local_bb4_gaussian_ROM_arrayidx44_output_regs_ready;
 reg [31:0] local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG;
wire [63:0] local_bb4_gaussian_ROM_arrayidx44$addr$ps;
wire local_bb4_gaussian_ROM_arrayidx44_causedstall;

assign local_bb4_gaussian_ROM_arrayidx44_inputs_ready = 1'b1;
assign local_bb4_gaussian_ROM_arrayidx44_output_regs_ready = 1'b1;
assign local_bb4_gaussian_ROM_arrayidx44$addr$ps = (local_bb4_arrayidx44_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign local_bb4_arrayidx44_stall_in = 1'b0;
assign local_bb4_gaussian_ROM_arrayidx44_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (local_bb4_gaussian_ROM_arrayidx44_output_regs_ready)
		begin
			case (local_bb4_gaussian_ROM_arrayidx44$addr$ps[4:2])
				3'h0:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h3F61EB85;
				end

				3'h1:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h3F781D7E;
				end

				3'h2:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h3F800000;
				end

				3'h3:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h3F781D7E;
				end

				3'h4:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h3F61EB85;
				end

				3'h5:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h3F413A93;
				end

				3'h6:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h0;
				end

				3'h7:
				begin
					local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG <= 32'h0;
				end

				default:
				begin
				end

			endcase
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_gaussian_ROM_arrayidx44_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_gaussian_ROM_arrayidx44_output_regs_ready)
		begin
			local_bb4_gaussian_ROM_arrayidx44_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_gaussian_ROM_arrayidx44_stall_in))
			begin
				local_bb4_gaussian_ROM_arrayidx44_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb4_cmp1_i5_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb4_cmp1_i5_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb4_cmp1_i5_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_cmp1_i5_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb4_cmp1_i5_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_cmp1_i5_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_cmp1_i5_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_cmp1_i5_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb4_cmp1_i5_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb4_cmp1_i5_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb4_cmp1_i5_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb4_cmp1_i5_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb4_cmp1_i5_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb4_cmp1_i5),
	.data_out(rnode_5to6_bb4_cmp1_i5_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb4_cmp1_i5_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb4_cmp1_i5_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb4_cmp1_i5_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb4_cmp1_i5_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb4_cmp1_i5_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp1_i5_stall_in = 1'b0;
assign rnode_5to6_bb4_cmp1_i5_0_NO_SHIFT_REG = rnode_5to6_bb4_cmp1_i5_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb4_cmp1_i5_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_cmp1_i5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb4_cmp20_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb4_cmp20_0_stall_in_NO_SHIFT_REG;
 logic rnode_4to5_bb4_cmp20_0_NO_SHIFT_REG;
 logic rnode_4to5_bb4_cmp20_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_4to5_bb4_cmp20_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb4_cmp20_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb4_cmp20_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb4_cmp20_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb4_cmp20_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb4_cmp20_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb4_cmp20_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb4_cmp20_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb4_cmp20_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb4_cmp20),
	.data_out(rnode_4to5_bb4_cmp20_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb4_cmp20_0_reg_5_fifo.DEPTH = 1;
defparam rnode_4to5_bb4_cmp20_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_4to5_bb4_cmp20_0_reg_5_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_4to5_bb4_cmp20_0_reg_5_fifo.IMPL = "shift_reg";

assign rnode_4to5_bb4_cmp20_0_reg_5_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp20_stall_in = 1'b0;
assign rnode_4to5_bb4_cmp20_0_NO_SHIFT_REG = rnode_4to5_bb4_cmp20_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb4_cmp20_0_stall_in_reg_5_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb4_cmp20_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_2_VALID_9_10_0_inputs_ready;
 reg SFC_2_VALID_9_10_0_valid_out_0_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_0;
 reg SFC_2_VALID_9_10_0_valid_out_1_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_1;
 reg SFC_2_VALID_9_10_0_valid_out_2_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_2;
 reg SFC_2_VALID_9_10_0_valid_out_3_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_3;
 reg SFC_2_VALID_9_10_0_valid_out_4_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_4;
 reg SFC_2_VALID_9_10_0_valid_out_5_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_5;
 reg SFC_2_VALID_9_10_0_valid_out_6_NO_SHIFT_REG;
wire SFC_2_VALID_9_10_0_stall_in_6;
wire SFC_2_VALID_9_10_0_output_regs_ready;
 reg SFC_2_VALID_9_10_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_9_10_0_causedstall;

assign SFC_2_VALID_9_10_0_inputs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_9_10_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_9_10_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_9_10_0_output_regs_ready)
		begin
			SFC_2_VALID_9_10_0_NO_SHIFT_REG <= SFC_2_VALID_8_9_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_keep_going_acl_pipeline_1_inputs_ready;
 reg local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG;
wire local_bb4_keep_going_acl_pipeline_1_stall_in;
wire local_bb4_keep_going_acl_pipeline_1_output_regs_ready;
wire local_bb4_keep_going_acl_pipeline_1_keep_going;
wire local_bb4_keep_going_acl_pipeline_1_fu_valid_out;
wire local_bb4_keep_going_acl_pipeline_1_fu_stall_out;
 reg local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG;
wire local_bb4_keep_going_acl_pipeline_1_feedback_pipelined;
wire local_bb4_keep_going_acl_pipeline_1_causedstall;

acl_pipeline local_bb4_keep_going_acl_pipeline_1_pipelined (
	.clock(clock),
	.resetn(resetn),
	.data_in(1'b1),
	.stall_out(local_bb4_keep_going_acl_pipeline_1_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_keep_going_acl_pipeline_1_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_keep_going_acl_pipeline_1_keep_going),
	.initeration_in(1'b0),
	.initeration_valid_in(1'b0),
	.initeration_stall_out(feedback_stall_out_0),
	.not_exitcond_in(feedback_data_in_1),
	.not_exitcond_valid_in(feedback_valid_in_1),
	.not_exitcond_stall_out(feedback_stall_out_1),
	.pipeline_valid_out(acl_pipelined_valid),
	.pipeline_stall_in(acl_pipelined_stall),
	.exiting_valid_out(acl_pipelined_exiting_valid)
);

defparam local_bb4_keep_going_acl_pipeline_1_pipelined.FIFO_DEPTH = 0;
defparam local_bb4_keep_going_acl_pipeline_1_pipelined.STYLE = "NON_SPECULATIVE";

assign local_bb4_keep_going_acl_pipeline_1_inputs_ready = 1'b1;
assign local_bb4_keep_going_acl_pipeline_1_output_regs_ready = 1'b1;
assign acl_pipelined_exiting_stall = acl_pipelined_stall;
assign SFC_2_VALID_8_9_0_stall_in_1 = 1'b0;
assign rnode_8to9_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb4_keep_going_acl_pipeline_1_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG <= 'x;
		local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_keep_going_acl_pipeline_1_output_regs_ready)
		begin
			local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG <= local_bb4_keep_going_acl_pipeline_1_keep_going;
			local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_keep_going_acl_pipeline_1_stall_in))
			begin
				local_bb4_keep_going_acl_pipeline_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_sub24_add2318_pop10_c0_ene2_stall_local;
wire [31:0] local_bb4_sub24_add2318_pop10_c0_ene2;
wire local_bb4_sub24_add2318_pop10_c0_ene2_fu_valid_out;
wire local_bb4_sub24_add2318_pop10_c0_ene2_fu_stall_out;

acl_pop local_bb4_sub24_add2318_pop10_c0_ene2_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_8to9_bb4_c0_ene123_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_8to9_bb4_c0_ene2_0_NO_SHIFT_REG),
	.stall_out(local_bb4_sub24_add2318_pop10_c0_ene2_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sub24_add2318_pop10_c0_ene2_fu_valid_out),
	.stall_in(local_bb4_sub24_add2318_pop10_c0_ene2_stall_local),
	.data_out(local_bb4_sub24_add2318_pop10_c0_ene2),
	.feedback_in(feedback_data_in_10),
	.feedback_valid_in(feedback_valid_in_10),
	.feedback_stall_out(feedback_stall_out_10)
);

defparam local_bb4_sub24_add2318_pop10_c0_ene2_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_sub24_add2318_pop10_c0_ene2_feedback.DATA_WIDTH = 32;
defparam local_bb4_sub24_add2318_pop10_c0_ene2_feedback.STYLE = "REGULAR";

assign local_bb4_sub24_add2318_pop10_c0_ene2_stall_local = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i411_stall_local;
wire [31:0] local_bb4_and_i411;

assign local_bb4_and_i411 = ((local_bb4_shr_i410 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i422_stall_local;
wire local_bb4_lnot14_i422;

assign local_bb4_lnot14_i422 = ((local_bb4_and5_i416 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i444_stall_local;
wire [31:0] local_bb4_or_i444;

assign local_bb4_or_i444 = ((local_bb4_and5_i416 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u21_stall_local;
wire [31:0] local_bb4_var__u21;

assign local_bb4_var__u21 = local_bb4_gaussian_ROM_arrayidx44_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_sub27_add26_valid_out;
wire local_bb4_sub27_add26_stall_in;
wire local_bb4_sub27_add26_inputs_ready;
wire local_bb4_sub27_add26_stall_local;
wire [31:0] local_bb4_sub27_add26;

assign local_bb4_sub27_add26_inputs_ready = (rnode_5to6_bb4_cmp1_i5_0_valid_out_NO_SHIFT_REG & rnode_5to6_bb4_add26_0_valid_out_NO_SHIFT_REG);
assign local_bb4_sub27_add26 = (rnode_5to6_bb4_cmp1_i5_0_NO_SHIFT_REG ? input_wii_sub27 : rnode_5to6_bb4_add26_0_NO_SHIFT_REG);
assign local_bb4_sub27_add26_valid_out = 1'b1;
assign rnode_5to6_bb4_cmp1_i5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_add26_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u22_stall_local;
wire local_bb4_var__u22;

assign local_bb4_var__u22 = (local_bb4__acl_ffwd_dest_i1_9_u17 | rnode_4to5_bb4_cmp20_0_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_2_VALID_10_11_0_inputs_ready;
 reg SFC_2_VALID_10_11_0_valid_out_NO_SHIFT_REG;
wire SFC_2_VALID_10_11_0_stall_in;
wire SFC_2_VALID_10_11_0_output_regs_ready;
 reg SFC_2_VALID_10_11_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_2_VALID_10_11_0_causedstall;

assign SFC_2_VALID_10_11_0_inputs_ready = 1'b1;
assign SFC_2_VALID_10_11_0_output_regs_ready = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_0 = 1'b0;
assign SFC_2_VALID_10_11_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_2_VALID_10_11_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_2_VALID_10_11_0_output_regs_ready)
		begin
			SFC_2_VALID_10_11_0_NO_SHIFT_REG <= SFC_2_VALID_9_10_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__pop12_c0_ene4_valid_out_0;
wire local_bb4__pop12_c0_ene4_stall_in_0;
wire local_bb4__pop12_c0_ene4_valid_out_1;
wire local_bb4__pop12_c0_ene4_stall_in_1;
wire local_bb4__pop12_c0_ene4_inputs_ready;
wire local_bb4__pop12_c0_ene4_stall_local;
wire local_bb4__pop12_c0_ene4;
wire local_bb4__pop12_c0_ene4_fu_valid_out;
wire local_bb4__pop12_c0_ene4_fu_stall_out;

acl_pop local_bb4__pop12_c0_ene4_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene123_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene4_0_NO_SHIFT_REG),
	.stall_out(local_bb4__pop12_c0_ene4_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__pop12_c0_ene4_fu_valid_out),
	.stall_in(local_bb4__pop12_c0_ene4_stall_local),
	.data_out(local_bb4__pop12_c0_ene4),
	.feedback_in(feedback_data_in_12),
	.feedback_valid_in(feedback_valid_in_12),
	.feedback_stall_out(feedback_stall_out_12)
);

defparam local_bb4__pop12_c0_ene4_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4__pop12_c0_ene4_feedback.DATA_WIDTH = 1;
defparam local_bb4__pop12_c0_ene4_feedback.STYLE = "REGULAR";

assign local_bb4__pop12_c0_ene4_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_1_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene4_0_valid_out_NO_SHIFT_REG);
assign local_bb4__pop12_c0_ene4_stall_local = 1'b0;
assign local_bb4__pop12_c0_ene4_valid_out_0 = 1'b1;
assign local_bb4__pop12_c0_ene4_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_1 = 1'b0;
assign rnode_9to10_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notexitcond1520_pop13_c0_ene5_valid_out_0;
wire local_bb4_notexitcond1520_pop13_c0_ene5_stall_in_0;
wire local_bb4_notexitcond1520_pop13_c0_ene5_valid_out_1;
wire local_bb4_notexitcond1520_pop13_c0_ene5_stall_in_1;
wire local_bb4_notexitcond1520_pop13_c0_ene5_inputs_ready;
wire local_bb4_notexitcond1520_pop13_c0_ene5_stall_local;
wire local_bb4_notexitcond1520_pop13_c0_ene5;
wire local_bb4_notexitcond1520_pop13_c0_ene5_fu_valid_out;
wire local_bb4_notexitcond1520_pop13_c0_ene5_fu_stall_out;

acl_pop local_bb4_notexitcond1520_pop13_c0_ene5_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_9to10_bb4_c0_ene123_1_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_c0_ene5_0_NO_SHIFT_REG),
	.stall_out(local_bb4_notexitcond1520_pop13_c0_ene5_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond1520_pop13_c0_ene5_fu_valid_out),
	.stall_in(local_bb4_notexitcond1520_pop13_c0_ene5_stall_local),
	.data_out(local_bb4_notexitcond1520_pop13_c0_ene5),
	.feedback_in(feedback_data_in_13),
	.feedback_valid_in(feedback_valid_in_13),
	.feedback_stall_out(feedback_stall_out_13)
);

defparam local_bb4_notexitcond1520_pop13_c0_ene5_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_notexitcond1520_pop13_c0_ene5_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond1520_pop13_c0_ene5_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond1520_pop13_c0_ene5_inputs_ready = (SFC_2_VALID_9_10_0_valid_out_2_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG & rnode_9to10_bb4_c0_ene5_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notexitcond1520_pop13_c0_ene5_stall_local = 1'b0;
assign local_bb4_notexitcond1520_pop13_c0_ene5_valid_out_0 = 1'b1;
assign local_bb4_notexitcond1520_pop13_c0_ene5_valid_out_1 = 1'b1;
assign SFC_2_VALID_9_10_0_stall_in_2 = 1'b0;
assign rnode_9to10_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_keep_going_acl_pipeline_1_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_keep_going_acl_pipeline_1_stall_in = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_NO_SHIFT_REG = rnode_10to11_bb4_keep_going_acl_pipeline_1_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i418_stall_local;
wire local_bb4_lnot_i418;

assign local_bb4_lnot_i418 = ((local_bb4_and_i411 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i420_stall_local;
wire local_bb4_cmp_i420;

assign local_bb4_cmp_i420 = ((local_bb4_and_i411 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_not_i441_stall_local;
wire local_bb4_lnot14_not_i441;

assign local_bb4_lnot14_not_i441 = (local_bb4_lnot14_i422 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_conv_i_i446_stall_local;
wire [63:0] local_bb4_conv_i_i446;

assign local_bb4_conv_i_i446[63:32] = 32'h0;
assign local_bb4_conv_i_i446[31:0] = ((local_bb4_or_i444 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i412_stall_local;
wire [31:0] local_bb4_shr2_i412;

assign local_bb4_shr2_i412 = (local_bb4_var__u21 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i414_stall_local;
wire [31:0] local_bb4_xor_i414;

assign local_bb4_xor_i414 = (local_bb4_var__u21 ^ local_bb4_var__u20);

// This section implements an unregistered operation.
// 
wire local_bb4_and6_i417_stall_local;
wire [31:0] local_bb4_and6_i417;

assign local_bb4_and6_i417 = (local_bb4_var__u21 & 32'h7FFFFF);

// This section implements a registered operation.
// 
wire local_bb4_mul30_inputs_ready;
 reg local_bb4_mul30_valid_out_NO_SHIFT_REG;
wire local_bb4_mul30_stall_in;
wire local_bb4_mul30_output_regs_ready;
wire [31:0] local_bb4_mul30;
 reg local_bb4_mul30_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul30_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul30_causedstall;

acl_int_mult int_module_local_bb4_mul30 (
	.clock(clock),
	.dataa(local_bb4_sub27_add26),
	.datab(input_global_size_0),
	.enable(local_bb4_mul30_output_regs_ready),
	.result(local_bb4_mul30)
);

defparam int_module_local_bb4_mul30.INPUT1_WIDTH = 32;
defparam int_module_local_bb4_mul30.INPUT2_WIDTH = 32;
defparam int_module_local_bb4_mul30.OUTPUT_WIDTH = 32;
defparam int_module_local_bb4_mul30.LATENCY = 3;
defparam int_module_local_bb4_mul30.SIGNED = 0;

assign local_bb4_mul30_inputs_ready = 1'b1;
assign local_bb4_mul30_output_regs_ready = 1'b1;
assign local_bb4_sub27_add26_stall_in = 1'b0;
assign local_bb4_mul30_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul30_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul30_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul30_output_regs_ready)
		begin
			local_bb4_mul30_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul30_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul30_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul30_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul30_output_regs_ready)
		begin
			local_bb4_mul30_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul30_stall_in))
			begin
				local_bb4_mul30_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u22_valid_out_1;
wire local_bb4_var__u22_stall_in_1;
wire local_bb4_notexit_valid_out_0;
wire local_bb4_notexit_stall_in_0;
wire local_bb4_notexit_valid_out_1;
wire local_bb4_notexit_stall_in_1;
wire local_bb4_notexit_inputs_ready;
wire local_bb4_notexit_stall_local;
wire local_bb4_notexit;

assign local_bb4_notexit_inputs_ready = (rnode_3to5_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG & rnode_4to5_bb4_cmp20_0_valid_out_NO_SHIFT_REG);
assign local_bb4_notexit = (local_bb4_var__u22 ^ 1'b1);
assign local_bb4_var__u22_valid_out_1 = 1'b1;
assign local_bb4_notexit_valid_out_0 = 1'b1;
assign local_bb4_notexit_valid_out_1 = 1'b1;
assign rnode_3to5_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_4to5_bb4_cmp20_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__pop12_c0_ene4_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4__pop12_c0_ene4_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4__pop12_c0_ene4),
	.data_out(rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__pop12_c0_ene4_stall_in_1 = 1'b0;
assign rnode_10to11_bb4__pop12_c0_ene4_0_NO_SHIFT_REG = rnode_10to11_bb4__pop12_c0_ene4_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond1520_pop13_c0_ene5),
	.data_out(rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond1520_pop13_c0_ene5_stall_in_1 = 1'b0;
assign rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_NO_SHIFT_REG = rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__28_i442_stall_local;
wire local_bb4__28_i442;

assign local_bb4__28_i442 = (local_bb4_cmp_i420 & local_bb4_lnot14_not_i441);

// This section implements an unregistered operation.
// 
wire local_bb4_and3_i413_stall_local;
wire [31:0] local_bb4_and3_i413;

assign local_bb4_and3_i413 = ((local_bb4_shr2_i412 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_i423_stall_local;
wire local_bb4_lnot17_i423;

assign local_bb4_lnot17_i423 = ((local_bb4_and6_i417 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u23_stall_local;
wire [31:0] local_bb4_var__u23;

assign local_bb4_var__u23 = ((local_bb4_and6_i417 & 32'h7FFFFF) | (local_bb4_and_i411 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_or47_i445_stall_local;
wire [31:0] local_bb4_or47_i445;

assign local_bb4_or47_i445 = ((local_bb4_and6_i417 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_sub24_add2318_pop10_c0_ene2_valid_out_1;
wire local_bb4_sub24_add2318_pop10_c0_ene2_stall_in_1;
wire local_bb4_add31_valid_out;
wire local_bb4_add31_stall_in;
wire local_bb4_add31_inputs_ready;
wire local_bb4_add31_stall_local;
wire [31:0] local_bb4_add31;

assign local_bb4_add31_inputs_ready = (SFC_2_VALID_8_9_0_valid_out_2_NO_SHIFT_REG & rnode_8to9_bb4_c0_ene2_0_valid_out_NO_SHIFT_REG & rnode_8to9_bb4_c0_ene123_0_valid_out_1_NO_SHIFT_REG & local_bb4_mul30_valid_out_NO_SHIFT_REG);
assign local_bb4_add31 = (local_bb4_mul30 + local_bb4_sub24_add2318_pop10_c0_ene2);
assign local_bb4_sub24_add2318_pop10_c0_ene2_valid_out_1 = 1'b1;
assign local_bb4_add31_valid_out = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in_2 = 1'b0;
assign rnode_8to9_bb4_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_c0_ene123_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign local_bb4_mul30_stall_in = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb4_var__u22_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb4_var__u22_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb4_var__u22_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_var__u22_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb4_var__u22_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_var__u22_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_var__u22_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_var__u22_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb4_var__u22_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb4_var__u22_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb4_var__u22_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb4_var__u22_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb4_var__u22_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb4_var__u22),
	.data_out(rnode_5to6_bb4_var__u22_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb4_var__u22_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb4_var__u22_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb4_var__u22_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb4_var__u22_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb4_var__u22_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u22_stall_in_1 = 1'b0;
assign rnode_5to6_bb4_var__u22_0_NO_SHIFT_REG = rnode_5to6_bb4_var__u22_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb4_var__u22_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_var__u22_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_indvars_iv_push7_indvars_iv_next_inputs_ready;
 reg local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG;
wire local_bb4_indvars_iv_push7_indvars_iv_next_stall_in;
wire local_bb4_indvars_iv_push7_indvars_iv_next_output_regs_ready;
wire [63:0] local_bb4_indvars_iv_push7_indvars_iv_next_result;
wire local_bb4_indvars_iv_push7_indvars_iv_next_fu_valid_out;
wire local_bb4_indvars_iv_push7_indvars_iv_next_fu_stall_out;
 reg [63:0] local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG;
wire local_bb4_indvars_iv_push7_indvars_iv_next_causedstall;

acl_push local_bb4_indvars_iv_push7_indvars_iv_next_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexit),
	.predicate(1'b0),
	.data_in(rnode_3to5_bb4_indvars_iv_next_0_NO_SHIFT_REG),
	.stall_out(local_bb4_indvars_iv_push7_indvars_iv_next_fu_stall_out),
	.valid_in(SFC_2_VALID_4_5_0_NO_SHIFT_REG),
	.valid_out(local_bb4_indvars_iv_push7_indvars_iv_next_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_indvars_iv_push7_indvars_iv_next_result),
	.feedback_out(feedback_data_out_7),
	.feedback_valid_out(feedback_valid_out_7),
	.feedback_stall_in(feedback_stall_in_7)
);

defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.STALLFREE = 1;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.DATA_WIDTH = 64;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.FIFO_DEPTH = 9;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.MIN_FIFO_LATENCY = 7;
defparam local_bb4_indvars_iv_push7_indvars_iv_next_feedback.STYLE = "REGULAR";

assign local_bb4_indvars_iv_push7_indvars_iv_next_inputs_ready = 1'b1;
assign local_bb4_indvars_iv_push7_indvars_iv_next_output_regs_ready = 1'b1;
assign local_bb4_notexit_stall_in_0 = 1'b0;
assign SFC_2_VALID_4_5_0_stall_in_1 = 1'b0;
assign rnode_3to5_bb4_indvars_iv_next_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_indvars_iv_push7_indvars_iv_next_causedstall = (SFC_2_VALID_4_5_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG <= 'x;
		local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_indvars_iv_push7_indvars_iv_next_output_regs_ready)
		begin
			local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG <= local_bb4_indvars_iv_push7_indvars_iv_next_result;
			local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_indvars_iv_push7_indvars_iv_next_stall_in))
			begin
				local_bb4_indvars_iv_push7_indvars_iv_next_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_5to6_bb4_notexit_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to6_bb4_notexit_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to6_bb4_notexit_0_NO_SHIFT_REG;
 logic rnode_5to6_bb4_notexit_0_reg_6_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to6_bb4_notexit_0_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_notexit_0_valid_out_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_notexit_0_stall_in_reg_6_NO_SHIFT_REG;
 logic rnode_5to6_bb4_notexit_0_stall_out_reg_6_NO_SHIFT_REG;

acl_data_fifo rnode_5to6_bb4_notexit_0_reg_6_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to6_bb4_notexit_0_reg_6_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to6_bb4_notexit_0_stall_in_reg_6_NO_SHIFT_REG),
	.valid_out(rnode_5to6_bb4_notexit_0_valid_out_reg_6_NO_SHIFT_REG),
	.stall_out(rnode_5to6_bb4_notexit_0_stall_out_reg_6_NO_SHIFT_REG),
	.data_in(local_bb4_notexit),
	.data_out(rnode_5to6_bb4_notexit_0_reg_6_NO_SHIFT_REG)
);

defparam rnode_5to6_bb4_notexit_0_reg_6_fifo.DEPTH = 1;
defparam rnode_5to6_bb4_notexit_0_reg_6_fifo.DATA_WIDTH = 1;
defparam rnode_5to6_bb4_notexit_0_reg_6_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_5to6_bb4_notexit_0_reg_6_fifo.IMPL = "shift_reg";

assign rnode_5to6_bb4_notexit_0_reg_6_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexit_stall_in_1 = 1'b0;
assign rnode_5to6_bb4_notexit_0_NO_SHIFT_REG = rnode_5to6_bb4_notexit_0_reg_6_NO_SHIFT_REG;
assign rnode_5to6_bb4_notexit_0_stall_in_reg_6_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_notexit_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot8_i419_stall_local;
wire local_bb4_lnot8_i419;

assign local_bb4_lnot8_i419 = ((local_bb4_and3_i413 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_i421_stall_local;
wire local_bb4_cmp11_i421;

assign local_bb4_cmp11_i421 = ((local_bb4_and3_i413 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u24_stall_local;
wire [31:0] local_bb4_var__u24;

assign local_bb4_var__u24 = ((local_bb4_and3_i413 & 32'hFF) | (local_bb4_and6_i417 & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i455_stall_local;
wire [31:0] local_bb4_add_i455;

assign local_bb4_add_i455 = ((local_bb4_and3_i413 & 32'hFF) + (local_bb4_and_i411 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_not_i427_stall_local;
wire local_bb4_lnot17_not_i427;

assign local_bb4_lnot17_not_i427 = (local_bb4_lnot17_i423 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u25_stall_local;
wire local_bb4_var__u25;

assign local_bb4_var__u25 = ((local_bb4_var__u23 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_conv1_i_i447_stall_local;
wire [63:0] local_bb4_conv1_i_i447;

assign local_bb4_conv1_i_i447[63:32] = 32'h0;
assign local_bb4_conv1_i_i447[31:0] = ((local_bb4_or47_i445 & 32'hFFFFFF) | 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(local_bb4_sub24_add2318_pop10_c0_ene2),
	.data_out(rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_sub24_add2318_pop10_c0_ene2_stall_in_1 = 1'b0;
assign rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_NO_SHIFT_REG = rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_add31_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add31_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_add31_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add31_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_add31_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add31_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add31_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_add31_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_add31_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_add31_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_add31_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_add31_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_add31_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(local_bb4_add31),
	.data_out(rnode_9to10_bb4_add31_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_add31_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_add31_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_add31_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_add31_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_add31_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add31_stall_in = 1'b0;
assign rnode_9to10_bb4_add31_0_NO_SHIFT_REG = rnode_9to10_bb4_add31_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_add31_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_add31_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_6to10_bb4_var__u22_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to10_bb4_var__u22_0_stall_in_NO_SHIFT_REG;
 logic rnode_6to10_bb4_var__u22_0_NO_SHIFT_REG;
 logic rnode_6to10_bb4_var__u22_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to10_bb4_var__u22_0_reg_10_NO_SHIFT_REG;
 logic rnode_6to10_bb4_var__u22_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_6to10_bb4_var__u22_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_6to10_bb4_var__u22_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_6to10_bb4_var__u22_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to10_bb4_var__u22_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to10_bb4_var__u22_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_6to10_bb4_var__u22_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_6to10_bb4_var__u22_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_5to6_bb4_var__u22_0_NO_SHIFT_REG),
	.data_out(rnode_6to10_bb4_var__u22_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_6to10_bb4_var__u22_0_reg_10_fifo.DEPTH = 4;
defparam rnode_6to10_bb4_var__u22_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_6to10_bb4_var__u22_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to10_bb4_var__u22_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_6to10_bb4_var__u22_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_5to6_bb4_var__u22_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_6to10_bb4_var__u22_0_NO_SHIFT_REG = rnode_6to10_bb4_var__u22_0_reg_10_NO_SHIFT_REG;
assign rnode_6to10_bb4_var__u22_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_6to10_bb4_var__u22_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb4_indvars_iv_push7_indvars_iv_next_NO_SHIFT_REG),
	.data_out(rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_fifo.DATA_WIDTH = 64;
defparam rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_indvars_iv_push7_indvars_iv_next_stall_in = 1'b0;
assign rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG = rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_6to8_bb4_notexit_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to8_bb4_notexit_0_stall_in_NO_SHIFT_REG;
 logic rnode_6to8_bb4_notexit_0_NO_SHIFT_REG;
 logic rnode_6to8_bb4_notexit_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to8_bb4_notexit_0_reg_8_NO_SHIFT_REG;
 logic rnode_6to8_bb4_notexit_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_6to8_bb4_notexit_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_6to8_bb4_notexit_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_6to8_bb4_notexit_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to8_bb4_notexit_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to8_bb4_notexit_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_6to8_bb4_notexit_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_6to8_bb4_notexit_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(rnode_5to6_bb4_notexit_0_NO_SHIFT_REG),
	.data_out(rnode_6to8_bb4_notexit_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_6to8_bb4_notexit_0_reg_8_fifo.DEPTH = 2;
defparam rnode_6to8_bb4_notexit_0_reg_8_fifo.DATA_WIDTH = 1;
defparam rnode_6to8_bb4_notexit_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to8_bb4_notexit_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_6to8_bb4_notexit_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_5to6_bb4_notexit_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_6to8_bb4_notexit_0_NO_SHIFT_REG = rnode_6to8_bb4_notexit_0_reg_8_NO_SHIFT_REG;
assign rnode_6to8_bb4_notexit_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_6to8_bb4_notexit_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i473_stall_local;
wire local_bb4_reduction_0_i473;

assign local_bb4_reduction_0_i473 = (local_bb4_lnot_i418 | local_bb4_lnot8_i419);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge8_demorgan_i424_stall_local;
wire local_bb4_brmerge8_demorgan_i424;

assign local_bb4_brmerge8_demorgan_i424 = (local_bb4_cmp11_i421 & local_bb4_lnot17_i423);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_not_i428_stall_local;
wire local_bb4_cmp11_not_i428;

assign local_bb4_cmp11_not_i428 = (local_bb4_cmp11_i421 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u26_stall_local;
wire local_bb4_var__u26;

assign local_bb4_var__u26 = (local_bb4_cmp_i420 | local_bb4_cmp11_i421);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u27_stall_local;
wire local_bb4_var__u27;

assign local_bb4_var__u27 = ((local_bb4_var__u24 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_idxprom32_stall_local;
wire [63:0] local_bb4_idxprom32;

assign local_bb4_idxprom32[63:32] = 32'h0;
assign local_bb4_idxprom32[31:0] = rnode_9to10_bb4_add31_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_var__u22_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_var__u22_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_var__u22_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_var__u22_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_var__u22_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_var__u22_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_var__u22_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_var__u22_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_var__u22_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_var__u22_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_var__u22_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_var__u22_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_var__u22_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(rnode_6to10_bb4_var__u22_0_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_var__u22_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_var__u22_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_var__u22_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_var__u22_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_var__u22_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_var__u22_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to10_bb4_var__u22_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_var__u22_0_NO_SHIFT_REG = rnode_10to11_bb4_var__u22_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_var__u22_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_var__u22_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG;
 logic rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG),
	.data_out(rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_fifo.DEPTH = 3;
defparam rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_fifo.DATA_WIDTH = 64;
defparam rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG = rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_reg_10_NO_SHIFT_REG;
assign rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_notexit_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_notexit_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to9_bb4_notexit_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_notexit_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_notexit_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_notexit_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_notexit_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_notexit_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_notexit_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_notexit_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_notexit_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_notexit_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_notexit_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_6to8_bb4_notexit_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_notexit_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_notexit_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_notexit_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_notexit_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_notexit_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_notexit_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to8_bb4_notexit_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_notexit_0_NO_SHIFT_REG = rnode_8to9_bb4_notexit_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_notexit_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_notexit_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge10_demorgan_i425_stall_local;
wire local_bb4_brmerge10_demorgan_i425;

assign local_bb4_brmerge10_demorgan_i425 = (local_bb4_brmerge8_demorgan_i424 & local_bb4_lnot_i418);

// This section implements an unregistered operation.
// 
wire local_bb4__mux9_mux_i426_stall_local;
wire local_bb4__mux9_mux_i426;

assign local_bb4__mux9_mux_i426 = (local_bb4_brmerge8_demorgan_i424 ^ local_bb4_cmp11_i421);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge3_i429_stall_local;
wire local_bb4_brmerge3_i429;

assign local_bb4_brmerge3_i429 = (local_bb4_var__u27 | local_bb4_cmp11_not_i428);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_i431_stall_local;
wire local_bb4__mux_mux_i431;

assign local_bb4__mux_mux_i431 = (local_bb4_var__u27 | local_bb4_cmp11_i421);

// This section implements an unregistered operation.
// 
wire local_bb4__not_i433_stall_local;
wire local_bb4__not_i433;

assign local_bb4__not_i433 = (local_bb4_var__u27 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_arrayidx33_valid_out;
wire local_bb4_arrayidx33_stall_in;
wire local_bb4_arrayidx33_inputs_ready;
wire local_bb4_arrayidx33_stall_local;
wire [63:0] local_bb4_arrayidx33;

assign local_bb4_arrayidx33_inputs_ready = rnode_9to10_bb4_add31_0_valid_out_NO_SHIFT_REG;
assign local_bb4_arrayidx33 = ((input_in & 64'hFFFFFFFFFFFFFC00) + ((local_bb4_idxprom32 & 64'hFFFFFFFF) << 6'h2));
assign local_bb4_arrayidx33_valid_out = 1'b1;
assign rnode_9to10_bb4_add31_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to10_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_NO_SHIFT_REG = rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_notexitcond_notexit_inputs_ready;
 reg local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_0;
 reg local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_1;
 reg local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_2;
 reg local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_3;
 reg local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_stall_in_4;
wire local_bb4_notexitcond_notexit_output_regs_ready;
wire local_bb4_notexitcond_notexit_result;
wire local_bb4_notexitcond_notexit_fu_valid_out;
wire local_bb4_notexitcond_notexit_fu_stall_out;
 reg local_bb4_notexitcond_notexit_NO_SHIFT_REG;
wire local_bb4_notexitcond_notexit_causedstall;

acl_push local_bb4_notexitcond_notexit_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(1'b1),
	.predicate(1'b0),
	.data_in(rnode_8to9_bb4_notexit_0_NO_SHIFT_REG),
	.stall_out(local_bb4_notexitcond_notexit_fu_stall_out),
	.valid_in(SFC_2_VALID_8_9_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond_notexit_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond_notexit_result),
	.feedback_out(feedback_data_out_1),
	.feedback_valid_out(feedback_valid_out_1),
	.feedback_stall_in(feedback_stall_in_1)
);

defparam local_bb4_notexitcond_notexit_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond_notexit_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond_notexit_feedback.FIFO_DEPTH = 8;
defparam local_bb4_notexitcond_notexit_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_notexitcond_notexit_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond_notexit_inputs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_output_regs_ready = 1'b1;
assign SFC_2_VALID_8_9_0_stall_in_3 = 1'b0;
assign rnode_8to9_bb4_notexit_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_notexitcond_notexit_causedstall = (SFC_2_VALID_8_9_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond_notexit_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond_notexit_output_regs_ready)
		begin
			local_bb4_notexitcond_notexit_NO_SHIFT_REG <= local_bb4_notexitcond_notexit_result;
			local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond_notexit_stall_in_0))
			begin
				local_bb4_notexitcond_notexit_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_1))
			begin
				local_bb4_notexitcond_notexit_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_2))
			begin
				local_bb4_notexitcond_notexit_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_3))
			begin
				local_bb4_notexitcond_notexit_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_notexitcond_notexit_stall_in_4))
			begin
				local_bb4_notexitcond_notexit_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__26_demorgan_i439_stall_local;
wire local_bb4__26_demorgan_i439;

assign local_bb4__26_demorgan_i439 = (local_bb4_cmp_i420 | local_bb4_brmerge10_demorgan_i425);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge5_i430_stall_local;
wire local_bb4_brmerge5_i430;

assign local_bb4_brmerge5_i430 = (local_bb4_brmerge3_i429 | local_bb4_lnot17_not_i427);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i434_stall_local;
wire local_bb4_reduction_3_i434;

assign local_bb4_reduction_3_i434 = (local_bb4_cmp11_i421 & local_bb4__not_i433);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_arrayidx33_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx33_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx33_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx33_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_10to11_bb4_arrayidx33_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx33_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx33_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_arrayidx33_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_arrayidx33_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_arrayidx33_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_arrayidx33_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_arrayidx33_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_arrayidx33_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in((local_bb4_arrayidx33 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_10to11_bb4_arrayidx33_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_arrayidx33_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_arrayidx33_0_reg_11_fifo.DATA_WIDTH = 64;
defparam rnode_10to11_bb4_arrayidx33_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_arrayidx33_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_arrayidx33_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_arrayidx33_stall_in = 1'b0;
assign rnode_10to11_bb4_arrayidx33_0_NO_SHIFT_REG = rnode_10to11_bb4_arrayidx33_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_arrayidx33_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx33_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_sub24_add2318_push10_sub24_add2318_pop10_inputs_ready;
 reg local_bb4_sub24_add2318_push10_sub24_add2318_pop10_valid_out_NO_SHIFT_REG;
wire local_bb4_sub24_add2318_push10_sub24_add2318_pop10_stall_in;
wire local_bb4_sub24_add2318_push10_sub24_add2318_pop10_output_regs_ready;
wire [31:0] local_bb4_sub24_add2318_push10_sub24_add2318_pop10_result;
wire local_bb4_sub24_add2318_push10_sub24_add2318_pop10_fu_valid_out;
wire local_bb4_sub24_add2318_push10_sub24_add2318_pop10_fu_stall_out;
 reg [31:0] local_bb4_sub24_add2318_push10_sub24_add2318_pop10_NO_SHIFT_REG;
wire local_bb4_sub24_add2318_push10_sub24_add2318_pop10_causedstall;

acl_push local_bb4_sub24_add2318_push10_sub24_add2318_pop10_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_NO_SHIFT_REG),
	.stall_out(local_bb4_sub24_add2318_push10_sub24_add2318_pop10_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sub24_add2318_push10_sub24_add2318_pop10_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_sub24_add2318_push10_sub24_add2318_pop10_result),
	.feedback_out(feedback_data_out_10),
	.feedback_valid_out(feedback_valid_out_10),
	.feedback_stall_in(feedback_stall_in_10)
);

defparam local_bb4_sub24_add2318_push10_sub24_add2318_pop10_feedback.STALLFREE = 1;
defparam local_bb4_sub24_add2318_push10_sub24_add2318_pop10_feedback.DATA_WIDTH = 32;
defparam local_bb4_sub24_add2318_push10_sub24_add2318_pop10_feedback.FIFO_DEPTH = 9;
defparam local_bb4_sub24_add2318_push10_sub24_add2318_pop10_feedback.MIN_FIFO_LATENCY = 8;
defparam local_bb4_sub24_add2318_push10_sub24_add2318_pop10_feedback.STYLE = "REGULAR";

assign local_bb4_sub24_add2318_push10_sub24_add2318_pop10_inputs_ready = 1'b1;
assign local_bb4_sub24_add2318_push10_sub24_add2318_pop10_output_regs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_1 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_4 = 1'b0;
assign rnode_9to10_bb4_sub24_add2318_pop10_c0_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_sub24_add2318_push10_sub24_add2318_pop10_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_sub24_add2318_push10_sub24_add2318_pop10_NO_SHIFT_REG <= 'x;
		local_bb4_sub24_add2318_push10_sub24_add2318_pop10_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_sub24_add2318_push10_sub24_add2318_pop10_output_regs_ready)
		begin
			local_bb4_sub24_add2318_push10_sub24_add2318_pop10_NO_SHIFT_REG <= local_bb4_sub24_add2318_push10_sub24_add2318_pop10_result;
			local_bb4_sub24_add2318_push10_sub24_add2318_pop10_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_sub24_add2318_push10_sub24_add2318_pop10_stall_in))
			begin
				local_bb4_sub24_add2318_push10_sub24_add2318_pop10_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4__push12__pop12_inputs_ready;
 reg local_bb4__push12__pop12_valid_out_NO_SHIFT_REG;
wire local_bb4__push12__pop12_stall_in;
wire local_bb4__push12__pop12_output_regs_ready;
wire local_bb4__push12__pop12_result;
wire local_bb4__push12__pop12_fu_valid_out;
wire local_bb4__push12__pop12_fu_stall_out;
 reg local_bb4__push12__pop12_NO_SHIFT_REG;
wire local_bb4__push12__pop12_causedstall;

acl_push local_bb4__push12__pop12_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4__pop12_c0_ene4),
	.stall_out(local_bb4__push12__pop12_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4__push12__pop12_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4__push12__pop12_result),
	.feedback_out(feedback_data_out_12),
	.feedback_valid_out(feedback_valid_out_12),
	.feedback_stall_in(feedback_stall_in_12)
);

defparam local_bb4__push12__pop12_feedback.STALLFREE = 1;
defparam local_bb4__push12__pop12_feedback.DATA_WIDTH = 1;
defparam local_bb4__push12__pop12_feedback.FIFO_DEPTH = 9;
defparam local_bb4__push12__pop12_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4__push12__pop12_feedback.STYLE = "REGULAR";

assign local_bb4__push12__pop12_inputs_ready = 1'b1;
assign local_bb4__push12__pop12_output_regs_ready = 1'b1;
assign local_bb4__pop12_c0_ene4_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_2 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_5 = 1'b0;
assign local_bb4__push12__pop12_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4__push12__pop12_NO_SHIFT_REG <= 'x;
		local_bb4__push12__pop12_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4__push12__pop12_output_regs_ready)
		begin
			local_bb4__push12__pop12_NO_SHIFT_REG <= local_bb4__push12__pop12_result;
			local_bb4__push12__pop12_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4__push12__pop12_stall_in))
			begin
				local_bb4__push12__pop12_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_notexitcond1520_push13_notexitcond1520_pop13_inputs_ready;
 reg local_bb4_notexitcond1520_push13_notexitcond1520_pop13_valid_out_NO_SHIFT_REG;
wire local_bb4_notexitcond1520_push13_notexitcond1520_pop13_stall_in;
wire local_bb4_notexitcond1520_push13_notexitcond1520_pop13_output_regs_ready;
wire local_bb4_notexitcond1520_push13_notexitcond1520_pop13_result;
wire local_bb4_notexitcond1520_push13_notexitcond1520_pop13_fu_valid_out;
wire local_bb4_notexitcond1520_push13_notexitcond1520_pop13_fu_stall_out;
 reg local_bb4_notexitcond1520_push13_notexitcond1520_pop13_NO_SHIFT_REG;
wire local_bb4_notexitcond1520_push13_notexitcond1520_pop13_causedstall;

acl_push local_bb4_notexitcond1520_push13_notexitcond1520_pop13_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb4_notexitcond1520_pop13_c0_ene5),
	.stall_out(local_bb4_notexitcond1520_push13_notexitcond1520_pop13_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_notexitcond1520_push13_notexitcond1520_pop13_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_notexitcond1520_push13_notexitcond1520_pop13_result),
	.feedback_out(feedback_data_out_13),
	.feedback_valid_out(feedback_valid_out_13),
	.feedback_stall_in(feedback_stall_in_13)
);

defparam local_bb4_notexitcond1520_push13_notexitcond1520_pop13_feedback.STALLFREE = 1;
defparam local_bb4_notexitcond1520_push13_notexitcond1520_pop13_feedback.DATA_WIDTH = 1;
defparam local_bb4_notexitcond1520_push13_notexitcond1520_pop13_feedback.FIFO_DEPTH = 9;
defparam local_bb4_notexitcond1520_push13_notexitcond1520_pop13_feedback.MIN_FIFO_LATENCY = 9;
defparam local_bb4_notexitcond1520_push13_notexitcond1520_pop13_feedback.STYLE = "REGULAR";

assign local_bb4_notexitcond1520_push13_notexitcond1520_pop13_inputs_ready = 1'b1;
assign local_bb4_notexitcond1520_push13_notexitcond1520_pop13_output_regs_ready = 1'b1;
assign local_bb4_notexitcond1520_pop13_c0_ene5_stall_in_0 = 1'b0;
assign local_bb4_notexitcond_notexit_stall_in_3 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_6 = 1'b0;
assign local_bb4_notexitcond1520_push13_notexitcond1520_pop13_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_notexitcond1520_push13_notexitcond1520_pop13_NO_SHIFT_REG <= 'x;
		local_bb4_notexitcond1520_push13_notexitcond1520_pop13_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_notexitcond1520_push13_notexitcond1520_pop13_output_regs_ready)
		begin
			local_bb4_notexitcond1520_push13_notexitcond1520_pop13_NO_SHIFT_REG <= local_bb4_notexitcond1520_push13_notexitcond1520_pop13_result;
			local_bb4_notexitcond1520_push13_notexitcond1520_pop13_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_notexitcond1520_push13_notexitcond1520_pop13_stall_in))
			begin
				local_bb4_notexitcond1520_push13_notexitcond1520_pop13_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_notexitcond_notexit_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_notexitcond_notexit_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_notexitcond_notexit_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_notexitcond_notexit_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_notexitcond_notexit_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_4 = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG = rnode_10to11_bb4_notexitcond_notexit_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_notexitcond_notexit_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_mux_i432_stall_local;
wire local_bb4__mux_mux_mux_i432;

assign local_bb4__mux_mux_mux_i432 = (local_bb4_brmerge5_i430 & local_bb4__mux_mux_i431);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i435_stall_local;
wire local_bb4_reduction_5_i435;

assign local_bb4_reduction_5_i435 = (local_bb4_lnot14_i422 & local_bb4_reduction_3_i434);

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi124_stall_local;
wire [191:0] local_bb4_c0_exi124;

assign local_bb4_c0_exi124[63:0] = 64'bx;
assign local_bb4_c0_exi124[127:64] = (rnode_10to11_bb4_arrayidx33_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
assign local_bb4_c0_exi124[191:128] = 64'bx;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i436_stall_local;
wire local_bb4_reduction_6_i436;

assign local_bb4_reduction_6_i436 = (local_bb4_var__u25 & local_bb4_reduction_5_i435);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i437_stall_local;
wire local_bb4__24_i437;

assign local_bb4__24_i437 = (local_bb4_cmp_i420 ? local_bb4_reduction_6_i436 : local_bb4_brmerge10_demorgan_i425);

// This section implements an unregistered operation.
// 
wire local_bb4__25_i438_stall_local;
wire local_bb4__25_i438;

assign local_bb4__25_i438 = (local_bb4__24_i437 ? local_bb4_lnot14_i422 : local_bb4__mux_mux_mux_i432);

// This section implements an unregistered operation.
// 
wire local_bb4_gaussian_ROM4119_pop11_c0_ene3_valid_out_1;
wire local_bb4_gaussian_ROM4119_pop11_c0_ene3_stall_in_1;
wire local_bb4_xor_i414_valid_out;
wire local_bb4_xor_i414_stall_in;
wire local_bb4_add_i455_valid_out;
wire local_bb4_add_i455_stall_in;
wire local_bb4_conv_i_i446_valid_out;
wire local_bb4_conv_i_i446_stall_in;
wire local_bb4_reduction_0_i473_valid_out;
wire local_bb4_reduction_0_i473_stall_in;
wire local_bb4__28_i442_valid_out;
wire local_bb4__28_i442_stall_in;
wire local_bb4_var__u26_valid_out;
wire local_bb4_var__u26_stall_in;
wire local_bb4__27_i440_valid_out;
wire local_bb4__27_i440_stall_in;
wire local_bb4_conv1_i_i447_valid_out;
wire local_bb4_conv1_i_i447_stall_in;
wire local_bb4__27_i440_inputs_ready;
wire local_bb4__27_i440_stall_local;
wire local_bb4__27_i440;

assign local_bb4__27_i440_inputs_ready = (SFC_2_VALID_5_6_0_valid_out_1_NO_SHIFT_REG & rnode_5to6_bb4_c0_ene123_0_valid_out_0_NO_SHIFT_REG & rnode_5to6_bb4_c0_ene3_0_valid_out_NO_SHIFT_REG & local_bb4_gaussian_ROM_arrayidx44_valid_out_NO_SHIFT_REG);
assign local_bb4__27_i440 = (local_bb4__26_demorgan_i439 ? local_bb4__25_i438 : local_bb4__mux9_mux_i426);
assign local_bb4_gaussian_ROM4119_pop11_c0_ene3_valid_out_1 = 1'b1;
assign local_bb4_xor_i414_valid_out = 1'b1;
assign local_bb4_add_i455_valid_out = 1'b1;
assign local_bb4_conv_i_i446_valid_out = 1'b1;
assign local_bb4_reduction_0_i473_valid_out = 1'b1;
assign local_bb4__28_i442_valid_out = 1'b1;
assign local_bb4_var__u26_valid_out = 1'b1;
assign local_bb4__27_i440_valid_out = 1'b1;
assign local_bb4_conv1_i_i447_valid_out = 1'b1;
assign SFC_2_VALID_5_6_0_stall_in_1 = 1'b0;
assign rnode_5to6_bb4_c0_ene123_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_5to6_bb4_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_gaussian_ROM_arrayidx44_stall_in = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb4_gaussian_ROM4119_pop11_c0_ene3),
	.data_out(rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_fifo.DATA_WIDTH = 32;
defparam rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_gaussian_ROM4119_pop11_c0_ene3_stall_in_1 = 1'b0;
assign rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG = rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_xor_i414_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_xor_i414_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_xor_i414_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_xor_i414_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_xor_i414_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_xor_i414_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_xor_i414_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_xor_i414_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_xor_i414_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_xor_i414_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_xor_i414_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_xor_i414_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_xor_i414_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i414),
	.data_out(rnode_6to7_bb4_xor_i414_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_xor_i414_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_xor_i414_0_reg_7_fifo.DATA_WIDTH = 32;
defparam rnode_6to7_bb4_xor_i414_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_xor_i414_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_xor_i414_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i414_stall_in = 1'b0;
assign rnode_6to7_bb4_xor_i414_0_NO_SHIFT_REG = rnode_6to7_bb4_xor_i414_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_xor_i414_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_xor_i414_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_add_i455_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_add_i455_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_add_i455_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_add_i455_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_6to7_bb4_add_i455_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_add_i455_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_add_i455_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_add_i455_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_add_i455_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_add_i455_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_add_i455_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_add_i455_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_add_i455_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in((local_bb4_add_i455 & 32'h1FF)),
	.data_out(rnode_6to7_bb4_add_i455_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_add_i455_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_add_i455_0_reg_7_fifo.DATA_WIDTH = 32;
defparam rnode_6to7_bb4_add_i455_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_add_i455_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_add_i455_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add_i455_stall_in = 1'b0;
assign rnode_6to7_bb4_add_i455_0_NO_SHIFT_REG = rnode_6to7_bb4_add_i455_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_add_i455_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_add_i455_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_reduction_0_i473_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_reduction_0_i473_0_stall_in_NO_SHIFT_REG;
 logic rnode_6to7_bb4_reduction_0_i473_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_reduction_0_i473_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to7_bb4_reduction_0_i473_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_reduction_0_i473_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_reduction_0_i473_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_reduction_0_i473_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_reduction_0_i473_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_reduction_0_i473_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_reduction_0_i473_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_reduction_0_i473_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_reduction_0_i473_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_0_i473),
	.data_out(rnode_6to7_bb4_reduction_0_i473_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_reduction_0_i473_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_reduction_0_i473_0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_6to7_bb4_reduction_0_i473_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_reduction_0_i473_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_reduction_0_i473_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_0_i473_stall_in = 1'b0;
assign rnode_6to7_bb4_reduction_0_i473_0_NO_SHIFT_REG = rnode_6to7_bb4_reduction_0_i473_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_reduction_0_i473_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_reduction_0_i473_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4__28_i442_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4__28_i442_0_stall_in_NO_SHIFT_REG;
 logic rnode_6to7_bb4__28_i442_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4__28_i442_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to7_bb4__28_i442_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4__28_i442_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4__28_i442_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4__28_i442_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4__28_i442_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4__28_i442_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4__28_i442_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4__28_i442_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4__28_i442_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb4__28_i442),
	.data_out(rnode_6to7_bb4__28_i442_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4__28_i442_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4__28_i442_0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_6to7_bb4__28_i442_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4__28_i442_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4__28_i442_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__28_i442_stall_in = 1'b0;
assign rnode_6to7_bb4__28_i442_0_NO_SHIFT_REG = rnode_6to7_bb4__28_i442_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4__28_i442_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4__28_i442_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4_var__u26_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4_var__u26_0_stall_in_NO_SHIFT_REG;
 logic rnode_6to7_bb4_var__u26_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4_var__u26_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to7_bb4_var__u26_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_var__u26_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_var__u26_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4_var__u26_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4_var__u26_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4_var__u26_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4_var__u26_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4_var__u26_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4_var__u26_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb4_var__u26),
	.data_out(rnode_6to7_bb4_var__u26_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4_var__u26_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4_var__u26_0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_6to7_bb4_var__u26_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4_var__u26_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4_var__u26_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u26_stall_in = 1'b0;
assign rnode_6to7_bb4_var__u26_0_NO_SHIFT_REG = rnode_6to7_bb4_var__u26_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4_var__u26_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4_var__u26_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_6to7_bb4__27_i440_0_valid_out_NO_SHIFT_REG;
 logic rnode_6to7_bb4__27_i440_0_stall_in_NO_SHIFT_REG;
 logic rnode_6to7_bb4__27_i440_0_NO_SHIFT_REG;
 logic rnode_6to7_bb4__27_i440_0_reg_7_inputs_ready_NO_SHIFT_REG;
 logic rnode_6to7_bb4__27_i440_0_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4__27_i440_0_valid_out_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4__27_i440_0_stall_in_reg_7_NO_SHIFT_REG;
 logic rnode_6to7_bb4__27_i440_0_stall_out_reg_7_NO_SHIFT_REG;

acl_data_fifo rnode_6to7_bb4__27_i440_0_reg_7_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_6to7_bb4__27_i440_0_reg_7_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_6to7_bb4__27_i440_0_stall_in_reg_7_NO_SHIFT_REG),
	.valid_out(rnode_6to7_bb4__27_i440_0_valid_out_reg_7_NO_SHIFT_REG),
	.stall_out(rnode_6to7_bb4__27_i440_0_stall_out_reg_7_NO_SHIFT_REG),
	.data_in(local_bb4__27_i440),
	.data_out(rnode_6to7_bb4__27_i440_0_reg_7_NO_SHIFT_REG)
);

defparam rnode_6to7_bb4__27_i440_0_reg_7_fifo.DEPTH = 1;
defparam rnode_6to7_bb4__27_i440_0_reg_7_fifo.DATA_WIDTH = 1;
defparam rnode_6to7_bb4__27_i440_0_reg_7_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_6to7_bb4__27_i440_0_reg_7_fifo.IMPL = "shift_reg";

assign rnode_6to7_bb4__27_i440_0_reg_7_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__27_i440_stall_in = 1'b0;
assign rnode_6to7_bb4__27_i440_0_NO_SHIFT_REG = rnode_6to7_bb4__27_i440_0_reg_7_NO_SHIFT_REG;
assign rnode_6to7_bb4__27_i440_0_stall_in_reg_7_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4__27_i440_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_mul_i_i448_inputs_ready;
 reg local_bb4_mul_i_i448_valid_out_0_NO_SHIFT_REG;
wire local_bb4_mul_i_i448_stall_in_0;
 reg local_bb4_mul_i_i448_valid_out_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i448_stall_in_1;
wire local_bb4_mul_i_i448_output_regs_ready;
wire [63:0] local_bb4_mul_i_i448;
 reg local_bb4_mul_i_i448_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul_i_i448_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i448_causedstall;

acl_int_mult int_module_local_bb4_mul_i_i448 (
	.clock(clock),
	.dataa(((local_bb4_conv1_i_i447 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb4_conv_i_i446 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb4_mul_i_i448_output_regs_ready),
	.result(local_bb4_mul_i_i448)
);

defparam int_module_local_bb4_mul_i_i448.INPUT1_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i448.INPUT2_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i448.OUTPUT_WIDTH = 64;
defparam int_module_local_bb4_mul_i_i448.LATENCY = 3;
defparam int_module_local_bb4_mul_i_i448.SIGNED = 0;

assign local_bb4_mul_i_i448_inputs_ready = 1'b1;
assign local_bb4_mul_i_i448_output_regs_ready = 1'b1;
assign local_bb4_conv1_i_i447_stall_in = 1'b0;
assign local_bb4_conv_i_i446_stall_in = 1'b0;
assign local_bb4_mul_i_i448_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i448_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i448_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i448_output_regs_ready)
		begin
			local_bb4_mul_i_i448_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i448_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul_i_i448_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i448_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i448_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i448_output_regs_ready)
		begin
			local_bb4_mul_i_i448_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i448_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul_i_i448_stall_in_0))
			begin
				local_bb4_mul_i_i448_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_mul_i_i448_stall_in_1))
			begin
				local_bb4_mul_i_i448_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_fifo.DEPTH = 2;
defparam rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG = rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_9_NO_SHIFT_REG;
assign rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_7to10_bb4_xor_i414_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to10_bb4_xor_i414_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_7to10_bb4_xor_i414_0_NO_SHIFT_REG;
 logic rnode_7to10_bb4_xor_i414_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to10_bb4_xor_i414_0_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_xor_i414_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_xor_i414_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_xor_i414_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_7to10_bb4_xor_i414_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to10_bb4_xor_i414_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to10_bb4_xor_i414_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_7to10_bb4_xor_i414_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_7to10_bb4_xor_i414_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_xor_i414_0_NO_SHIFT_REG),
	.data_out(rnode_7to10_bb4_xor_i414_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_7to10_bb4_xor_i414_0_reg_10_fifo.DEPTH = 3;
defparam rnode_7to10_bb4_xor_i414_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_7to10_bb4_xor_i414_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to10_bb4_xor_i414_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_7to10_bb4_xor_i414_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_xor_i414_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_7to10_bb4_xor_i414_0_NO_SHIFT_REG = rnode_7to10_bb4_xor_i414_0_reg_10_NO_SHIFT_REG;
assign rnode_7to10_bb4_xor_i414_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_7to10_bb4_xor_i414_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_add_i455_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add_i455_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add_i455_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add_i455_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_7to8_bb4_add_i455_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add_i455_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add_i455_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_add_i455_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_add_i455_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_add_i455_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_add_i455_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_add_i455_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_add_i455_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in((rnode_6to7_bb4_add_i455_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_7to8_bb4_add_i455_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_add_i455_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_add_i455_0_reg_8_fifo.DATA_WIDTH = 32;
defparam rnode_7to8_bb4_add_i455_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_add_i455_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_add_i455_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_add_i455_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_add_i455_0_NO_SHIFT_REG = rnode_7to8_bb4_add_i455_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_add_i455_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_add_i455_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_7to10_bb4_reduction_0_i473_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to10_bb4_reduction_0_i473_0_stall_in_NO_SHIFT_REG;
 logic rnode_7to10_bb4_reduction_0_i473_0_NO_SHIFT_REG;
 logic rnode_7to10_bb4_reduction_0_i473_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_7to10_bb4_reduction_0_i473_0_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_reduction_0_i473_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_reduction_0_i473_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_7to10_bb4_reduction_0_i473_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_7to10_bb4_reduction_0_i473_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to10_bb4_reduction_0_i473_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to10_bb4_reduction_0_i473_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_7to10_bb4_reduction_0_i473_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_7to10_bb4_reduction_0_i473_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_reduction_0_i473_0_NO_SHIFT_REG),
	.data_out(rnode_7to10_bb4_reduction_0_i473_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_7to10_bb4_reduction_0_i473_0_reg_10_fifo.DEPTH = 3;
defparam rnode_7to10_bb4_reduction_0_i473_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_7to10_bb4_reduction_0_i473_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to10_bb4_reduction_0_i473_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_7to10_bb4_reduction_0_i473_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_reduction_0_i473_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_7to10_bb4_reduction_0_i473_0_NO_SHIFT_REG = rnode_7to10_bb4_reduction_0_i473_0_reg_10_NO_SHIFT_REG;
assign rnode_7to10_bb4_reduction_0_i473_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_7to10_bb4_reduction_0_i473_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4_var__u26_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u26_0_stall_in_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u26_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u26_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u26_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u26_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u26_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4_var__u26_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4_var__u26_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4_var__u26_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4_var__u26_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4_var__u26_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4_var__u26_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(rnode_6to7_bb4_var__u26_0_NO_SHIFT_REG),
	.data_out(rnode_7to8_bb4_var__u26_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4_var__u26_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4_var__u26_0_reg_8_fifo.DATA_WIDTH = 1;
defparam rnode_7to8_bb4_var__u26_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4_var__u26_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4_var__u26_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_6to7_bb4_var__u26_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_var__u26_0_NO_SHIFT_REG = rnode_7to8_bb4_var__u26_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4_var__u26_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4_var__u26_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i443_valid_out;
wire local_bb4__29_i443_stall_in;
wire local_bb4__29_i443_inputs_ready;
wire local_bb4__29_i443_stall_local;
wire local_bb4__29_i443;

assign local_bb4__29_i443_inputs_ready = (rnode_6to7_bb4__28_i442_0_valid_out_NO_SHIFT_REG & rnode_6to7_bb4__27_i440_0_valid_out_NO_SHIFT_REG);
assign local_bb4__29_i443 = (rnode_6to7_bb4__28_i442_0_NO_SHIFT_REG | rnode_6to7_bb4__27_i440_0_NO_SHIFT_REG);
assign local_bb4__29_i443_valid_out = 1'b1;
assign rnode_6to7_bb4__28_i442_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_6to7_bb4__27_i440_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_conv3_i_i449_stall_local;
wire [31:0] local_bb4_conv3_i_i449;
wire [63:0] local_bb4_conv3_i_i449$ps;

assign local_bb4_conv3_i_i449$ps = (local_bb4_mul_i_i448 & 64'hFFFFFFFFFFFF);
assign local_bb4_conv3_i_i449 = local_bb4_conv3_i_i449$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u28_stall_local;
wire [63:0] local_bb4_var__u28;

assign local_bb4_var__u28 = ((local_bb4_mul_i_i448 & 64'hFFFFFFFFFFFF) >> 64'h18);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to9_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG = rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_xor_i414_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_xor_i414_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_xor_i414_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_xor_i414_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_xor_i414_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_xor_i414_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_xor_i414_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_xor_i414_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_xor_i414_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_xor_i414_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_xor_i414_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_xor_i414_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_xor_i414_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(rnode_7to10_bb4_xor_i414_0_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_xor_i414_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_xor_i414_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_xor_i414_0_reg_11_fifo.DATA_WIDTH = 32;
defparam rnode_10to11_bb4_xor_i414_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_xor_i414_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_xor_i414_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to10_bb4_xor_i414_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_xor_i414_0_NO_SHIFT_REG = rnode_10to11_bb4_xor_i414_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_xor_i414_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_xor_i414_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_add_i455_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_add_i455_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_add_i455_1_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_add_i455_2_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_8to9_bb4_add_i455_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_valid_out_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_stall_in_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_add_i455_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_add_i455_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_add_i455_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_add_i455_0_stall_in_0_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_add_i455_0_valid_out_0_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_add_i455_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in((rnode_7to8_bb4_add_i455_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_8to9_bb4_add_i455_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_add_i455_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_add_i455_0_reg_9_fifo.DATA_WIDTH = 32;
defparam rnode_8to9_bb4_add_i455_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_add_i455_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_add_i455_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_add_i455_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_add_i455_0_stall_in_0_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_add_i455_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_add_i455_0_NO_SHIFT_REG = rnode_8to9_bb4_add_i455_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_add_i455_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_add_i455_1_NO_SHIFT_REG = rnode_8to9_bb4_add_i455_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_add_i455_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_8to9_bb4_add_i455_2_NO_SHIFT_REG = rnode_8to9_bb4_add_i455_0_reg_9_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_reduction_0_i473_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_reduction_0_i473_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4_reduction_0_i473_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_reduction_0_i473_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4_reduction_0_i473_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_reduction_0_i473_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_reduction_0_i473_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_reduction_0_i473_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_reduction_0_i473_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_reduction_0_i473_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_reduction_0_i473_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_reduction_0_i473_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_reduction_0_i473_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(rnode_7to10_bb4_reduction_0_i473_0_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4_reduction_0_i473_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_reduction_0_i473_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_reduction_0_i473_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4_reduction_0_i473_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_reduction_0_i473_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_reduction_0_i473_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to10_bb4_reduction_0_i473_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_reduction_0_i473_0_NO_SHIFT_REG = rnode_10to11_bb4_reduction_0_i473_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_reduction_0_i473_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_reduction_0_i473_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_8to9_bb4_var__u26_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to9_bb4_var__u26_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to9_bb4_var__u26_0_NO_SHIFT_REG;
 logic rnode_8to9_bb4_var__u26_0_reg_9_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to9_bb4_var__u26_0_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_var__u26_0_valid_out_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_var__u26_0_stall_in_reg_9_NO_SHIFT_REG;
 logic rnode_8to9_bb4_var__u26_0_stall_out_reg_9_NO_SHIFT_REG;

acl_data_fifo rnode_8to9_bb4_var__u26_0_reg_9_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to9_bb4_var__u26_0_reg_9_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to9_bb4_var__u26_0_stall_in_reg_9_NO_SHIFT_REG),
	.valid_out(rnode_8to9_bb4_var__u26_0_valid_out_reg_9_NO_SHIFT_REG),
	.stall_out(rnode_8to9_bb4_var__u26_0_stall_out_reg_9_NO_SHIFT_REG),
	.data_in(rnode_7to8_bb4_var__u26_0_NO_SHIFT_REG),
	.data_out(rnode_8to9_bb4_var__u26_0_reg_9_NO_SHIFT_REG)
);

defparam rnode_8to9_bb4_var__u26_0_reg_9_fifo.DEPTH = 1;
defparam rnode_8to9_bb4_var__u26_0_reg_9_fifo.DATA_WIDTH = 1;
defparam rnode_8to9_bb4_var__u26_0_reg_9_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to9_bb4_var__u26_0_reg_9_fifo.IMPL = "shift_reg";

assign rnode_8to9_bb4_var__u26_0_reg_9_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4_var__u26_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_var__u26_0_NO_SHIFT_REG = rnode_8to9_bb4_var__u26_0_reg_9_NO_SHIFT_REG;
assign rnode_8to9_bb4_var__u26_0_stall_in_reg_9_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_var__u26_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_7to8_bb4__29_i443_0_valid_out_NO_SHIFT_REG;
 logic rnode_7to8_bb4__29_i443_0_stall_in_NO_SHIFT_REG;
 logic rnode_7to8_bb4__29_i443_0_NO_SHIFT_REG;
 logic rnode_7to8_bb4__29_i443_0_reg_8_inputs_ready_NO_SHIFT_REG;
 logic rnode_7to8_bb4__29_i443_0_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4__29_i443_0_valid_out_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4__29_i443_0_stall_in_reg_8_NO_SHIFT_REG;
 logic rnode_7to8_bb4__29_i443_0_stall_out_reg_8_NO_SHIFT_REG;

acl_data_fifo rnode_7to8_bb4__29_i443_0_reg_8_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_7to8_bb4__29_i443_0_reg_8_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_7to8_bb4__29_i443_0_stall_in_reg_8_NO_SHIFT_REG),
	.valid_out(rnode_7to8_bb4__29_i443_0_valid_out_reg_8_NO_SHIFT_REG),
	.stall_out(rnode_7to8_bb4__29_i443_0_stall_out_reg_8_NO_SHIFT_REG),
	.data_in(local_bb4__29_i443),
	.data_out(rnode_7to8_bb4__29_i443_0_reg_8_NO_SHIFT_REG)
);

defparam rnode_7to8_bb4__29_i443_0_reg_8_fifo.DEPTH = 1;
defparam rnode_7to8_bb4__29_i443_0_reg_8_fifo.DATA_WIDTH = 1;
defparam rnode_7to8_bb4__29_i443_0_reg_8_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_7to8_bb4__29_i443_0_reg_8_fifo.IMPL = "shift_reg";

assign rnode_7to8_bb4__29_i443_0_reg_8_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__29_i443_stall_in = 1'b0;
assign rnode_7to8_bb4__29_i443_0_NO_SHIFT_REG = rnode_7to8_bb4__29_i443_0_reg_8_NO_SHIFT_REG;
assign rnode_7to8_bb4__29_i443_0_stall_in_reg_8_NO_SHIFT_REG = 1'b0;
assign rnode_7to8_bb4__29_i443_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i16_i452_stall_local;
wire [31:0] local_bb4_shr_i16_i452;

assign local_bb4_shr_i16_i452 = (local_bb4_conv3_i_i449 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i18_i454_stall_local;
wire [31:0] local_bb4_shl1_i18_i454;

assign local_bb4_shl1_i18_i454 = (local_bb4_conv3_i_i449 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u29_stall_local;
wire [31:0] local_bb4_var__u29;

assign local_bb4_var__u29 = (local_bb4_conv3_i_i449 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i_i462_stall_local;
wire [31:0] local_bb4_shl1_i_i462;

assign local_bb4_shl1_i_i462 = (local_bb4_conv3_i_i449 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb4__tr_i450_stall_local;
wire [31:0] local_bb4__tr_i450;
wire [63:0] local_bb4__tr_i450$ps;

assign local_bb4__tr_i450$ps = (local_bb4_var__u28 & 64'hFFFFFF);
assign local_bb4__tr_i450 = local_bb4__tr_i450$ps[31:0];

// This section implements a registered operation.
// 
wire local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_inputs_ready;
 reg local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_valid_out_NO_SHIFT_REG;
wire local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_stall_in;
wire local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_output_regs_ready;
wire [31:0] local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_result;
wire local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_fu_valid_out;
wire local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_fu_stall_out;
 reg [31:0] local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_NO_SHIFT_REG;
wire local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_causedstall;

acl_push local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_bb4_notexitcond_notexit_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_NO_SHIFT_REG),
	.stall_out(local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_fu_stall_out),
	.valid_in(SFC_2_VALID_9_10_0_NO_SHIFT_REG),
	.valid_out(local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_result),
	.feedback_out(feedback_data_out_11),
	.feedback_valid_out(feedback_valid_out_11),
	.feedback_stall_in(feedback_stall_in_11)
);

defparam local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_feedback.STALLFREE = 1;
defparam local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_feedback.DATA_WIDTH = 32;
defparam local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_feedback.FIFO_DEPTH = 9;
defparam local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_feedback.MIN_FIFO_LATENCY = 5;
defparam local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_feedback.STYLE = "REGULAR";

assign local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_inputs_ready = 1'b1;
assign local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_output_regs_ready = 1'b1;
assign local_bb4_notexitcond_notexit_stall_in_0 = 1'b0;
assign SFC_2_VALID_9_10_0_stall_in_3 = 1'b0;
assign rnode_9to10_bb4_gaussian_ROM4119_pop11_c0_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_causedstall = (SFC_2_VALID_9_10_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_NO_SHIFT_REG <= 'x;
		local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_output_regs_ready)
		begin
			local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_NO_SHIFT_REG <= local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_result;
			local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_stall_in))
			begin
				local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and4_i415_stall_local;
wire [31:0] local_bb4_and4_i415;

assign local_bb4_and4_i415 = (rnode_10to11_bb4_xor_i414_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_inc_i458_stall_local;
wire [31:0] local_bb4_inc_i458;

assign local_bb4_inc_i458 = ((rnode_8to9_bb4_add_i455_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp50_not_i463_stall_local;
wire local_bb4_cmp50_not_i463;

assign local_bb4_cmp50_not_i463 = ((rnode_8to9_bb4_add_i455_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_8to10_bb4__29_i443_0_valid_out_NO_SHIFT_REG;
 logic rnode_8to10_bb4__29_i443_0_stall_in_NO_SHIFT_REG;
 logic rnode_8to10_bb4__29_i443_0_NO_SHIFT_REG;
 logic rnode_8to10_bb4__29_i443_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic rnode_8to10_bb4__29_i443_0_reg_10_NO_SHIFT_REG;
 logic rnode_8to10_bb4__29_i443_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_8to10_bb4__29_i443_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_8to10_bb4__29_i443_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_8to10_bb4__29_i443_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_8to10_bb4__29_i443_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_8to10_bb4__29_i443_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_8to10_bb4__29_i443_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_8to10_bb4__29_i443_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in(rnode_7to8_bb4__29_i443_0_NO_SHIFT_REG),
	.data_out(rnode_8to10_bb4__29_i443_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_8to10_bb4__29_i443_0_reg_10_fifo.DEPTH = 2;
defparam rnode_8to10_bb4__29_i443_0_reg_10_fifo.DATA_WIDTH = 1;
defparam rnode_8to10_bb4__29_i443_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_8to10_bb4__29_i443_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_8to10_bb4__29_i443_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_7to8_bb4__29_i443_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_8to10_bb4__29_i443_0_NO_SHIFT_REG = rnode_8to10_bb4__29_i443_0_reg_10_NO_SHIFT_REG;
assign rnode_8to10_bb4__29_i443_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_8to10_bb4__29_i443_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i460_stall_local;
wire [31:0] local_bb4_shr_i_i460;

assign local_bb4_shr_i_i460 = ((local_bb4_var__u29 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i15_i451_stall_local;
wire [31:0] local_bb4_shl_i15_i451;

assign local_bb4_shl_i15_i451 = ((local_bb4__tr_i450 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb4_and48_i456_stall_local;
wire [31:0] local_bb4_and48_i456;

assign local_bb4_and48_i456 = ((local_bb4__tr_i450 & 32'hFFFFFF) & 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4__29_i443_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4__29_i443_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4__29_i443_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4__29_i443_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4__29_i443_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__29_i443_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__29_i443_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__29_i443_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4__29_i443_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4__29_i443_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4__29_i443_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4__29_i443_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4__29_i443_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(rnode_8to10_bb4__29_i443_0_NO_SHIFT_REG),
	.data_out(rnode_10to11_bb4__29_i443_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4__29_i443_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4__29_i443_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4__29_i443_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4__29_i443_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4__29_i443_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_8to10_bb4__29_i443_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__29_i443_0_NO_SHIFT_REG = rnode_10to11_bb4__29_i443_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4__29_i443_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__29_i443_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_i17_i453_stall_local;
wire [31:0] local_bb4_or_i17_i453;

assign local_bb4_or_i17_i453 = ((local_bb4_shl_i15_i451 & 32'hFFFF00) | (local_bb4_shr_i16_i452 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool49_i457_stall_local;
wire local_bb4_tobool49_i457;

assign local_bb4_tobool49_i457 = ((local_bb4_and48_i456 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_i459_stall_local;
wire [31:0] local_bb4_shl_i_i459;

assign local_bb4_shl_i_i459 = ((local_bb4_or_i17_i453 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__31_i464_stall_local;
wire local_bb4__31_i464;

assign local_bb4__31_i464 = (local_bb4_tobool49_i457 & local_bb4_cmp50_not_i463);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i461_stall_local;
wire [31:0] local_bb4_or_i_i461;

assign local_bb4_or_i_i461 = ((local_bb4_shl_i_i459 & 32'h1FFFFFE) | (local_bb4_shr_i_i460 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i465_stall_local;
wire [31:0] local_bb4__32_i465;

assign local_bb4__32_i465 = (local_bb4__31_i464 ? (local_bb4_shl1_i_i462 & 32'hFFFFFE00) : (local_bb4_shl1_i18_i454 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__36_i469_stall_local;
wire [31:0] local_bb4__36_i469;

assign local_bb4__36_i469 = (local_bb4__31_i464 ? (rnode_8to9_bb4_add_i455_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4__34_i467_stall_local;
wire [31:0] local_bb4__34_i467;

assign local_bb4__34_i467 = (local_bb4__31_i464 ? (local_bb4_or_i_i461 & 32'h1FFFFFF) : (local_bb4_or_i17_i453 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i466_stall_local;
wire [31:0] local_bb4__33_i466;

assign local_bb4__33_i466 = (local_bb4_tobool49_i457 ? (local_bb4__32_i465 & 32'hFFFFFF00) : (local_bb4_shl1_i18_i454 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__37_i470_stall_local;
wire [31:0] local_bb4__37_i470;

assign local_bb4__37_i470 = (local_bb4_tobool49_i457 ? (local_bb4__36_i469 & 32'h1FF) : (local_bb4_inc_i458 & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb4__35_i468_stall_local;
wire [31:0] local_bb4__35_i468;

assign local_bb4__35_i468 = (local_bb4_tobool49_i457 ? (local_bb4__34_i467 & 32'h1FFFFFF) : (local_bb4_or_i17_i453 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp53_i471_stall_local;
wire local_bb4_cmp53_i471;

assign local_bb4_cmp53_i471 = ((local_bb4__37_i470 & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp68_i475_stall_local;
wire local_bb4_cmp68_i475;

assign local_bb4_cmp68_i475 = ((local_bb4__37_i470 & 32'h3FF) < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i477_stall_local;
wire [31:0] local_bb4_sub_i477;

assign local_bb4_sub_i477 = ((local_bb4__37_i470 & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp71_not_i492_stall_local;
wire local_bb4_cmp71_not_i492;

assign local_bb4_cmp71_not_i492 = ((local_bb4__37_i470 & 32'h3FF) != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i476_stall_local;
wire [31:0] local_bb4_and75_i476;

assign local_bb4_and75_i476 = ((local_bb4__35_i468 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and83_i482_stall_local;
wire [31:0] local_bb4_and83_i482;

assign local_bb4_and83_i482 = ((local_bb4__35_i468 & 32'h1FFFFFF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or581_i472_stall_local;
wire local_bb4_or581_i472;

assign local_bb4_or581_i472 = (rnode_8to9_bb4_var__u26_0_NO_SHIFT_REG | local_bb4_cmp53_i471);

// This section implements an unregistered operation.
// 
wire local_bb4_and74_i478_stall_local;
wire [31:0] local_bb4_and74_i478;

assign local_bb4_and74_i478 = ((local_bb4_sub_i477 & 32'hFF800000) + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i466_valid_out;
wire local_bb4__33_i466_stall_in;
wire local_bb4_cmp68_i475_valid_out;
wire local_bb4_cmp68_i475_stall_in;
wire local_bb4_cmp71_not_i492_valid_out;
wire local_bb4_cmp71_not_i492_stall_in;
wire local_bb4_and75_i476_valid_out;
wire local_bb4_and75_i476_stall_in;
wire local_bb4_and83_i482_valid_out;
wire local_bb4_and83_i482_stall_in;
wire local_bb4_or581_i472_valid_out;
wire local_bb4_or581_i472_stall_in;
wire local_bb4_shl_i479_valid_out;
wire local_bb4_shl_i479_stall_in;
wire local_bb4_shl_i479_inputs_ready;
wire local_bb4_shl_i479_stall_local;
wire [31:0] local_bb4_shl_i479;

assign local_bb4_shl_i479_inputs_ready = (local_bb4_mul_i_i448_valid_out_0_NO_SHIFT_REG & local_bb4_mul_i_i448_valid_out_1_NO_SHIFT_REG & rnode_8to9_bb4_add_i455_0_valid_out_1_NO_SHIFT_REG & rnode_8to9_bb4_add_i455_0_valid_out_0_NO_SHIFT_REG & rnode_8to9_bb4_add_i455_0_valid_out_2_NO_SHIFT_REG & rnode_8to9_bb4_var__u26_0_valid_out_NO_SHIFT_REG);
assign local_bb4_shl_i479 = ((local_bb4_and74_i478 & 32'hFF800000) & 32'h7F800000);
assign local_bb4__33_i466_valid_out = 1'b1;
assign local_bb4_cmp68_i475_valid_out = 1'b1;
assign local_bb4_cmp71_not_i492_valid_out = 1'b1;
assign local_bb4_and75_i476_valid_out = 1'b1;
assign local_bb4_and83_i482_valid_out = 1'b1;
assign local_bb4_or581_i472_valid_out = 1'b1;
assign local_bb4_shl_i479_valid_out = 1'b1;
assign local_bb4_mul_i_i448_stall_in_0 = 1'b0;
assign local_bb4_mul_i_i448_stall_in_1 = 1'b0;
assign rnode_8to9_bb4_add_i455_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_add_i455_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_add_i455_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_8to9_bb4_var__u26_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4__33_i466_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4__33_i466_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4__33_i466_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4__33_i466_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4__33_i466_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4__33_i466_1_NO_SHIFT_REG;
 logic rnode_9to10_bb4__33_i466_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4__33_i466_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4__33_i466_0_valid_out_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4__33_i466_0_stall_in_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4__33_i466_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4__33_i466_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4__33_i466_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4__33_i466_0_stall_in_0_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4__33_i466_0_valid_out_0_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4__33_i466_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in((local_bb4__33_i466 & 32'hFFFFFF00)),
	.data_out(rnode_9to10_bb4__33_i466_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4__33_i466_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4__33_i466_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4__33_i466_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4__33_i466_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4__33_i466_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__33_i466_stall_in = 1'b0;
assign rnode_9to10_bb4__33_i466_0_stall_in_0_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4__33_i466_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4__33_i466_0_NO_SHIFT_REG = rnode_9to10_bb4__33_i466_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4__33_i466_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_9to10_bb4__33_i466_1_NO_SHIFT_REG = rnode_9to10_bb4__33_i466_0_reg_10_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_9to11_bb4_cmp68_i475_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp68_i475_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp68_i475_0_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp68_i475_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp68_i475_0_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp68_i475_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp68_i475_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp68_i475_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_9to11_bb4_cmp68_i475_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to11_bb4_cmp68_i475_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to11_bb4_cmp68_i475_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_9to11_bb4_cmp68_i475_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_9to11_bb4_cmp68_i475_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_cmp68_i475),
	.data_out(rnode_9to11_bb4_cmp68_i475_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_9to11_bb4_cmp68_i475_0_reg_11_fifo.DEPTH = 2;
defparam rnode_9to11_bb4_cmp68_i475_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_9to11_bb4_cmp68_i475_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to11_bb4_cmp68_i475_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_9to11_bb4_cmp68_i475_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp68_i475_stall_in = 1'b0;
assign rnode_9to11_bb4_cmp68_i475_0_NO_SHIFT_REG = rnode_9to11_bb4_cmp68_i475_0_reg_11_NO_SHIFT_REG;
assign rnode_9to11_bb4_cmp68_i475_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_cmp68_i475_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_9to11_bb4_cmp71_not_i492_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp71_not_i492_0_stall_in_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp71_not_i492_0_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp71_not_i492_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp71_not_i492_0_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp71_not_i492_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp71_not_i492_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_cmp71_not_i492_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_9to11_bb4_cmp71_not_i492_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to11_bb4_cmp71_not_i492_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to11_bb4_cmp71_not_i492_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_9to11_bb4_cmp71_not_i492_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_9to11_bb4_cmp71_not_i492_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_cmp71_not_i492),
	.data_out(rnode_9to11_bb4_cmp71_not_i492_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_9to11_bb4_cmp71_not_i492_0_reg_11_fifo.DEPTH = 2;
defparam rnode_9to11_bb4_cmp71_not_i492_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_9to11_bb4_cmp71_not_i492_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to11_bb4_cmp71_not_i492_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_9to11_bb4_cmp71_not_i492_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp71_not_i492_stall_in = 1'b0;
assign rnode_9to11_bb4_cmp71_not_i492_0_NO_SHIFT_REG = rnode_9to11_bb4_cmp71_not_i492_0_reg_11_NO_SHIFT_REG;
assign rnode_9to11_bb4_cmp71_not_i492_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_cmp71_not_i492_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_and75_i476_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and75_i476_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_and75_i476_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and75_i476_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_and75_i476_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and75_i476_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and75_i476_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and75_i476_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_and75_i476_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_and75_i476_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_and75_i476_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_and75_i476_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_and75_i476_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in((local_bb4_and75_i476 & 32'h7FFFFF)),
	.data_out(rnode_9to10_bb4_and75_i476_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_and75_i476_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_and75_i476_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_and75_i476_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_and75_i476_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_and75_i476_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and75_i476_stall_in = 1'b0;
assign rnode_9to10_bb4_and75_i476_0_NO_SHIFT_REG = rnode_9to10_bb4_and75_i476_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_and75_i476_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_and75_i476_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_and83_i482_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and83_i482_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_and83_i482_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and83_i482_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_and83_i482_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and83_i482_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and83_i482_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_and83_i482_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_and83_i482_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_and83_i482_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_and83_i482_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_and83_i482_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_and83_i482_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in((local_bb4_and83_i482 & 32'h1)),
	.data_out(rnode_9to10_bb4_and83_i482_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_and83_i482_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_and83_i482_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_and83_i482_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_and83_i482_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_and83_i482_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and83_i482_stall_in = 1'b0;
assign rnode_9to10_bb4_and83_i482_0_NO_SHIFT_REG = rnode_9to10_bb4_and83_i482_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_and83_i482_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_and83_i482_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_9to11_bb4_or581_i472_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_1_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_valid_out_0_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_stall_in_0_reg_11_NO_SHIFT_REG;
 logic rnode_9to11_bb4_or581_i472_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_9to11_bb4_or581_i472_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to11_bb4_or581_i472_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to11_bb4_or581_i472_0_stall_in_0_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_9to11_bb4_or581_i472_0_valid_out_0_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_9to11_bb4_or581_i472_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4_or581_i472),
	.data_out(rnode_9to11_bb4_or581_i472_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_9to11_bb4_or581_i472_0_reg_11_fifo.DEPTH = 2;
defparam rnode_9to11_bb4_or581_i472_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_9to11_bb4_or581_i472_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to11_bb4_or581_i472_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_9to11_bb4_or581_i472_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or581_i472_stall_in = 1'b0;
assign rnode_9to11_bb4_or581_i472_0_stall_in_0_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_or581_i472_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_9to11_bb4_or581_i472_0_NO_SHIFT_REG = rnode_9to11_bb4_or581_i472_0_reg_11_NO_SHIFT_REG;
assign rnode_9to11_bb4_or581_i472_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_9to11_bb4_or581_i472_1_NO_SHIFT_REG = rnode_9to11_bb4_or581_i472_0_reg_11_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_9to10_bb4_shl_i479_0_valid_out_NO_SHIFT_REG;
 logic rnode_9to10_bb4_shl_i479_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_shl_i479_0_NO_SHIFT_REG;
 logic rnode_9to10_bb4_shl_i479_0_reg_10_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_9to10_bb4_shl_i479_0_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_shl_i479_0_valid_out_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_shl_i479_0_stall_in_reg_10_NO_SHIFT_REG;
 logic rnode_9to10_bb4_shl_i479_0_stall_out_reg_10_NO_SHIFT_REG;

acl_data_fifo rnode_9to10_bb4_shl_i479_0_reg_10_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_9to10_bb4_shl_i479_0_reg_10_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_9to10_bb4_shl_i479_0_stall_in_reg_10_NO_SHIFT_REG),
	.valid_out(rnode_9to10_bb4_shl_i479_0_valid_out_reg_10_NO_SHIFT_REG),
	.stall_out(rnode_9to10_bb4_shl_i479_0_stall_out_reg_10_NO_SHIFT_REG),
	.data_in((local_bb4_shl_i479 & 32'h7F800000)),
	.data_out(rnode_9to10_bb4_shl_i479_0_reg_10_NO_SHIFT_REG)
);

defparam rnode_9to10_bb4_shl_i479_0_reg_10_fifo.DEPTH = 1;
defparam rnode_9to10_bb4_shl_i479_0_reg_10_fifo.DATA_WIDTH = 32;
defparam rnode_9to10_bb4_shl_i479_0_reg_10_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_9to10_bb4_shl_i479_0_reg_10_fifo.IMPL = "shift_reg";

assign rnode_9to10_bb4_shl_i479_0_reg_10_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shl_i479_stall_in = 1'b0;
assign rnode_9to10_bb4_shl_i479_0_NO_SHIFT_REG = rnode_9to10_bb4_shl_i479_0_reg_10_NO_SHIFT_REG;
assign rnode_9to10_bb4_shl_i479_0_stall_in_reg_10_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_shl_i479_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i481_stall_local;
wire local_bb4_cmp77_i481;

assign local_bb4_cmp77_i481 = ((rnode_9to10_bb4__33_i466_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u30_stall_local;
wire local_bb4_var__u30;

assign local_bb4_var__u30 = ($signed((rnode_9to10_bb4__33_i466_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u31_stall_local;
wire [31:0] local_bb4_var__u31;

assign local_bb4_var__u31[31:1] = 31'h0;
assign local_bb4_var__u31[0] = rnode_9to11_bb4_cmp68_i475_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool84_i483_stall_local;
wire local_bb4_tobool84_i483;

assign local_bb4_tobool84_i483 = ((rnode_9to10_bb4_and83_i482_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i474_stall_local;
wire local_bb4_reduction_2_i474;

assign local_bb4_reduction_2_i474 = (rnode_10to11_bb4_reduction_0_i473_0_NO_SHIFT_REG | rnode_9to11_bb4_or581_i472_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cond111_i500_stall_local;
wire [31:0] local_bb4_cond111_i500;

assign local_bb4_cond111_i500 = (rnode_9to11_bb4_or581_i472_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or76_i480_valid_out;
wire local_bb4_or76_i480_stall_in;
wire local_bb4_or76_i480_inputs_ready;
wire local_bb4_or76_i480_stall_local;
wire [31:0] local_bb4_or76_i480;

assign local_bb4_or76_i480_inputs_ready = (rnode_9to10_bb4_shl_i479_0_valid_out_NO_SHIFT_REG & rnode_9to10_bb4_and75_i476_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or76_i480 = ((rnode_9to10_bb4_shl_i479_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_9to10_bb4_and75_i476_0_NO_SHIFT_REG & 32'h7FFFFF));
assign local_bb4_or76_i480_valid_out = 1'b1;
assign rnode_9to10_bb4_shl_i479_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_and75_i476_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__39_i484_stall_local;
wire local_bb4__39_i484;

assign local_bb4__39_i484 = (local_bb4_tobool84_i483 & local_bb4_var__u30);

// This section implements an unregistered operation.
// 
wire local_bb4_conv101_i495_stall_local;
wire [31:0] local_bb4_conv101_i495;

assign local_bb4_conv101_i495[31:1] = 31'h0;
assign local_bb4_conv101_i495[0] = local_bb4_reduction_2_i474;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4_or76_i480_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4_or76_i480_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_or76_i480_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4_or76_i480_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_10to11_bb4_or76_i480_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_or76_i480_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_or76_i480_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4_or76_i480_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4_or76_i480_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4_or76_i480_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4_or76_i480_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4_or76_i480_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4_or76_i480_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in((local_bb4_or76_i480 & 32'h7FFFFFFF)),
	.data_out(rnode_10to11_bb4_or76_i480_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4_or76_i480_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4_or76_i480_0_reg_11_fifo.DATA_WIDTH = 32;
defparam rnode_10to11_bb4_or76_i480_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4_or76_i480_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4_or76_i480_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or76_i480_stall_in = 1'b0;
assign rnode_10to11_bb4_or76_i480_0_NO_SHIFT_REG = rnode_10to11_bb4_or76_i480_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4_or76_i480_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_or76_i480_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__40_i485_valid_out;
wire local_bb4__40_i485_stall_in;
wire local_bb4__40_i485_inputs_ready;
wire local_bb4__40_i485_stall_local;
wire local_bb4__40_i485;

assign local_bb4__40_i485_inputs_ready = (rnode_9to10_bb4__33_i466_0_valid_out_0_NO_SHIFT_REG & rnode_9to10_bb4__33_i466_0_valid_out_1_NO_SHIFT_REG & rnode_9to10_bb4_and83_i482_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40_i485 = (local_bb4_cmp77_i481 | local_bb4__39_i484);
assign local_bb4__40_i485_valid_out = 1'b1;
assign rnode_9to10_bb4__33_i466_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4__33_i466_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_9to10_bb4_and83_i482_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_10to11_bb4__40_i485_0_valid_out_NO_SHIFT_REG;
 logic rnode_10to11_bb4__40_i485_0_stall_in_NO_SHIFT_REG;
 logic rnode_10to11_bb4__40_i485_0_NO_SHIFT_REG;
 logic rnode_10to11_bb4__40_i485_0_reg_11_inputs_ready_NO_SHIFT_REG;
 logic rnode_10to11_bb4__40_i485_0_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__40_i485_0_valid_out_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__40_i485_0_stall_in_reg_11_NO_SHIFT_REG;
 logic rnode_10to11_bb4__40_i485_0_stall_out_reg_11_NO_SHIFT_REG;

acl_data_fifo rnode_10to11_bb4__40_i485_0_reg_11_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_10to11_bb4__40_i485_0_reg_11_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_10to11_bb4__40_i485_0_stall_in_reg_11_NO_SHIFT_REG),
	.valid_out(rnode_10to11_bb4__40_i485_0_valid_out_reg_11_NO_SHIFT_REG),
	.stall_out(rnode_10to11_bb4__40_i485_0_stall_out_reg_11_NO_SHIFT_REG),
	.data_in(local_bb4__40_i485),
	.data_out(rnode_10to11_bb4__40_i485_0_reg_11_NO_SHIFT_REG)
);

defparam rnode_10to11_bb4__40_i485_0_reg_11_fifo.DEPTH = 1;
defparam rnode_10to11_bb4__40_i485_0_reg_11_fifo.DATA_WIDTH = 1;
defparam rnode_10to11_bb4__40_i485_0_reg_11_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_10to11_bb4__40_i485_0_reg_11_fifo.IMPL = "shift_reg";

assign rnode_10to11_bb4__40_i485_0_reg_11_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_i485_stall_in = 1'b0;
assign rnode_10to11_bb4__40_i485_0_NO_SHIFT_REG = rnode_10to11_bb4__40_i485_0_reg_11_NO_SHIFT_REG;
assign rnode_10to11_bb4__40_i485_0_stall_in_reg_11_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__40_i485_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cond_i486_stall_local;
wire [31:0] local_bb4_cond_i486;

assign local_bb4_cond_i486[31:1] = 31'h0;
assign local_bb4_cond_i486[0] = rnode_10to11_bb4__40_i485_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add87_i487_stall_local;
wire [31:0] local_bb4_add87_i487;

assign local_bb4_add87_i487 = ((local_bb4_cond_i486 & 32'h1) + (rnode_10to11_bb4_or76_i480_0_NO_SHIFT_REG & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i488_stall_local;
wire [31:0] local_bb4_and88_i488;

assign local_bb4_and88_i488 = (local_bb4_add87_i487 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i490_stall_local;
wire [31:0] local_bb4_and90_i490;

assign local_bb4_and90_i490 = (local_bb4_add87_i487 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_or89_i489_stall_local;
wire [31:0] local_bb4_or89_i489;

assign local_bb4_or89_i489 = ((local_bb4_and88_i488 & 32'h7FFFFFFF) | (local_bb4_and4_i415 & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i491_stall_local;
wire local_bb4_cmp91_i491;

assign local_bb4_cmp91_i491 = ((local_bb4_and90_i490 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge14_i493_stall_local;
wire local_bb4_brmerge14_i493;

assign local_bb4_brmerge14_i493 = (local_bb4_cmp91_i491 | rnode_9to11_bb4_cmp71_not_i492_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_conv99_i494_stall_local;
wire [31:0] local_bb4_conv99_i494;

assign local_bb4_conv99_i494 = (local_bb4_brmerge14_i493 ? (local_bb4_var__u31 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or102_i496_stall_local;
wire [31:0] local_bb4_or102_i496;

assign local_bb4_or102_i496 = ((local_bb4_conv99_i494 & 32'h1) | (local_bb4_conv101_i495 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool103_i497_stall_local;
wire local_bb4_tobool103_i497;

assign local_bb4_tobool103_i497 = ((local_bb4_or102_i496 & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cond107_i498_stall_local;
wire [31:0] local_bb4_cond107_i498;

assign local_bb4_cond107_i498 = (local_bb4_tobool103_i497 ? (local_bb4_and4_i415 & 32'h80000000) : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and108_i499_stall_local;
wire [31:0] local_bb4_and108_i499;

assign local_bb4_and108_i499 = (local_bb4_cond107_i498 & local_bb4_or89_i489);

// This section implements an unregistered operation.
// 
wire local_bb4_or112_i501_stall_local;
wire [31:0] local_bb4_or112_i501;

assign local_bb4_or112_i501 = (local_bb4_and108_i499 | (local_bb4_cond111_i500 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u32_stall_local;
wire [31:0] local_bb4_var__u32;

assign local_bb4_var__u32 = local_bb4_or112_i501;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u33_stall_local;
wire [31:0] local_bb4_var__u33;

assign local_bb4_var__u33 = (rnode_10to11_bb4__29_i443_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb4_var__u32);

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi225_stall_local;
wire [191:0] local_bb4_c0_exi225;

assign local_bb4_c0_exi225[127:0] = local_bb4_c0_exi124[127:0];
assign local_bb4_c0_exi225[159:128] = local_bb4_var__u33;
assign local_bb4_c0_exi225[191:160] = local_bb4_c0_exi124[191:160];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi326_stall_local;
wire [191:0] local_bb4_c0_exi326;

assign local_bb4_c0_exi326[159:0] = local_bb4_c0_exi225[159:0];
assign local_bb4_c0_exi326[160] = rnode_10to11_bb4_var__u22_0_NO_SHIFT_REG;
assign local_bb4_c0_exi326[191:161] = local_bb4_c0_exi225[191:161];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi427_stall_local;
wire [191:0] local_bb4_c0_exi427;

assign local_bb4_c0_exi427[167:0] = local_bb4_c0_exi326[167:0];
assign local_bb4_c0_exi427[168] = rnode_10to11_bb4_notexitcond_notexit_0_NO_SHIFT_REG;
assign local_bb4_c0_exi427[191:169] = local_bb4_c0_exi326[191:169];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi5_stall_local;
wire [191:0] local_bb4_c0_exi5;

assign local_bb4_c0_exi5[175:0] = local_bb4_c0_exi427[175:0];
assign local_bb4_c0_exi5[176] = rnode_10to11_bb4__pop12_c0_ene4_0_NO_SHIFT_REG;
assign local_bb4_c0_exi5[191:177] = local_bb4_c0_exi427[191:177];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exi6_valid_out;
wire local_bb4_c0_exi6_stall_in;
wire local_bb4_c0_exi6_inputs_ready;
wire local_bb4_c0_exi6_stall_local;
wire [191:0] local_bb4_c0_exi6;

assign local_bb4_c0_exi6_inputs_ready = (rnode_10to11_bb4__pop12_c0_ene4_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_var__u22_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_notexitcond_notexit_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_arrayidx33_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_xor_i414_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4__29_i443_0_valid_out_NO_SHIFT_REG & rnode_9to11_bb4_or581_i472_0_valid_out_1_NO_SHIFT_REG & rnode_9to11_bb4_or581_i472_0_valid_out_0_NO_SHIFT_REG & rnode_10to11_bb4_reduction_0_i473_0_valid_out_NO_SHIFT_REG & rnode_9to11_bb4_cmp68_i475_0_valid_out_NO_SHIFT_REG & rnode_9to11_bb4_cmp71_not_i492_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4__40_i485_0_valid_out_NO_SHIFT_REG & rnode_10to11_bb4_or76_i480_0_valid_out_NO_SHIFT_REG);
assign local_bb4_c0_exi6[183:0] = local_bb4_c0_exi5[183:0];
assign local_bb4_c0_exi6[184] = rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_NO_SHIFT_REG;
assign local_bb4_c0_exi6[191:185] = local_bb4_c0_exi5[191:185];
assign local_bb4_c0_exi6_valid_out = 1'b1;
assign rnode_10to11_bb4__pop12_c0_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond1520_pop13_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_var__u22_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_notexitcond_notexit_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_arrayidx33_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_xor_i414_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__29_i443_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_or581_i472_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_or581_i472_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_reduction_0_i473_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_cmp68_i475_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_9to11_bb4_cmp71_not_i492_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4__40_i485_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_or76_i480_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_c0_exit28_c0_exi6_inputs_ready;
 reg local_bb4_c0_exit28_c0_exi6_valid_out_0_NO_SHIFT_REG;
wire local_bb4_c0_exit28_c0_exi6_stall_in_0;
 reg local_bb4_c0_exit28_c0_exi6_valid_out_1_NO_SHIFT_REG;
wire local_bb4_c0_exit28_c0_exi6_stall_in_1;
 reg [191:0] local_bb4_c0_exit28_c0_exi6_NO_SHIFT_REG;
wire [191:0] local_bb4_c0_exit28_c0_exi6_in;
wire local_bb4_c0_exit28_c0_exi6_valid;
wire local_bb4_c0_exit28_c0_exi6_causedstall;

acl_stall_free_sink local_bb4_c0_exit28_c0_exi6_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb4_c0_exi6),
	.data_out(local_bb4_c0_exit28_c0_exi6_in),
	.input_accepted(local_bb4_c0_enter22_c0_eni5_input_accepted),
	.valid_out(local_bb4_c0_exit28_c0_exi6_valid),
	.stall_in(~(local_bb4_c0_exit28_c0_exi6_output_regs_ready)),
	.stall_entry(local_bb4_c0_exit28_c0_exi6_entry_stall),
	.valid_in(local_bb4_c0_exit28_c0_exi6_valid_in),
	.IIphases(local_bb4_c0_exit28_c0_exi6_phases),
	.inc_pipelined_thread(local_bb4_c0_enter22_c0_eni5_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb4_c0_enter22_c0_eni5_dec_pipelined_thread)
);

defparam local_bb4_c0_exit28_c0_exi6_instance.DATA_WIDTH = 192;
defparam local_bb4_c0_exit28_c0_exi6_instance.PIPELINE_DEPTH = 15;
defparam local_bb4_c0_exit28_c0_exi6_instance.SHARINGII = 1;
defparam local_bb4_c0_exit28_c0_exi6_instance.SCHEDULEII = 1;
defparam local_bb4_c0_exit28_c0_exi6_instance.ALWAYS_THROTTLE = 0;

assign local_bb4_c0_exit28_c0_exi6_inputs_ready = 1'b1;
assign local_bb4_c0_exit28_c0_exi6_output_regs_ready = ((~(local_bb4_c0_exit28_c0_exi6_valid_out_0_NO_SHIFT_REG) | ~(local_bb4_c0_exit28_c0_exi6_stall_in_0)) & (~(local_bb4_c0_exit28_c0_exi6_valid_out_1_NO_SHIFT_REG) | ~(local_bb4_c0_exit28_c0_exi6_stall_in_1)));
assign local_bb4_c0_exit28_c0_exi6_valid_in = SFC_2_VALID_10_11_0_NO_SHIFT_REG;
assign local_bb4_c0_exi6_stall_in = 1'b0;
assign local_bb4_gaussian_ROM4119_push11_gaussian_ROM4119_pop11_stall_in = 1'b0;
assign local_bb4_sub24_add2318_push10_sub24_add2318_pop10_stall_in = 1'b0;
assign local_bb4__push12__pop12_stall_in = 1'b0;
assign local_bb4_notexitcond1520_push13_notexitcond1520_pop13_stall_in = 1'b0;
assign SFC_2_VALID_10_11_0_stall_in = 1'b0;
assign rnode_10to11_bb4_keep_going_acl_pipeline_1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_10to11_bb4_indvars_iv_push7_indvars_iv_next_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_c0_exit28_c0_exi6_causedstall = (1'b1 && (1'b0 && !(~(local_bb4_c0_exit28_c0_exi6_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c0_exit28_c0_exi6_NO_SHIFT_REG <= 'x;
		local_bb4_c0_exit28_c0_exi6_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_c0_exit28_c0_exi6_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c0_exit28_c0_exi6_output_regs_ready)
		begin
			local_bb4_c0_exit28_c0_exi6_NO_SHIFT_REG <= local_bb4_c0_exit28_c0_exi6_in;
			local_bb4_c0_exit28_c0_exi6_valid_out_0_NO_SHIFT_REG <= local_bb4_c0_exit28_c0_exi6_valid;
			local_bb4_c0_exit28_c0_exi6_valid_out_1_NO_SHIFT_REG <= local_bb4_c0_exit28_c0_exi6_valid;
		end
		else
		begin
			if (~(local_bb4_c0_exit28_c0_exi6_stall_in_0))
			begin
				local_bb4_c0_exit28_c0_exi6_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c0_exit28_c0_exi6_stall_in_1))
			begin
				local_bb4_c0_exit28_c0_exi6_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe129_valid_out;
wire local_bb4_c0_exe129_stall_in;
wire local_bb4_c0_exe129_inputs_ready;
wire local_bb4_c0_exe129_stall_local;
wire [63:0] local_bb4_c0_exe129;

assign local_bb4_c0_exe129_inputs_ready = local_bb4_c0_exit28_c0_exi6_valid_out_0_NO_SHIFT_REG;
assign local_bb4_c0_exe129 = local_bb4_c0_exit28_c0_exi6_NO_SHIFT_REG[127:64];
assign local_bb4_c0_exe129_valid_out = local_bb4_c0_exe129_inputs_ready;
assign local_bb4_c0_exe129_stall_local = local_bb4_c0_exe129_stall_in;
assign local_bb4_c0_exit28_c0_exi6_stall_in_0 = (|local_bb4_c0_exe129_stall_local);

// Register node:
//  * latency = 159
//  * capacity = 159
 logic rnode_16to175_bb4_c0_exit28_c0_exi6_0_valid_out_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_in_NO_SHIFT_REG;
 logic [191:0] rnode_16to175_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [191:0] rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit28_c0_exi6_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_16to175_bb4_c0_exit28_c0_exi6_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb4_c0_exit28_c0_exi6_NO_SHIFT_REG),
	.data_out(rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_fifo.DEPTH = 160;
defparam rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_fifo.DATA_WIDTH = 192;
defparam rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_fifo.IMPL = "ram";

assign rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_inputs_ready_NO_SHIFT_REG = local_bb4_c0_exit28_c0_exi6_valid_out_1_NO_SHIFT_REG;
assign local_bb4_c0_exit28_c0_exi6_stall_in_1 = rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_out_reg_175_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit28_c0_exi6_0_reg_175_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_in_reg_175_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_in_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit28_c0_exi6_0_valid_out_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit28_c0_exi6_0_valid_out_reg_175_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_ld__inputs_ready;
 reg local_bb4_ld__valid_out_NO_SHIFT_REG;
wire local_bb4_ld__stall_in;
wire local_bb4_ld__output_regs_ready;
wire local_bb4_ld__fu_stall_out;
wire local_bb4_ld__fu_valid_out;
wire [31:0] local_bb4_ld__lsu_dataout;
 reg [31:0] local_bb4_ld__NO_SHIFT_REG;
wire local_bb4_ld__causedstall;

lsu_top lsu_local_bb4_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb4_ld__fu_stall_out),
	.i_valid(local_bb4_ld__inputs_ready),
	.i_address((local_bb4_c0_exe129 & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(local_bb4__acl_ffwd_dest_i1_9),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb4_ld__output_regs_ready)),
	.o_valid(local_bb4_ld__fu_valid_out),
	.o_readdata(local_bb4_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb4_ld__active),
	.avm_address(avm_local_bb4_ld__address),
	.avm_read(avm_local_bb4_ld__read),
	.avm_readdata(avm_local_bb4_ld__readdata),
	.avm_write(avm_local_bb4_ld__write),
	.avm_writeack(avm_local_bb4_ld__writeack),
	.avm_burstcount(avm_local_bb4_ld__burstcount),
	.avm_writedata(avm_local_bb4_ld__writedata),
	.avm_byteenable(avm_local_bb4_ld__byteenable),
	.avm_waitrequest(avm_local_bb4_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb4_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb4_ld_.AWIDTH = 33;
defparam lsu_local_bb4_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb4_ld_.MWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb4_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb4_ld_.READ = 1;
defparam lsu_local_bb4_ld_.ATOMIC = 0;
defparam lsu_local_bb4_ld_.WIDTH = 32;
defparam lsu_local_bb4_ld_.MWIDTH = 512;
defparam lsu_local_bb4_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb4_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb4_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb4_ld_.MEMORY_SIDE_MEM_LATENCY = 115;
defparam lsu_local_bb4_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb4_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb4_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb4_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb4_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb4_ld_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb4_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb4_ld_.USECACHING = 1;
defparam lsu_local_bb4_ld_.CACHESIZE = 1024;
defparam lsu_local_bb4_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb4_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb4_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb4_ld_.ADDRSPACE = 1;
defparam lsu_local_bb4_ld_.STYLE = "BURST-COALESCED";

assign local_bb4_ld__inputs_ready = (local_bb4_c0_exe129_valid_out & local_bb4__acl_ffwd_dest_i1_9_valid_out);
assign local_bb4_ld__output_regs_ready = (&(~(local_bb4_ld__valid_out_NO_SHIFT_REG) | ~(local_bb4_ld__stall_in)));
assign local_bb4_c0_exe129_stall_in = (local_bb4_ld__fu_stall_out | ~(local_bb4_ld__inputs_ready));
assign local_bb4__acl_ffwd_dest_i1_9_stall_in = (local_bb4_ld__fu_stall_out | ~(local_bb4_ld__inputs_ready));
assign local_bb4_ld__causedstall = (local_bb4_ld__inputs_ready && (local_bb4_ld__fu_stall_out && !(~(local_bb4_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_ld__NO_SHIFT_REG <= 'x;
		local_bb4_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_ld__output_regs_ready)
		begin
			local_bb4_ld__NO_SHIFT_REG <= local_bb4_ld__lsu_dataout;
			local_bb4_ld__valid_out_NO_SHIFT_REG <= local_bb4_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb4_ld__stall_in))
			begin
				local_bb4_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_NO_SHIFT_REG;
 logic [191:0] rnode_175to176_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_1_NO_SHIFT_REG;
 logic [191:0] rnode_175to176_bb4_c0_exit28_c0_exi6_1_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_2_NO_SHIFT_REG;
 logic [191:0] rnode_175to176_bb4_c0_exit28_c0_exi6_2_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [191:0] rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_out_reg_176_NO_SHIFT_REG;
 reg rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_0_NO_SHIFT_REG;
 reg rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_2_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_16to175_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_fifo.DATA_WIDTH = 192;
defparam rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_fifo.IMPL = "ll_reg";

assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_inputs_ready_NO_SHIFT_REG = rnode_16to175_bb4_c0_exit28_c0_exi6_0_valid_out_NO_SHIFT_REG;
assign rnode_16to175_bb4_c0_exit28_c0_exi6_0_stall_in_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_out_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_176_NO_SHIFT_REG = ((rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_0_NO_SHIFT_REG)) | 1'b0 | (rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_2_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_2_NO_SHIFT_REG)));
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_NO_SHIFT_REG = (rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_176_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_0_NO_SHIFT_REG));
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_1_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_2_NO_SHIFT_REG = (rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_176_NO_SHIFT_REG & ~(rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_2_NO_SHIFT_REG));
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit28_c0_exi6_1_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit28_c0_exi6_2_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit28_c0_exi6_0_reg_176_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_0_NO_SHIFT_REG <= (rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_176_NO_SHIFT_REG & (rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_0_NO_SHIFT_REG | ~(rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_NO_SHIFT_REG)) & rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_176_NO_SHIFT_REG);
		rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_2_NO_SHIFT_REG <= (rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_176_NO_SHIFT_REG & (rnode_175to176_bb4_c0_exit28_c0_exi6_0_consumed_2_NO_SHIFT_REG | ~(rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_2_NO_SHIFT_REG)) & rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_176_NO_SHIFT_REG);
	end
end


// This section implements a staging register.
// 
wire rstag_176to176_bb4_ld__valid_out;
wire rstag_176to176_bb4_ld__stall_in;
wire rstag_176to176_bb4_ld__inputs_ready;
wire rstag_176to176_bb4_ld__stall_local;
 reg rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG;
wire rstag_176to176_bb4_ld__combined_valid;
 reg [31:0] rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_176to176_bb4_ld_;

assign rstag_176to176_bb4_ld__inputs_ready = local_bb4_ld__valid_out_NO_SHIFT_REG;
assign rstag_176to176_bb4_ld_ = (rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG ? rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG : local_bb4_ld__NO_SHIFT_REG);
assign rstag_176to176_bb4_ld__combined_valid = (rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG | rstag_176to176_bb4_ld__inputs_ready);
assign rstag_176to176_bb4_ld__valid_out = rstag_176to176_bb4_ld__combined_valid;
assign rstag_176to176_bb4_ld__stall_local = rstag_176to176_bb4_ld__stall_in;
assign local_bb4_ld__stall_in = (|rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_176to176_bb4_ld__stall_local)
		begin
			if (~(rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= rstag_176to176_bb4_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_176to176_bb4_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_176to176_bb4_ld__staging_reg_NO_SHIFT_REG <= local_bb4_ld__NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe230_stall_local;
wire [31:0] local_bb4_c0_exe230;

assign local_bb4_c0_exe230 = rnode_175to176_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG[159:128];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe432_stall_local;
wire local_bb4_c0_exe432;

assign local_bb4_c0_exe432 = rnode_175to176_bb4_c0_exit28_c0_exi6_1_NO_SHIFT_REG[168];

// Register node:
//  * latency = 73
//  * capacity = 73
 logic rnode_176to249_bb4_c0_exit28_c0_exi6_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_in_NO_SHIFT_REG;
 logic [191:0] rnode_176to249_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG;
 logic rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_inputs_ready_NO_SHIFT_REG;
 logic [191:0] rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_NO_SHIFT_REG;
 logic rnode_176to249_bb4_c0_exit28_c0_exi6_0_valid_out_reg_249_NO_SHIFT_REG;
 logic rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_in_reg_249_NO_SHIFT_REG;
 logic rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_out_reg_249_NO_SHIFT_REG;

acl_data_fifo rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_in_reg_249_NO_SHIFT_REG),
	.valid_out(rnode_176to249_bb4_c0_exit28_c0_exi6_0_valid_out_reg_249_NO_SHIFT_REG),
	.stall_out(rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_out_reg_249_NO_SHIFT_REG),
	.data_in(rnode_175to176_bb4_c0_exit28_c0_exi6_2_NO_SHIFT_REG),
	.data_out(rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_NO_SHIFT_REG)
);

defparam rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_fifo.DEPTH = 74;
defparam rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_fifo.DATA_WIDTH = 192;
defparam rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_fifo.IMPL = "ram";

assign rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_inputs_ready_NO_SHIFT_REG = rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_2_NO_SHIFT_REG;
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_2_NO_SHIFT_REG = rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_out_reg_249_NO_SHIFT_REG;
assign rnode_176to249_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG = rnode_176to249_bb4_c0_exit28_c0_exi6_0_reg_249_NO_SHIFT_REG;
assign rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_in_reg_249_NO_SHIFT_REG = rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_in_NO_SHIFT_REG;
assign rnode_176to249_bb4_c0_exit28_c0_exi6_0_valid_out_NO_SHIFT_REG = rnode_176to249_bb4_c0_exit28_c0_exi6_0_valid_out_reg_249_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni1_stall_local;
wire [223:0] local_bb4_c1_eni1;

assign local_bb4_c1_eni1[31:0] = 32'bx;
assign local_bb4_c1_eni1[63:32] = rstag_176to176_bb4_ld_;
assign local_bb4_c1_eni1[223:64] = 160'bx;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_0_NO_SHIFT_REG;
 logic [191:0] rnode_249to250_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_1_NO_SHIFT_REG;
 logic [191:0] rnode_249to250_bb4_c0_exit28_c0_exi6_1_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_2_NO_SHIFT_REG;
 logic [191:0] rnode_249to250_bb4_c0_exit28_c0_exi6_2_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_inputs_ready_NO_SHIFT_REG;
 logic [191:0] rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_250_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_250_NO_SHIFT_REG;
 logic rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_out_reg_250_NO_SHIFT_REG;

acl_data_fifo rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_250_NO_SHIFT_REG),
	.valid_out(rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_250_NO_SHIFT_REG),
	.stall_out(rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_out_reg_250_NO_SHIFT_REG),
	.data_in(rnode_176to249_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG),
	.data_out(rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_NO_SHIFT_REG)
);

defparam rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_fifo.DEPTH = 1;
defparam rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_fifo.DATA_WIDTH = 192;
defparam rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_fifo.IMPL = "ll_reg";

assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_inputs_ready_NO_SHIFT_REG = rnode_176to249_bb4_c0_exit28_c0_exi6_0_valid_out_NO_SHIFT_REG;
assign rnode_176to249_bb4_c0_exit28_c0_exi6_0_stall_in_NO_SHIFT_REG = rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_out_reg_250_NO_SHIFT_REG;
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_0_reg_250_NO_SHIFT_REG = (rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_0_NO_SHIFT_REG | rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_1_NO_SHIFT_REG | rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_2_NO_SHIFT_REG);
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_NO_SHIFT_REG = rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_250_NO_SHIFT_REG;
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_1_NO_SHIFT_REG = rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_250_NO_SHIFT_REG;
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_2_NO_SHIFT_REG = rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_reg_250_NO_SHIFT_REG;
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG = rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_NO_SHIFT_REG;
assign rnode_249to250_bb4_c0_exit28_c0_exi6_1_NO_SHIFT_REG = rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_NO_SHIFT_REG;
assign rnode_249to250_bb4_c0_exit28_c0_exi6_2_NO_SHIFT_REG = rnode_249to250_bb4_c0_exit28_c0_exi6_0_reg_250_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni2_stall_local;
wire [223:0] local_bb4_c1_eni2;

assign local_bb4_c1_eni2[63:0] = local_bb4_c1_eni1[63:0];
assign local_bb4_c1_eni2[95:64] = local_bb4_c0_exe230;
assign local_bb4_c1_eni2[223:96] = local_bb4_c1_eni1[223:96];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe331_stall_local;
wire local_bb4_c0_exe331;

assign local_bb4_c0_exe331 = rnode_249to250_bb4_c0_exit28_c0_exi6_0_NO_SHIFT_REG[160];

// This section implements an unregistered operation.
// 
wire local_bb4_c0_exe6_valid_out;
wire local_bb4_c0_exe6_stall_in;
wire local_bb4_c0_exe331_valid_out;
wire local_bb4_c0_exe331_stall_in;
wire local_bb4_c0_exe6_inputs_ready;
wire local_bb4_c0_exe6_stall_local;
wire local_bb4_c0_exe6;

assign local_bb4_c0_exe6_inputs_ready = (rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_1_NO_SHIFT_REG & rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_c0_exe6 = rnode_249to250_bb4_c0_exit28_c0_exi6_1_NO_SHIFT_REG[184];
assign local_bb4_c0_exe6_stall_local = (local_bb4_c0_exe6_stall_in | local_bb4_c0_exe331_stall_in);
assign local_bb4_c0_exe6_valid_out = local_bb4_c0_exe6_inputs_ready;
assign local_bb4_c0_exe331_valid_out = local_bb4_c0_exe6_inputs_ready;
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_1_NO_SHIFT_REG = (local_bb4_c0_exe6_stall_local | ~(local_bb4_c0_exe6_inputs_ready));
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c0_exe6_stall_local | ~(local_bb4_c0_exe6_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni3_stall_local;
wire [223:0] local_bb4_c1_eni3;

assign local_bb4_c1_eni3[95:0] = local_bb4_c1_eni2[95:0];
assign local_bb4_c1_eni3[127:96] = rcnode_175to176_rc0_t_322_0_NO_SHIFT_REG[31:0];
assign local_bb4_c1_eni3[223:128] = local_bb4_c1_eni2[223:128];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni4_stall_local;
wire [223:0] local_bb4_c1_eni4;

assign local_bb4_c1_eni4[127:0] = local_bb4_c1_eni3[127:0];
assign local_bb4_c1_eni4[128] = rcnode_175to176_rc0_t_322_0_NO_SHIFT_REG[32];
assign local_bb4_c1_eni4[223:129] = local_bb4_c1_eni3[223:129];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni5_stall_local;
wire [223:0] local_bb4_c1_eni5;

assign local_bb4_c1_eni5[159:0] = local_bb4_c1_eni4[159:0];
assign local_bb4_c1_eni5[191:160] = rcnode_175to176_rc0_t_322_0_NO_SHIFT_REG[64:33];
assign local_bb4_c1_eni5[223:192] = local_bb4_c1_eni4[223:192];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_eni6_valid_out;
wire local_bb4_c1_eni6_stall_in;
wire local_bb4_c0_exe432_valid_out_1;
wire local_bb4_c0_exe432_stall_in_1;
wire local_bb4_c1_eni6_inputs_ready;
wire local_bb4_c1_eni6_stall_local;
wire [223:0] local_bb4_c1_eni6;

assign local_bb4_c1_eni6_inputs_ready = (rcnode_175to176_rc0_t_322_0_valid_out_0_NO_SHIFT_REG & rcnode_175to176_rc0_t_322_0_valid_out_1_NO_SHIFT_REG & rcnode_175to176_rc0_t_322_0_valid_out_3_NO_SHIFT_REG & rstag_176to176_bb4_ld__valid_out & rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb4_c0_exit28_c0_exi6_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_c1_eni6[191:0] = local_bb4_c1_eni5[191:0];
assign local_bb4_c1_eni6[192] = local_bb4_c0_exe432;
assign local_bb4_c1_eni6[223:193] = local_bb4_c1_eni5[223:193];
assign local_bb4_c1_eni6_stall_local = (local_bb4_c1_eni6_stall_in | local_bb4_c0_exe432_stall_in_1);
assign local_bb4_c1_eni6_valid_out = local_bb4_c1_eni6_inputs_ready;
assign local_bb4_c0_exe432_valid_out_1 = local_bb4_c1_eni6_inputs_ready;
assign rcnode_175to176_rc0_t_322_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rcnode_175to176_rc0_t_322_0_stall_in_1_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rcnode_175to176_rc0_t_322_0_stall_in_3_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rstag_176to176_bb4_ld__stall_in = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_0_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));
assign rnode_175to176_bb4_c0_exit28_c0_exi6_0_stall_in_1_NO_SHIFT_REG = (local_bb4_c1_eni6_stall_local | ~(local_bb4_c1_eni6_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb4_c1_enter_c1_eni6_inputs_ready;
 reg local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_0;
 reg local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_1;
 reg local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_2;
 reg local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_3;
 reg local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_4;
 reg local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_5;
 reg local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_stall_in_6;
wire local_bb4_c1_enter_c1_eni6_output_regs_ready;
 reg [223:0] local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG;
wire local_bb4_c1_enter_c1_eni6_input_accepted;
 reg local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG;
wire local_bb4_c1_exit_c1_exi2_entry_stall;
wire local_bb4_c1_exit_c1_exi2_output_regs_ready;
wire [69:0] local_bb4_c1_exit_c1_exi2_valid_bits;
wire local_bb4_c1_exit_c1_exi2_valid_in;
wire local_bb4_c1_exit_c1_exi2_phases;
wire local_bb4_c1_enter_c1_eni6_inc_pipelined_thread;
wire local_bb4_c1_enter_c1_eni6_dec_pipelined_thread;
wire local_bb4_c1_enter_c1_eni6_causedstall;

assign local_bb4_c1_enter_c1_eni6_inputs_ready = (local_bb4_c1_eni6_valid_out & local_bb4_c0_exe432_valid_out_1 & rcnode_175to176_rc0_t_322_0_valid_out_2_NO_SHIFT_REG);
assign local_bb4_c1_enter_c1_eni6_output_regs_ready = 1'b1;
assign local_bb4_c1_enter_c1_eni6_input_accepted = (local_bb4_c1_enter_c1_eni6_inputs_ready && !(local_bb4_c1_exit_c1_exi2_entry_stall));
assign local_bb4_c1_enter_c1_eni6_inc_pipelined_thread = rcnode_175to176_rc0_t_322_0_NO_SHIFT_REG[32];
assign local_bb4_c1_enter_c1_eni6_dec_pipelined_thread = ~(local_bb4_c0_exe432);
assign local_bb4_c1_eni6_stall_in = ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign local_bb4_c0_exe432_stall_in_1 = ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign rcnode_175to176_rc0_t_322_0_stall_in_2_NO_SHIFT_REG = ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) | ~(1'b1));
assign local_bb4_c1_enter_c1_eni6_causedstall = (1'b1 && ((~(local_bb4_c1_enter_c1_eni6_inputs_ready) | local_bb4_c1_exit_c1_exi2_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG <= local_bb4_c1_enter_c1_eni6_input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG <= 'x;
		local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c1_enter_c1_eni6_output_regs_ready)
		begin
			local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG <= local_bb4_c1_eni6;
			local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_0))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_1))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_2))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_3))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_4))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_5))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_c1_enter_c1_eni6_stall_in_6))
			begin
				local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene1_stall_local;
wire [31:0] local_bb4_c1_ene1;

assign local_bb4_c1_ene1 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[63:32];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene2_valid_out;
wire local_bb4_c1_ene2_stall_in;
wire local_bb4_c1_ene2_inputs_ready;
wire local_bb4_c1_ene2_stall_local;
wire [31:0] local_bb4_c1_ene2;

assign local_bb4_c1_ene2_inputs_ready = local_bb4_c1_enter_c1_eni6_valid_out_1_NO_SHIFT_REG;
assign local_bb4_c1_ene2 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[95:64];
assign local_bb4_c1_ene2_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_1 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene3_valid_out;
wire local_bb4_c1_ene3_stall_in;
wire local_bb4_c1_ene3_inputs_ready;
wire local_bb4_c1_ene3_stall_local;
wire [31:0] local_bb4_c1_ene3;

assign local_bb4_c1_ene3_inputs_ready = local_bb4_c1_enter_c1_eni6_valid_out_2_NO_SHIFT_REG;
assign local_bb4_c1_ene3 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[127:96];
assign local_bb4_c1_ene3_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_2 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene4_stall_local;
wire local_bb4_c1_ene4;

assign local_bb4_c1_ene4 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[128];

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene5_valid_out;
wire local_bb4_c1_ene5_stall_in;
wire local_bb4_c1_ene5_inputs_ready;
wire local_bb4_c1_ene5_stall_local;
wire [31:0] local_bb4_c1_ene5;

assign local_bb4_c1_ene5_inputs_ready = local_bb4_c1_enter_c1_eni6_valid_out_4_NO_SHIFT_REG;
assign local_bb4_c1_ene5 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[191:160];
assign local_bb4_c1_ene5_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_4 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene6_valid_out;
wire local_bb4_c1_ene6_stall_in;
wire local_bb4_c1_ene6_inputs_ready;
wire local_bb4_c1_ene6_stall_local;
wire local_bb4_c1_ene6;

assign local_bb4_c1_ene6_inputs_ready = local_bb4_c1_enter_c1_eni6_valid_out_5_NO_SHIFT_REG;
assign local_bb4_c1_ene6 = local_bb4_c1_enter_c1_eni6_NO_SHIFT_REG[192];
assign local_bb4_c1_ene6_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_5 = 1'b0;

// This section implements an unregistered operation.
// 
wire SFC_3_VALID_177_177_0_valid_out;
wire SFC_3_VALID_177_177_0_stall_in;
wire SFC_3_VALID_177_177_0_inputs_ready;
wire SFC_3_VALID_177_177_0_stall_local;
wire SFC_3_VALID_177_177_0;

assign SFC_3_VALID_177_177_0_inputs_ready = local_bb4_c1_enter_c1_eni6_valid_out_6_NO_SHIFT_REG;
assign SFC_3_VALID_177_177_0 = local_bb4_c1_enter_c1_eni6_valid_bit_NO_SHIFT_REG;
assign SFC_3_VALID_177_177_0_valid_out = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_6 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u34_stall_local;
wire [31:0] local_bb4_var__u34;

assign local_bb4_var__u34 = local_bb4_c1_ene1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_c1_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene2_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene2_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene2_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene2_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene2_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene2_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_c1_ene2_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_c1_ene2_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_c1_ene2_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_c1_ene2_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_c1_ene2_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene2),
	.data_out(rnode_177to178_bb4_c1_ene2_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_c1_ene2_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_c1_ene2_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_c1_ene2_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_c1_ene2_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_c1_ene2_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene2_stall_in = 1'b0;
assign rnode_177to178_bb4_c1_ene2_0_NO_SHIFT_REG = rnode_177to178_bb4_c1_ene2_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_c1_ene2_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_c1_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene3_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene3_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene3_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene3_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene3_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_c1_ene3_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_c1_ene3_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_c1_ene3_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_c1_ene3_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_c1_ene3_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene3),
	.data_out(rnode_177to178_bb4_c1_ene3_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_c1_ene3_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_c1_ene3_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_c1_ene3_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_c1_ene3_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_c1_ene3_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene3_stall_in = 1'b0;
assign rnode_177to178_bb4_c1_ene3_0_NO_SHIFT_REG = rnode_177to178_bb4_c1_ene3_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_c1_ene3_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__acl_ffwd_dest_f_7_stall_local;
wire [31:0] local_bb4__acl_ffwd_dest_f_7;

assign local_bb4__acl_ffwd_dest_f_7 = ffwd_7_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene5_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene5_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene5_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene5_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene5_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_c1_ene5_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_c1_ene5_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_c1_ene5_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_c1_ene5_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_c1_ene5_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene5),
	.data_out(rnode_177to178_bb4_c1_ene5_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_c1_ene5_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_c1_ene5_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_c1_ene5_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_c1_ene5_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_c1_ene5_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene5_stall_in = 1'b0;
assign rnode_177to178_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_177to178_bb4_c1_ene5_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_c1_ene5_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene6_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene6_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene6_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene6_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene6_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_c1_ene6_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_c1_ene6_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_c1_ene6_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_c1_ene6_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_c1_ene6_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene6),
	.data_out(rnode_177to178_bb4_c1_ene6_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_c1_ene6_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_c1_ene6_0_reg_178_fifo.DATA_WIDTH = 1;
defparam rnode_177to178_bb4_c1_ene6_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_c1_ene6_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_c1_ene6_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene6_stall_in = 1'b0;
assign rnode_177to178_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_177to178_bb4_c1_ene6_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_c1_ene6_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_177_178_0_inputs_ready;
 reg SFC_3_VALID_177_178_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_177_178_0_stall_in;
wire SFC_3_VALID_177_178_0_output_regs_ready;
 reg SFC_3_VALID_177_178_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_177_178_0_causedstall;

assign SFC_3_VALID_177_178_0_inputs_ready = 1'b1;
assign SFC_3_VALID_177_178_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_177_177_0_stall_in = 1'b0;
assign SFC_3_VALID_177_178_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_177_178_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_177_178_0_output_regs_ready)
		begin
			SFC_3_VALID_177_178_0_NO_SHIFT_REG <= SFC_3_VALID_177_177_0;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and2_i315_stall_local;
wire [31:0] local_bb4_and2_i315;

assign local_bb4_and2_i315 = (local_bb4_var__u34 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i320_stall_local;
wire [31:0] local_bb4_and12_i320;

assign local_bb4_and12_i320 = (local_bb4_var__u34 & 32'hFFFF);

// Register node:
//  * latency = 46
//  * capacity = 46
 logic rnode_178to224_bb4_c1_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to224_bb4_c1_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_178to224_bb4_c1_ene2_0_NO_SHIFT_REG;
 logic rnode_178to224_bb4_c1_ene2_0_reg_224_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to224_bb4_c1_ene2_0_reg_224_NO_SHIFT_REG;
 logic rnode_178to224_bb4_c1_ene2_0_valid_out_reg_224_NO_SHIFT_REG;
 logic rnode_178to224_bb4_c1_ene2_0_stall_in_reg_224_NO_SHIFT_REG;
 logic rnode_178to224_bb4_c1_ene2_0_stall_out_reg_224_NO_SHIFT_REG;

acl_data_fifo rnode_178to224_bb4_c1_ene2_0_reg_224_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to224_bb4_c1_ene2_0_reg_224_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to224_bb4_c1_ene2_0_stall_in_reg_224_NO_SHIFT_REG),
	.valid_out(rnode_178to224_bb4_c1_ene2_0_valid_out_reg_224_NO_SHIFT_REG),
	.stall_out(rnode_178to224_bb4_c1_ene2_0_stall_out_reg_224_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_c1_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_178to224_bb4_c1_ene2_0_reg_224_NO_SHIFT_REG)
);

defparam rnode_178to224_bb4_c1_ene2_0_reg_224_fifo.DEPTH = 46;
defparam rnode_178to224_bb4_c1_ene2_0_reg_224_fifo.DATA_WIDTH = 32;
defparam rnode_178to224_bb4_c1_ene2_0_reg_224_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to224_bb4_c1_ene2_0_reg_224_fifo.IMPL = "shift_reg";

assign rnode_178to224_bb4_c1_ene2_0_reg_224_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_c1_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to224_bb4_c1_ene2_0_NO_SHIFT_REG = rnode_178to224_bb4_c1_ene2_0_reg_224_NO_SHIFT_REG;
assign rnode_178to224_bb4_c1_ene2_0_stall_in_reg_224_NO_SHIFT_REG = 1'b0;
assign rnode_178to224_bb4_c1_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 56
//  * capacity = 56
 logic rnode_178to234_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to234_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_178to234_bb4_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_178to234_bb4_c1_ene3_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to234_bb4_c1_ene3_0_reg_234_NO_SHIFT_REG;
 logic rnode_178to234_bb4_c1_ene3_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_178to234_bb4_c1_ene3_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_178to234_bb4_c1_ene3_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_178to234_bb4_c1_ene3_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to234_bb4_c1_ene3_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to234_bb4_c1_ene3_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_178to234_bb4_c1_ene3_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_178to234_bb4_c1_ene3_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_c1_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_178to234_bb4_c1_ene3_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_178to234_bb4_c1_ene3_0_reg_234_fifo.DEPTH = 56;
defparam rnode_178to234_bb4_c1_ene3_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_178to234_bb4_c1_ene3_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to234_bb4_c1_ene3_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_178to234_bb4_c1_ene3_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to234_bb4_c1_ene3_0_NO_SHIFT_REG = rnode_178to234_bb4_c1_ene3_0_reg_234_NO_SHIFT_REG;
assign rnode_178to234_bb4_c1_ene3_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_178to234_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u35_stall_local;
wire [31:0] local_bb4_var__u35;

assign local_bb4_var__u35 = local_bb4__acl_ffwd_dest_f_7;

// Register node:
//  * latency = 51
//  * capacity = 51
 logic rnode_178to229_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_178to229_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene5_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to229_bb4_c1_ene5_0_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene5_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene5_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene5_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_178to229_bb4_c1_ene5_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to229_bb4_c1_ene5_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to229_bb4_c1_ene5_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_178to229_bb4_c1_ene5_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_178to229_bb4_c1_ene5_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_178to229_bb4_c1_ene5_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_178to229_bb4_c1_ene5_0_reg_229_fifo.DEPTH = 51;
defparam rnode_178to229_bb4_c1_ene5_0_reg_229_fifo.DATA_WIDTH = 32;
defparam rnode_178to229_bb4_c1_ene5_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to229_bb4_c1_ene5_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_178to229_bb4_c1_ene5_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to229_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_178to229_bb4_c1_ene5_0_reg_229_NO_SHIFT_REG;
assign rnode_178to229_bb4_c1_ene5_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_178to229_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 60
//  * capacity = 60
 logic rnode_178to238_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to238_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to238_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_178to238_bb4_c1_ene6_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to238_bb4_c1_ene6_0_reg_238_NO_SHIFT_REG;
 logic rnode_178to238_bb4_c1_ene6_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_178to238_bb4_c1_ene6_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_178to238_bb4_c1_ene6_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_178to238_bb4_c1_ene6_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to238_bb4_c1_ene6_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to238_bb4_c1_ene6_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_178to238_bb4_c1_ene6_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_178to238_bb4_c1_ene6_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_178to238_bb4_c1_ene6_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_178to238_bb4_c1_ene6_0_reg_238_fifo.DEPTH = 60;
defparam rnode_178to238_bb4_c1_ene6_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_178to238_bb4_c1_ene6_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to238_bb4_c1_ene6_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_178to238_bb4_c1_ene6_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to238_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_178to238_bb4_c1_ene6_0_reg_238_NO_SHIFT_REG;
assign rnode_178to238_bb4_c1_ene6_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_178to238_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_178_179_0_inputs_ready;
 reg SFC_3_VALID_178_179_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_178_179_0_stall_in;
wire SFC_3_VALID_178_179_0_output_regs_ready;
 reg SFC_3_VALID_178_179_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_178_179_0_causedstall;

assign SFC_3_VALID_178_179_0_inputs_ready = 1'b1;
assign SFC_3_VALID_178_179_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_177_178_0_stall_in = 1'b0;
assign SFC_3_VALID_178_179_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_178_179_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_178_179_0_output_regs_ready)
		begin
			SFC_3_VALID_178_179_0_NO_SHIFT_REG <= SFC_3_VALID_177_178_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i316_stall_local;
wire [31:0] local_bb4_shr3_i316;

assign local_bb4_shr3_i316 = ((local_bb4_and2_i315 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_224to225_bb4_c1_ene2_0_valid_out_NO_SHIFT_REG;
 logic rnode_224to225_bb4_c1_ene2_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_224to225_bb4_c1_ene2_0_NO_SHIFT_REG;
 logic rnode_224to225_bb4_c1_ene2_0_reg_225_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_224to225_bb4_c1_ene2_0_reg_225_NO_SHIFT_REG;
 logic rnode_224to225_bb4_c1_ene2_0_valid_out_reg_225_NO_SHIFT_REG;
 logic rnode_224to225_bb4_c1_ene2_0_stall_in_reg_225_NO_SHIFT_REG;
 logic rnode_224to225_bb4_c1_ene2_0_stall_out_reg_225_NO_SHIFT_REG;

acl_data_fifo rnode_224to225_bb4_c1_ene2_0_reg_225_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_224to225_bb4_c1_ene2_0_reg_225_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_224to225_bb4_c1_ene2_0_stall_in_reg_225_NO_SHIFT_REG),
	.valid_out(rnode_224to225_bb4_c1_ene2_0_valid_out_reg_225_NO_SHIFT_REG),
	.stall_out(rnode_224to225_bb4_c1_ene2_0_stall_out_reg_225_NO_SHIFT_REG),
	.data_in(rnode_178to224_bb4_c1_ene2_0_NO_SHIFT_REG),
	.data_out(rnode_224to225_bb4_c1_ene2_0_reg_225_NO_SHIFT_REG)
);

defparam rnode_224to225_bb4_c1_ene2_0_reg_225_fifo.DEPTH = 1;
defparam rnode_224to225_bb4_c1_ene2_0_reg_225_fifo.DATA_WIDTH = 32;
defparam rnode_224to225_bb4_c1_ene2_0_reg_225_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_224to225_bb4_c1_ene2_0_reg_225_fifo.IMPL = "shift_reg";

assign rnode_224to225_bb4_c1_ene2_0_reg_225_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to224_bb4_c1_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_224to225_bb4_c1_ene2_0_NO_SHIFT_REG = rnode_224to225_bb4_c1_ene2_0_reg_225_NO_SHIFT_REG;
assign rnode_224to225_bb4_c1_ene2_0_stall_in_reg_225_NO_SHIFT_REG = 1'b0;
assign rnode_224to225_bb4_c1_ene2_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene3_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_c1_ene3_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene3_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene3_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene3_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_c1_ene3_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_c1_ene3_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_c1_ene3_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_c1_ene3_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_c1_ene3_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(rnode_178to234_bb4_c1_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_234to235_bb4_c1_ene3_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_c1_ene3_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_c1_ene3_0_reg_235_fifo.DATA_WIDTH = 32;
defparam rnode_234to235_bb4_c1_ene3_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_c1_ene3_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_c1_ene3_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to234_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_c1_ene3_0_NO_SHIFT_REG = rnode_234to235_bb4_c1_ene3_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_c1_ene3_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i312_stall_local;
wire [31:0] local_bb4_xor_i312;

assign local_bb4_xor_i312 = (local_bb4_var__u35 ^ 32'h80000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene5_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_c1_ene5_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene5_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene5_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene5_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_c1_ene5_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_c1_ene5_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_c1_ene5_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_c1_ene5_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_c1_ene5_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(rnode_178to229_bb4_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_229to230_bb4_c1_ene5_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_c1_ene5_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_c1_ene5_0_reg_230_fifo.DATA_WIDTH = 32;
defparam rnode_229to230_bb4_c1_ene5_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_c1_ene5_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_c1_ene5_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to229_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_c1_ene5_0_NO_SHIFT_REG = rnode_229to230_bb4_c1_ene5_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_c1_ene5_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_c1_ene6_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_valid_out_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_stall_in_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_c1_ene6_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_c1_ene6_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_c1_ene6_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_c1_ene6_0_stall_in_0_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_c1_ene6_0_valid_out_0_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_c1_ene6_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in(rnode_178to238_bb4_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_238to239_bb4_c1_ene6_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_c1_ene6_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_c1_ene6_0_reg_239_fifo.DATA_WIDTH = 1;
defparam rnode_238to239_bb4_c1_ene6_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_c1_ene6_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_c1_ene6_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to238_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_c1_ene6_0_stall_in_0_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_c1_ene6_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_238to239_bb4_c1_ene6_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_c1_ene6_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_c1_ene6_1_NO_SHIFT_REG = rnode_238to239_bb4_c1_ene6_0_reg_239_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_179_180_0_inputs_ready;
 reg SFC_3_VALID_179_180_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_179_180_0_stall_in;
wire SFC_3_VALID_179_180_0_output_regs_ready;
 reg SFC_3_VALID_179_180_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_179_180_0_causedstall;

assign SFC_3_VALID_179_180_0_inputs_ready = 1'b1;
assign SFC_3_VALID_179_180_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_178_179_0_stall_in = 1'b0;
assign SFC_3_VALID_179_180_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_179_180_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_179_180_0_output_regs_ready)
		begin
			SFC_3_VALID_179_180_0_NO_SHIFT_REG <= SFC_3_VALID_178_179_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u36_stall_local;
wire [31:0] local_bb4_var__u36;

assign local_bb4_var__u36 = rnode_224to225_bb4_c1_ene2_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i313_stall_local;
wire [31:0] local_bb4_and_i313;

assign local_bb4_and_i313 = (local_bb4_xor_i312 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i319_stall_local;
wire [31:0] local_bb4_and10_i319;

assign local_bb4_and10_i319 = (local_bb4_xor_i312 & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_239to240_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_239to240_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_239to240_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_239to240_bb4_c1_ene6_0_reg_240_inputs_ready_NO_SHIFT_REG;
 logic rnode_239to240_bb4_c1_ene6_0_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_c1_ene6_0_valid_out_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_c1_ene6_0_stall_in_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_c1_ene6_0_stall_out_reg_240_NO_SHIFT_REG;

acl_data_fifo rnode_239to240_bb4_c1_ene6_0_reg_240_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to240_bb4_c1_ene6_0_reg_240_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to240_bb4_c1_ene6_0_stall_in_reg_240_NO_SHIFT_REG),
	.valid_out(rnode_239to240_bb4_c1_ene6_0_valid_out_reg_240_NO_SHIFT_REG),
	.stall_out(rnode_239to240_bb4_c1_ene6_0_stall_out_reg_240_NO_SHIFT_REG),
	.data_in(rnode_238to239_bb4_c1_ene6_1_NO_SHIFT_REG),
	.data_out(rnode_239to240_bb4_c1_ene6_0_reg_240_NO_SHIFT_REG)
);

defparam rnode_239to240_bb4_c1_ene6_0_reg_240_fifo.DEPTH = 1;
defparam rnode_239to240_bb4_c1_ene6_0_reg_240_fifo.DATA_WIDTH = 1;
defparam rnode_239to240_bb4_c1_ene6_0_reg_240_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to240_bb4_c1_ene6_0_reg_240_fifo.IMPL = "shift_reg";

assign rnode_239to240_bb4_c1_ene6_0_reg_240_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_c1_ene6_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_239to240_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_239to240_bb4_c1_ene6_0_reg_240_NO_SHIFT_REG;
assign rnode_239to240_bb4_c1_ene6_0_stall_in_reg_240_NO_SHIFT_REG = 1'b0;
assign rnode_239to240_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_180_181_0_inputs_ready;
 reg SFC_3_VALID_180_181_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_180_181_0_stall_in;
wire SFC_3_VALID_180_181_0_output_regs_ready;
 reg SFC_3_VALID_180_181_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_180_181_0_causedstall;

assign SFC_3_VALID_180_181_0_inputs_ready = 1'b1;
assign SFC_3_VALID_180_181_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_179_180_0_stall_in = 1'b0;
assign SFC_3_VALID_180_181_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_180_181_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_180_181_0_output_regs_ready)
		begin
			SFC_3_VALID_180_181_0_NO_SHIFT_REG <= SFC_3_VALID_179_180_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr_i220_stall_local;
wire [31:0] local_bb4_shr_i220;

assign local_bb4_shr_i220 = (local_bb4_var__u36 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and5_i226_stall_local;
wire [31:0] local_bb4_and5_i226;

assign local_bb4_and5_i226 = (local_bb4_var__u36 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i314_stall_local;
wire [31:0] local_bb4_shr_i314;

assign local_bb4_shr_i314 = ((local_bb4_and_i313 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i321_stall_local;
wire local_bb4_cmp13_i321;

assign local_bb4_cmp13_i321 = ((local_bb4_and10_i319 & 32'hFFFF) > (local_bb4_and12_i320 & 32'hFFFF));

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_240to243_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_240to243_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_240to243_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_240to243_bb4_c1_ene6_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic rnode_240to243_bb4_c1_ene6_0_reg_243_NO_SHIFT_REG;
 logic rnode_240to243_bb4_c1_ene6_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_240to243_bb4_c1_ene6_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_240to243_bb4_c1_ene6_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_240to243_bb4_c1_ene6_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to243_bb4_c1_ene6_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to243_bb4_c1_ene6_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_240to243_bb4_c1_ene6_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_240to243_bb4_c1_ene6_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(rnode_239to240_bb4_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_240to243_bb4_c1_ene6_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_240to243_bb4_c1_ene6_0_reg_243_fifo.DEPTH = 3;
defparam rnode_240to243_bb4_c1_ene6_0_reg_243_fifo.DATA_WIDTH = 1;
defparam rnode_240to243_bb4_c1_ene6_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to243_bb4_c1_ene6_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_240to243_bb4_c1_ene6_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_240to243_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_240to243_bb4_c1_ene6_0_reg_243_NO_SHIFT_REG;
assign rnode_240to243_bb4_c1_ene6_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_240to243_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_181_182_0_inputs_ready;
 reg SFC_3_VALID_181_182_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_181_182_0_stall_in;
wire SFC_3_VALID_181_182_0_output_regs_ready;
 reg SFC_3_VALID_181_182_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_181_182_0_causedstall;

assign SFC_3_VALID_181_182_0_inputs_ready = 1'b1;
assign SFC_3_VALID_181_182_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_180_181_0_stall_in = 1'b0;
assign SFC_3_VALID_181_182_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_181_182_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_181_182_0_output_regs_ready)
		begin
			SFC_3_VALID_181_182_0_NO_SHIFT_REG <= SFC_3_VALID_180_181_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and_i221_stall_local;
wire [31:0] local_bb4_and_i221;

assign local_bb4_and_i221 = ((local_bb4_shr_i220 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i232_stall_local;
wire local_bb4_lnot14_i232;

assign local_bb4_lnot14_i232 = ((local_bb4_and5_i226 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i254_stall_local;
wire [31:0] local_bb4_or_i254;

assign local_bb4_or_i254 = ((local_bb4_and5_i226 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i317_stall_local;
wire local_bb4_cmp_i317;

assign local_bb4_cmp_i317 = ((local_bb4_shr_i314 & 32'h7FFF) > (local_bb4_shr3_i316 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i318_stall_local;
wire local_bb4_cmp8_i318;

assign local_bb4_cmp8_i318 = ((local_bb4_shr_i314 & 32'h7FFF) == (local_bb4_shr3_i316 & 32'h7FFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_243to244_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_243to244_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG;
 logic rnode_243to244_bb4_c1_ene6_0_NO_SHIFT_REG;
 logic rnode_243to244_bb4_c1_ene6_0_reg_244_inputs_ready_NO_SHIFT_REG;
 logic rnode_243to244_bb4_c1_ene6_0_reg_244_NO_SHIFT_REG;
 logic rnode_243to244_bb4_c1_ene6_0_valid_out_reg_244_NO_SHIFT_REG;
 logic rnode_243to244_bb4_c1_ene6_0_stall_in_reg_244_NO_SHIFT_REG;
 logic rnode_243to244_bb4_c1_ene6_0_stall_out_reg_244_NO_SHIFT_REG;

acl_data_fifo rnode_243to244_bb4_c1_ene6_0_reg_244_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_243to244_bb4_c1_ene6_0_reg_244_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_243to244_bb4_c1_ene6_0_stall_in_reg_244_NO_SHIFT_REG),
	.valid_out(rnode_243to244_bb4_c1_ene6_0_valid_out_reg_244_NO_SHIFT_REG),
	.stall_out(rnode_243to244_bb4_c1_ene6_0_stall_out_reg_244_NO_SHIFT_REG),
	.data_in(rnode_240to243_bb4_c1_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_243to244_bb4_c1_ene6_0_reg_244_NO_SHIFT_REG)
);

defparam rnode_243to244_bb4_c1_ene6_0_reg_244_fifo.DEPTH = 1;
defparam rnode_243to244_bb4_c1_ene6_0_reg_244_fifo.DATA_WIDTH = 1;
defparam rnode_243to244_bb4_c1_ene6_0_reg_244_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_243to244_bb4_c1_ene6_0_reg_244_fifo.IMPL = "shift_reg";

assign rnode_243to244_bb4_c1_ene6_0_reg_244_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_240to243_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_243to244_bb4_c1_ene6_0_NO_SHIFT_REG = rnode_243to244_bb4_c1_ene6_0_reg_244_NO_SHIFT_REG;
assign rnode_243to244_bb4_c1_ene6_0_stall_in_reg_244_NO_SHIFT_REG = 1'b0;
assign rnode_243to244_bb4_c1_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_182_183_0_inputs_ready;
 reg SFC_3_VALID_182_183_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_182_183_0_stall_in;
wire SFC_3_VALID_182_183_0_output_regs_ready;
 reg SFC_3_VALID_182_183_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_182_183_0_causedstall;

assign SFC_3_VALID_182_183_0_inputs_ready = 1'b1;
assign SFC_3_VALID_182_183_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_181_182_0_stall_in = 1'b0;
assign SFC_3_VALID_182_183_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_182_183_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_182_183_0_output_regs_ready)
		begin
			SFC_3_VALID_182_183_0_NO_SHIFT_REG <= SFC_3_VALID_181_182_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i228_stall_local;
wire local_bb4_lnot_i228;

assign local_bb4_lnot_i228 = ((local_bb4_and_i221 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i230_stall_local;
wire local_bb4_cmp_i230;

assign local_bb4_cmp_i230 = ((local_bb4_and_i221 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_conv_i_i256_stall_local;
wire [63:0] local_bb4_conv_i_i256;

assign local_bb4_conv_i_i256[63:32] = 32'h0;
assign local_bb4_conv_i_i256[31:0] = ((local_bb4_or_i254 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4___i322_stall_local;
wire local_bb4___i322;

assign local_bb4___i322 = (local_bb4_cmp8_i318 & local_bb4_cmp13_i321);

// This section implements a registered operation.
// 
wire SFC_3_VALID_183_184_0_inputs_ready;
 reg SFC_3_VALID_183_184_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_183_184_0_stall_in;
wire SFC_3_VALID_183_184_0_output_regs_ready;
 reg SFC_3_VALID_183_184_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_183_184_0_causedstall;

assign SFC_3_VALID_183_184_0_inputs_ready = 1'b1;
assign SFC_3_VALID_183_184_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_182_183_0_stall_in = 1'b0;
assign SFC_3_VALID_183_184_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_183_184_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_183_184_0_output_regs_ready)
		begin
			SFC_3_VALID_183_184_0_NO_SHIFT_REG <= SFC_3_VALID_182_183_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_ene1_valid_out_1;
wire local_bb4_c1_ene1_stall_in_1;
wire local_bb4_var__u34_valid_out_2;
wire local_bb4_var__u34_stall_in_2;
wire local_bb4__21_i323_valid_out;
wire local_bb4__21_i323_stall_in;
wire local_bb4_c1_ene4_valid_out_1;
wire local_bb4_c1_ene4_stall_in_1;
wire local_bb4_xor_i312_valid_out_2;
wire local_bb4_xor_i312_stall_in_2;
wire local_bb4__21_i323_inputs_ready;
wire local_bb4__21_i323_stall_local;
wire local_bb4__21_i323;

assign local_bb4__21_i323_inputs_ready = (local_bb4_c1_enter_c1_eni6_valid_out_0_NO_SHIFT_REG & local_bb4_c1_enter_c1_eni6_valid_out_3_NO_SHIFT_REG);
assign local_bb4__21_i323 = (local_bb4_cmp_i317 | local_bb4___i322);
assign local_bb4_c1_ene1_valid_out_1 = 1'b1;
assign local_bb4_var__u34_valid_out_2 = 1'b1;
assign local_bb4__21_i323_valid_out = 1'b1;
assign local_bb4_c1_ene4_valid_out_1 = 1'b1;
assign local_bb4_xor_i312_valid_out_2 = 1'b1;
assign local_bb4_c1_enter_c1_eni6_stall_in_0 = 1'b0;
assign local_bb4_c1_enter_c1_eni6_stall_in_3 = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_184_185_0_inputs_ready;
 reg SFC_3_VALID_184_185_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_184_185_0_stall_in;
wire SFC_3_VALID_184_185_0_output_regs_ready;
 reg SFC_3_VALID_184_185_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_184_185_0_causedstall;

assign SFC_3_VALID_184_185_0_inputs_ready = 1'b1;
assign SFC_3_VALID_184_185_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_183_184_0_stall_in = 1'b0;
assign SFC_3_VALID_184_185_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_184_185_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_184_185_0_output_regs_ready)
		begin
			SFC_3_VALID_184_185_0_NO_SHIFT_REG <= SFC_3_VALID_183_184_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene1_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene1_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_c1_ene1_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene1_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene1_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene1_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_c1_ene1_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_c1_ene1_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_c1_ene1_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_c1_ene1_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_c1_ene1_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene1),
	.data_out(rnode_177to178_bb4_c1_ene1_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_c1_ene1_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_c1_ene1_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_c1_ene1_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_c1_ene1_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_c1_ene1_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene1_stall_in_1 = 1'b0;
assign rnode_177to178_bb4_c1_ene1_0_NO_SHIFT_REG = rnode_177to178_bb4_c1_ene1_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_c1_ene1_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_var__u34_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u34_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_var__u34_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u34_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u34_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_var__u34_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u34_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_var__u34_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u34_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u34_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_var__u34_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_var__u34_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_var__u34_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_var__u34_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_var__u34_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_var__u34_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_var__u34),
	.data_out(rnode_177to178_bb4_var__u34_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_var__u34_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_var__u34_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_var__u34_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_var__u34_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_var__u34_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u34_stall_in_2 = 1'b0;
assign rnode_177to178_bb4_var__u34_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_var__u34_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_var__u34_0_NO_SHIFT_REG = rnode_177to178_bb4_var__u34_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_var__u34_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_var__u34_1_NO_SHIFT_REG = rnode_177to178_bb4_var__u34_0_reg_178_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4__21_i323_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4__21_i323_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4__21_i323_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4__21_i323_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4__21_i323_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4__21_i323_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4__21_i323_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4__21_i323),
	.data_out(rnode_177to178_bb4__21_i323_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4__21_i323_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4__21_i323_0_reg_178_fifo.DATA_WIDTH = 1;
defparam rnode_177to178_bb4__21_i323_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4__21_i323_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4__21_i323_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i323_stall_in = 1'b0;
assign rnode_177to178_bb4__21_i323_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4__21_i323_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4__21_i323_0_NO_SHIFT_REG = rnode_177to178_bb4__21_i323_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4__21_i323_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4__21_i323_1_NO_SHIFT_REG = rnode_177to178_bb4__21_i323_0_reg_178_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene4_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene4_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene4_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene4_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_c1_ene4_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_c1_ene4_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_c1_ene4_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_c1_ene4_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_c1_ene4_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_c1_ene4_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_c1_ene4),
	.data_out(rnode_177to178_bb4_c1_ene4_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_c1_ene4_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_c1_ene4_0_reg_178_fifo.DATA_WIDTH = 1;
defparam rnode_177to178_bb4_c1_ene4_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_c1_ene4_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_c1_ene4_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_c1_ene4_stall_in_1 = 1'b0;
assign rnode_177to178_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_177to178_bb4_c1_ene4_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_c1_ene4_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb4_xor_i312_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i312_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_xor_i312_0_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i312_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i312_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_xor_i312_1_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i312_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb4_xor_i312_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i312_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i312_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb4_xor_i312_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb4_xor_i312_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb4_xor_i312_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb4_xor_i312_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb4_xor_i312_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb4_xor_i312_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i312),
	.data_out(rnode_177to178_bb4_xor_i312_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb4_xor_i312_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb4_xor_i312_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb4_xor_i312_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb4_xor_i312_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb4_xor_i312_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i312_stall_in_2 = 1'b0;
assign rnode_177to178_bb4_xor_i312_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_xor_i312_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_xor_i312_0_NO_SHIFT_REG = rnode_177to178_bb4_xor_i312_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb4_xor_i312_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_xor_i312_1_NO_SHIFT_REG = rnode_177to178_bb4_xor_i312_0_reg_178_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_185_186_0_inputs_ready;
 reg SFC_3_VALID_185_186_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_185_186_0_stall_in;
wire SFC_3_VALID_185_186_0_output_regs_ready;
 reg SFC_3_VALID_185_186_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_185_186_0_causedstall;

assign SFC_3_VALID_185_186_0_inputs_ready = 1'b1;
assign SFC_3_VALID_185_186_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_184_185_0_stall_in = 1'b0;
assign SFC_3_VALID_185_186_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_185_186_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_185_186_0_output_regs_ready)
		begin
			SFC_3_VALID_185_186_0_NO_SHIFT_REG <= SFC_3_VALID_184_185_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 51
//  * capacity = 51
 logic rnode_178to229_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_178to229_bb4_c1_ene1_0_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene1_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to229_bb4_c1_ene1_0_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene1_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene1_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene1_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_178to229_bb4_c1_ene1_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to229_bb4_c1_ene1_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to229_bb4_c1_ene1_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_178to229_bb4_c1_ene1_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_178to229_bb4_c1_ene1_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_c1_ene1_0_NO_SHIFT_REG),
	.data_out(rnode_178to229_bb4_c1_ene1_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_178to229_bb4_c1_ene1_0_reg_229_fifo.DEPTH = 51;
defparam rnode_178to229_bb4_c1_ene1_0_reg_229_fifo.DATA_WIDTH = 32;
defparam rnode_178to229_bb4_c1_ene1_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to229_bb4_c1_ene1_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_178to229_bb4_c1_ene1_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to229_bb4_c1_ene1_0_NO_SHIFT_REG = rnode_178to229_bb4_c1_ene1_0_reg_229_NO_SHIFT_REG;
assign rnode_178to229_bb4_c1_ene1_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_178to229_bb4_c1_ene1_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 51
//  * capacity = 51
 logic rnode_178to229_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene4_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene4_0_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene4_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene4_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_178to229_bb4_c1_ene4_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_178to229_bb4_c1_ene4_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to229_bb4_c1_ene4_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to229_bb4_c1_ene4_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_178to229_bb4_c1_ene4_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_178to229_bb4_c1_ene4_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb4_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_178to229_bb4_c1_ene4_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_178to229_bb4_c1_ene4_0_reg_229_fifo.DEPTH = 51;
defparam rnode_178to229_bb4_c1_ene4_0_reg_229_fifo.DATA_WIDTH = 1;
defparam rnode_178to229_bb4_c1_ene4_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to229_bb4_c1_ene4_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_178to229_bb4_c1_ene4_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to229_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_178to229_bb4_c1_ene4_0_reg_229_NO_SHIFT_REG;
assign rnode_178to229_bb4_c1_ene4_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_178to229_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__22_i324_stall_local;
wire [31:0] local_bb4__22_i324;

assign local_bb4__22_i324 = (rnode_177to178_bb4__21_i323_0_NO_SHIFT_REG ? rnode_177to178_bb4_var__u34_0_NO_SHIFT_REG : rnode_177to178_bb4_xor_i312_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i325_stall_local;
wire [31:0] local_bb4__23_i325;

assign local_bb4__23_i325 = (rnode_177to178_bb4__21_i323_1_NO_SHIFT_REG ? rnode_177to178_bb4_xor_i312_1_NO_SHIFT_REG : rnode_177to178_bb4_var__u34_1_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_3_VALID_186_187_0_inputs_ready;
 reg SFC_3_VALID_186_187_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_186_187_0_stall_in;
wire SFC_3_VALID_186_187_0_output_regs_ready;
 reg SFC_3_VALID_186_187_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_186_187_0_causedstall;

assign SFC_3_VALID_186_187_0_inputs_ready = 1'b1;
assign SFC_3_VALID_186_187_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_185_186_0_stall_in = 1'b0;
assign SFC_3_VALID_186_187_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_186_187_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_186_187_0_output_regs_ready)
		begin
			SFC_3_VALID_186_187_0_NO_SHIFT_REG <= SFC_3_VALID_185_186_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_c1_ene1_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene1_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_c1_ene1_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene1_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene1_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_c1_ene1_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene1_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_c1_ene1_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene1_0_valid_out_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene1_0_stall_in_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene1_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_c1_ene1_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_c1_ene1_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_c1_ene1_0_stall_in_0_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_c1_ene1_0_valid_out_0_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_c1_ene1_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(rnode_178to229_bb4_c1_ene1_0_NO_SHIFT_REG),
	.data_out(rnode_229to230_bb4_c1_ene1_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_c1_ene1_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_c1_ene1_0_reg_230_fifo.DATA_WIDTH = 32;
defparam rnode_229to230_bb4_c1_ene1_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_c1_ene1_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_c1_ene1_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to229_bb4_c1_ene1_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_c1_ene1_0_stall_in_0_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_c1_ene1_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_229to230_bb4_c1_ene1_0_NO_SHIFT_REG = rnode_229to230_bb4_c1_ene1_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_c1_ene1_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_229to230_bb4_c1_ene1_1_NO_SHIFT_REG = rnode_229to230_bb4_c1_ene1_0_reg_230_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_c1_ene4_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_valid_out_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_stall_in_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_c1_ene4_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_c1_ene4_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_c1_ene4_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_c1_ene4_0_stall_in_0_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_c1_ene4_0_valid_out_0_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_c1_ene4_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(rnode_178to229_bb4_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_229to230_bb4_c1_ene4_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_c1_ene4_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_c1_ene4_0_reg_230_fifo.DATA_WIDTH = 1;
defparam rnode_229to230_bb4_c1_ene4_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_c1_ene4_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_c1_ene4_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to229_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_c1_ene4_0_stall_in_0_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_c1_ene4_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_229to230_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_229to230_bb4_c1_ene4_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_c1_ene4_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_229to230_bb4_c1_ene4_1_NO_SHIFT_REG = rnode_229to230_bb4_c1_ene4_0_reg_230_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i328_stall_local;
wire [31:0] local_bb4_shr18_i328;

assign local_bb4_shr18_i328 = (local_bb4__22_i324 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i326_stall_local;
wire [31:0] local_bb4_shr16_i326;

assign local_bb4_shr16_i326 = (local_bb4__23_i325 >> 32'h17);

// This section implements a registered operation.
// 
wire SFC_3_VALID_187_188_0_inputs_ready;
 reg SFC_3_VALID_187_188_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_187_188_0_stall_in;
wire SFC_3_VALID_187_188_0_output_regs_ready;
 reg SFC_3_VALID_187_188_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_187_188_0_causedstall;

assign SFC_3_VALID_187_188_0_inputs_ready = 1'b1;
assign SFC_3_VALID_187_188_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_186_187_0_stall_in = 1'b0;
assign SFC_3_VALID_187_188_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_187_188_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_187_188_0_output_regs_ready)
		begin
			SFC_3_VALID_187_188_0_NO_SHIFT_REG <= SFC_3_VALID_186_187_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_cmp34_inputs_ready;
 reg local_bb4_cmp34_valid_out_NO_SHIFT_REG;
wire local_bb4_cmp34_stall_in;
wire local_bb4_cmp34_output_regs_ready;
wire local_bb4_cmp34;
 reg local_bb4_cmp34_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_cmp34_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_cmp34_causedstall;

acl_fp_cmp fp_module_local_bb4_cmp34 (
	.clock(clock),
	.dataa(rnode_229to230_bb4_c1_ene1_0_NO_SHIFT_REG),
	.datab(32'h0),
	.enable(local_bb4_cmp34_output_regs_ready),
	.result(local_bb4_cmp34)
);

defparam fp_module_local_bb4_cmp34.COMPARISON_MODE = 3;

assign local_bb4_cmp34_inputs_ready = 1'b1;
assign local_bb4_cmp34_output_regs_ready = 1'b1;
assign rnode_229to230_bb4_c1_ene1_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb4_cmp34_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_cmp34_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_cmp34_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_cmp34_output_regs_ready)
		begin
			local_bb4_cmp34_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_cmp34_valid_pipe_1_NO_SHIFT_REG <= local_bb4_cmp34_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_cmp34_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_cmp34_output_regs_ready)
		begin
			local_bb4_cmp34_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_cmp34_stall_in))
			begin
				local_bb4_cmp34_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u37_stall_local;
wire [31:0] local_bb4_var__u37;

assign local_bb4_var__u37 = rnode_229to230_bb4_c1_ene1_1_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_230to231_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_230to231_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_c1_ene4_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic rnode_230to231_bb4_c1_ene4_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_c1_ene4_0_valid_out_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_c1_ene4_0_stall_in_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_c1_ene4_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_c1_ene4_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_c1_ene4_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_c1_ene4_0_stall_in_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_c1_ene4_0_valid_out_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_c1_ene4_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in(rnode_229to230_bb4_c1_ene4_1_NO_SHIFT_REG),
	.data_out(rnode_230to231_bb4_c1_ene4_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_c1_ene4_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_c1_ene4_0_reg_231_fifo.DATA_WIDTH = 1;
defparam rnode_230to231_bb4_c1_ene4_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_c1_ene4_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_c1_ene4_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_229to230_bb4_c1_ene4_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_230to231_bb4_c1_ene4_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_c1_ene4_0_stall_in_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i329_stall_local;
wire [31:0] local_bb4_and19_i329;

assign local_bb4_and19_i329 = ((local_bb4_shr18_i328 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i354_stall_local;
wire [31:0] local_bb4_sub_i354;

assign local_bb4_sub_i354 = ((local_bb4_shr16_i326 & 32'h1FF) - (local_bb4_shr18_i328 & 32'h1FF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_188_189_0_inputs_ready;
 reg SFC_3_VALID_188_189_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_188_189_0_stall_in;
wire SFC_3_VALID_188_189_0_output_regs_ready;
 reg SFC_3_VALID_188_189_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_188_189_0_causedstall;

assign SFC_3_VALID_188_189_0_inputs_ready = 1'b1;
assign SFC_3_VALID_188_189_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_187_188_0_stall_in = 1'b0;
assign SFC_3_VALID_188_189_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_188_189_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_188_189_0_output_regs_ready)
		begin
			SFC_3_VALID_188_189_0_NO_SHIFT_REG <= SFC_3_VALID_187_188_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_cmp34_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp34_0_stall_in_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp34_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp34_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp34_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp34_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp34_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp34_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_cmp34_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_cmp34_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_cmp34_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_cmp34_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_cmp34_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(local_bb4_cmp34),
	.data_out(rnode_233to234_bb4_cmp34_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_cmp34_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_cmp34_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_233to234_bb4_cmp34_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_cmp34_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_cmp34_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp34_stall_in = 1'b0;
assign rnode_233to234_bb4_cmp34_0_NO_SHIFT_REG = rnode_233to234_bb4_cmp34_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_cmp34_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_cmp34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i_stall_local;
wire [31:0] local_bb4_shr2_i;

assign local_bb4_shr2_i = (local_bb4_var__u37 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and6_i_stall_local;
wire [31:0] local_bb4_and6_i;

assign local_bb4_and6_i = (local_bb4_var__u37 & 32'h7FFFFF);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_231to234_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_231to234_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_231to234_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_231to234_bb4_c1_ene4_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_231to234_bb4_c1_ene4_0_reg_234_NO_SHIFT_REG;
 logic rnode_231to234_bb4_c1_ene4_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_231to234_bb4_c1_ene4_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_231to234_bb4_c1_ene4_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_231to234_bb4_c1_ene4_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to234_bb4_c1_ene4_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to234_bb4_c1_ene4_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_231to234_bb4_c1_ene4_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_231to234_bb4_c1_ene4_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(rnode_230to231_bb4_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_231to234_bb4_c1_ene4_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_231to234_bb4_c1_ene4_0_reg_234_fifo.DEPTH = 3;
defparam rnode_231to234_bb4_c1_ene4_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_231to234_bb4_c1_ene4_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to234_bb4_c1_ene4_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_231to234_bb4_c1_ene4_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_231to234_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_231to234_bb4_c1_ene4_0_reg_234_NO_SHIFT_REG;
assign rnode_231to234_bb4_c1_ene4_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_231to234_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i333_stall_local;
wire local_bb4_lnot23_i333;

assign local_bb4_lnot23_i333 = ((local_bb4_and19_i329 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i335_stall_local;
wire local_bb4_cmp27_i335;

assign local_bb4_cmp27_i335 = ((local_bb4_and19_i329 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and69_i_stall_local;
wire [31:0] local_bb4_and69_i;

assign local_bb4_and69_i = (local_bb4_sub_i354 & 32'hFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_189_190_0_inputs_ready;
 reg SFC_3_VALID_189_190_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_189_190_0_stall_in;
wire SFC_3_VALID_189_190_0_output_regs_ready;
 reg SFC_3_VALID_189_190_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_189_190_0_causedstall;

assign SFC_3_VALID_189_190_0_inputs_ready = 1'b1;
assign SFC_3_VALID_189_190_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_188_189_0_stall_in = 1'b0;
assign SFC_3_VALID_189_190_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_189_190_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_189_190_0_output_regs_ready)
		begin
			SFC_3_VALID_189_190_0_NO_SHIFT_REG <= SFC_3_VALID_188_189_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_234to237_bb4_cmp34_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to237_bb4_cmp34_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to237_bb4_cmp34_0_NO_SHIFT_REG;
 logic rnode_234to237_bb4_cmp34_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to237_bb4_cmp34_0_reg_237_NO_SHIFT_REG;
 logic rnode_234to237_bb4_cmp34_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_234to237_bb4_cmp34_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_234to237_bb4_cmp34_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_234to237_bb4_cmp34_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to237_bb4_cmp34_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to237_bb4_cmp34_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_234to237_bb4_cmp34_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_234to237_bb4_cmp34_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(rnode_233to234_bb4_cmp34_0_NO_SHIFT_REG),
	.data_out(rnode_234to237_bb4_cmp34_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_234to237_bb4_cmp34_0_reg_237_fifo.DEPTH = 3;
defparam rnode_234to237_bb4_cmp34_0_reg_237_fifo.DATA_WIDTH = 1;
defparam rnode_234to237_bb4_cmp34_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to237_bb4_cmp34_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_234to237_bb4_cmp34_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4_cmp34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to237_bb4_cmp34_0_NO_SHIFT_REG = rnode_234to237_bb4_cmp34_0_reg_237_NO_SHIFT_REG;
assign rnode_234to237_bb4_cmp34_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_234to237_bb4_cmp34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or47_i_stall_local;
wire [31:0] local_bb4_or47_i;

assign local_bb4_or47_i = ((local_bb4_and6_i & 32'h7FFFFF) | 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene4_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene4_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene4_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene4_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene4_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_c1_ene4_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_c1_ene4_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_c1_ene4_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_c1_ene4_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_c1_ene4_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_c1_ene4_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(rnode_231to234_bb4_c1_ene4_0_NO_SHIFT_REG),
	.data_out(rnode_234to235_bb4_c1_ene4_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_c1_ene4_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_c1_ene4_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4_c1_ene4_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_c1_ene4_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_c1_ene4_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_231to234_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_c1_ene4_0_NO_SHIFT_REG = rnode_234to235_bb4_c1_ene4_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_c1_ene4_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp70_i_stall_local;
wire local_bb4_cmp70_i;

assign local_bb4_cmp70_i = ((local_bb4_and69_i & 32'hFF) > 32'h1F);

// This section implements a registered operation.
// 
wire SFC_3_VALID_190_191_0_inputs_ready;
 reg SFC_3_VALID_190_191_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_190_191_0_stall_in;
wire SFC_3_VALID_190_191_0_output_regs_ready;
 reg SFC_3_VALID_190_191_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_190_191_0_causedstall;

assign SFC_3_VALID_190_191_0_inputs_ready = 1'b1;
assign SFC_3_VALID_190_191_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_189_190_0_stall_in = 1'b0;
assign SFC_3_VALID_190_191_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_190_191_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_190_191_0_output_regs_ready)
		begin
			SFC_3_VALID_190_191_0_NO_SHIFT_REG <= SFC_3_VALID_189_190_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_cmp34_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_valid_out_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_stall_in_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp34_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_cmp34_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_cmp34_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_cmp34_0_stall_in_0_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_cmp34_0_valid_out_0_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_cmp34_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(rnode_234to237_bb4_cmp34_0_NO_SHIFT_REG),
	.data_out(rnode_237to238_bb4_cmp34_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_cmp34_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_cmp34_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_237to238_bb4_cmp34_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_cmp34_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_cmp34_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_234to237_bb4_cmp34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_cmp34_0_stall_in_0_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_cmp34_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_cmp34_0_NO_SHIFT_REG = rnode_237to238_bb4_cmp34_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_cmp34_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_cmp34_1_NO_SHIFT_REG = rnode_237to238_bb4_cmp34_0_reg_238_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv1_i_i_stall_local;
wire [63:0] local_bb4_conv1_i_i;

assign local_bb4_conv1_i_i[63:32] = 32'h0;
assign local_bb4_conv1_i_i[31:0] = ((local_bb4_or47_i & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i324_valid_out_1;
wire local_bb4__22_i324_stall_in_1;
wire local_bb4__23_i325_valid_out_1;
wire local_bb4__23_i325_stall_in_1;
wire local_bb4_shr16_i326_valid_out_1;
wire local_bb4_shr16_i326_stall_in_1;
wire local_bb4_lnot23_i333_valid_out;
wire local_bb4_lnot23_i333_stall_in;
wire local_bb4_cmp27_i335_valid_out;
wire local_bb4_cmp27_i335_stall_in;
wire local_bb4_align_0_i355_valid_out;
wire local_bb4_align_0_i355_stall_in;
wire local_bb4_align_0_i355_inputs_ready;
wire local_bb4_align_0_i355_stall_local;
wire [31:0] local_bb4_align_0_i355;

assign local_bb4_align_0_i355_inputs_ready = (rnode_177to178_bb4__21_i323_0_valid_out_0_NO_SHIFT_REG & rnode_177to178_bb4_var__u34_0_valid_out_0_NO_SHIFT_REG & rnode_177to178_bb4_xor_i312_0_valid_out_0_NO_SHIFT_REG & rnode_177to178_bb4__21_i323_0_valid_out_1_NO_SHIFT_REG & rnode_177to178_bb4_xor_i312_0_valid_out_1_NO_SHIFT_REG & rnode_177to178_bb4_var__u34_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_align_0_i355 = (local_bb4_cmp70_i ? 32'h1F : (local_bb4_and69_i & 32'hFF));
assign local_bb4__22_i324_valid_out_1 = 1'b1;
assign local_bb4__23_i325_valid_out_1 = 1'b1;
assign local_bb4_shr16_i326_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i333_valid_out = 1'b1;
assign local_bb4_cmp27_i335_valid_out = 1'b1;
assign local_bb4_align_0_i355_valid_out = 1'b1;
assign rnode_177to178_bb4__21_i323_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_var__u34_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_xor_i312_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4__21_i323_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_xor_i312_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb4_var__u34_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_191_192_0_inputs_ready;
 reg SFC_3_VALID_191_192_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_191_192_0_stall_in;
wire SFC_3_VALID_191_192_0_output_regs_ready;
 reg SFC_3_VALID_191_192_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_191_192_0_causedstall;

assign SFC_3_VALID_191_192_0_inputs_ready = 1'b1;
assign SFC_3_VALID_191_192_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_190_191_0_stall_in = 1'b0;
assign SFC_3_VALID_191_192_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_191_192_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_191_192_0_output_regs_ready)
		begin
			SFC_3_VALID_191_192_0_NO_SHIFT_REG <= SFC_3_VALID_190_191_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_cmp34_0_valid_out_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp34_0_stall_in_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp34_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp34_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp34_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp34_0_valid_out_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp34_0_stall_in_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp34_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_cmp34_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_cmp34_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_cmp34_0_stall_in_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_cmp34_0_valid_out_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_cmp34_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in(rnode_237to238_bb4_cmp34_1_NO_SHIFT_REG),
	.data_out(rnode_238to239_bb4_cmp34_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_cmp34_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_cmp34_0_reg_239_fifo.DATA_WIDTH = 1;
defparam rnode_238to239_bb4_cmp34_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_cmp34_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_cmp34_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_cmp34_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_cmp34_0_NO_SHIFT_REG = rnode_238to239_bb4_cmp34_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_cmp34_0_stall_in_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_cmp34_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4__22_i324_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i324_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__22_i324_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i324_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i324_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__22_i324_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i324_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__22_i324_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i324_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i324_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__22_i324_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4__22_i324_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4__22_i324_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4__22_i324_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4__22_i324_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4__22_i324_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4__22_i324),
	.data_out(rnode_178to179_bb4__22_i324_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4__22_i324_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4__22_i324_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb4__22_i324_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4__22_i324_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4__22_i324_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i324_stall_in_1 = 1'b0;
assign rnode_178to179_bb4__22_i324_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__22_i324_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__22_i324_0_NO_SHIFT_REG = rnode_178to179_bb4__22_i324_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4__22_i324_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__22_i324_1_NO_SHIFT_REG = rnode_178to179_bb4__22_i324_0_reg_179_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4__23_i325_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i325_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i325_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i325_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4__23_i325_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4__23_i325_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4__23_i325_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4__23_i325_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4__23_i325_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4__23_i325_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4__23_i325_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4__23_i325),
	.data_out(rnode_178to179_bb4__23_i325_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4__23_i325_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4__23_i325_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb4__23_i325_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4__23_i325_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4__23_i325_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i325_stall_in_1 = 1'b0;
assign rnode_178to179_bb4__23_i325_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__23_i325_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__23_i325_0_NO_SHIFT_REG = rnode_178to179_bb4__23_i325_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4__23_i325_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__23_i325_1_NO_SHIFT_REG = rnode_178to179_bb4__23_i325_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4__23_i325_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4__23_i325_2_NO_SHIFT_REG = rnode_178to179_bb4__23_i325_0_reg_179_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_178to180_bb4_shr16_i326_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i326_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to180_bb4_shr16_i326_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i326_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i326_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to180_bb4_shr16_i326_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i326_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to180_bb4_shr16_i326_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i326_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i326_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_shr16_i326_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_178to180_bb4_shr16_i326_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to180_bb4_shr16_i326_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to180_bb4_shr16_i326_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_178to180_bb4_shr16_i326_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_178to180_bb4_shr16_i326_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i326 & 32'h1FF)),
	.data_out(rnode_178to180_bb4_shr16_i326_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_178to180_bb4_shr16_i326_0_reg_180_fifo.DEPTH = 2;
defparam rnode_178to180_bb4_shr16_i326_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_178to180_bb4_shr16_i326_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to180_bb4_shr16_i326_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_178to180_bb4_shr16_i326_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i326_stall_in_1 = 1'b0;
assign rnode_178to180_bb4_shr16_i326_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_shr16_i326_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_shr16_i326_0_NO_SHIFT_REG = rnode_178to180_bb4_shr16_i326_0_reg_180_NO_SHIFT_REG;
assign rnode_178to180_bb4_shr16_i326_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_shr16_i326_1_NO_SHIFT_REG = rnode_178to180_bb4_shr16_i326_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_lnot23_i333_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i333_0_stall_in_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i333_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i333_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i333_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i333_0_valid_out_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i333_0_stall_in_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_lnot23_i333_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_lnot23_i333_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_lnot23_i333_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_lnot23_i333_0_stall_in_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_lnot23_i333_0_valid_out_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_lnot23_i333_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i333),
	.data_out(rnode_178to179_bb4_lnot23_i333_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_lnot23_i333_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4_lnot23_i333_0_reg_179_fifo.DATA_WIDTH = 1;
defparam rnode_178to179_bb4_lnot23_i333_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4_lnot23_i333_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4_lnot23_i333_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i333_stall_in = 1'b0;
assign rnode_178to179_bb4_lnot23_i333_0_NO_SHIFT_REG = rnode_178to179_bb4_lnot23_i333_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_lnot23_i333_0_stall_in_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_lnot23_i333_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_178to180_bb4_cmp27_i335_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_1_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_2_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_178to180_bb4_cmp27_i335_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_178to180_bb4_cmp27_i335_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to180_bb4_cmp27_i335_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to180_bb4_cmp27_i335_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_178to180_bb4_cmp27_i335_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_178to180_bb4_cmp27_i335_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i335),
	.data_out(rnode_178to180_bb4_cmp27_i335_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_178to180_bb4_cmp27_i335_0_reg_180_fifo.DEPTH = 2;
defparam rnode_178to180_bb4_cmp27_i335_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_178to180_bb4_cmp27_i335_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to180_bb4_cmp27_i335_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_178to180_bb4_cmp27_i335_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i335_stall_in = 1'b0;
assign rnode_178to180_bb4_cmp27_i335_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i335_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_cmp27_i335_0_NO_SHIFT_REG = rnode_178to180_bb4_cmp27_i335_0_reg_180_NO_SHIFT_REG;
assign rnode_178to180_bb4_cmp27_i335_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_cmp27_i335_1_NO_SHIFT_REG = rnode_178to180_bb4_cmp27_i335_0_reg_180_NO_SHIFT_REG;
assign rnode_178to180_bb4_cmp27_i335_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_cmp27_i335_2_NO_SHIFT_REG = rnode_178to180_bb4_cmp27_i335_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb4_align_0_i355_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i355_0_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i355_1_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i355_2_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i355_3_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i355_4_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb4_align_0_i355_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb4_align_0_i355_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb4_align_0_i355_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb4_align_0_i355_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb4_align_0_i355_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb4_align_0_i355_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb4_align_0_i355_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in((local_bb4_align_0_i355 & 32'hFF)),
	.data_out(rnode_178to179_bb4_align_0_i355_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb4_align_0_i355_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb4_align_0_i355_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb4_align_0_i355_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb4_align_0_i355_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb4_align_0_i355_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_align_0_i355_stall_in = 1'b0;
assign rnode_178to179_bb4_align_0_i355_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i355_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i355_0_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i355_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i355_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i355_1_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i355_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i355_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i355_2_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i355_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i355_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i355_3_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i355_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb4_align_0_i355_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb4_align_0_i355_4_NO_SHIFT_REG = rnode_178to179_bb4_align_0_i355_0_reg_179_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_192_193_0_inputs_ready;
 reg SFC_3_VALID_192_193_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_192_193_0_stall_in;
wire SFC_3_VALID_192_193_0_output_regs_ready;
 reg SFC_3_VALID_192_193_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_192_193_0_causedstall;

assign SFC_3_VALID_192_193_0_inputs_ready = 1'b1;
assign SFC_3_VALID_192_193_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_191_192_0_stall_in = 1'b0;
assign SFC_3_VALID_192_193_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_192_193_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_192_193_0_output_regs_ready)
		begin
			SFC_3_VALID_192_193_0_NO_SHIFT_REG <= SFC_3_VALID_191_192_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_239to242_bb4_cmp34_0_valid_out_NO_SHIFT_REG;
 logic rnode_239to242_bb4_cmp34_0_stall_in_NO_SHIFT_REG;
 logic rnode_239to242_bb4_cmp34_0_NO_SHIFT_REG;
 logic rnode_239to242_bb4_cmp34_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic rnode_239to242_bb4_cmp34_0_reg_242_NO_SHIFT_REG;
 logic rnode_239to242_bb4_cmp34_0_valid_out_reg_242_NO_SHIFT_REG;
 logic rnode_239to242_bb4_cmp34_0_stall_in_reg_242_NO_SHIFT_REG;
 logic rnode_239to242_bb4_cmp34_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_239to242_bb4_cmp34_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to242_bb4_cmp34_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to242_bb4_cmp34_0_stall_in_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_239to242_bb4_cmp34_0_valid_out_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_239to242_bb4_cmp34_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in(rnode_238to239_bb4_cmp34_0_NO_SHIFT_REG),
	.data_out(rnode_239to242_bb4_cmp34_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_239to242_bb4_cmp34_0_reg_242_fifo.DEPTH = 3;
defparam rnode_239to242_bb4_cmp34_0_reg_242_fifo.DATA_WIDTH = 1;
defparam rnode_239to242_bb4_cmp34_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to242_bb4_cmp34_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_239to242_bb4_cmp34_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_cmp34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_239to242_bb4_cmp34_0_NO_SHIFT_REG = rnode_239to242_bb4_cmp34_0_reg_242_NO_SHIFT_REG;
assign rnode_239to242_bb4_cmp34_0_stall_in_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_239to242_bb4_cmp34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i331_stall_local;
wire [31:0] local_bb4_and21_i331;

assign local_bb4_and21_i331 = (rnode_178to179_bb4__22_i324_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i330_valid_out;
wire local_bb4_and20_i330_stall_in;
wire local_bb4_and20_i330_inputs_ready;
wire local_bb4_and20_i330_stall_local;
wire [31:0] local_bb4_and20_i330;

assign local_bb4_and20_i330_inputs_ready = rnode_178to179_bb4__23_i325_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i330 = (rnode_178to179_bb4__23_i325_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i330_valid_out = 1'b1;
assign rnode_178to179_bb4__23_i325_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i336_valid_out;
wire local_bb4_and35_i336_stall_in;
wire local_bb4_and35_i336_inputs_ready;
wire local_bb4_and35_i336_stall_local;
wire [31:0] local_bb4_and35_i336;

assign local_bb4_and35_i336_inputs_ready = rnode_178to179_bb4__23_i325_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i336 = (rnode_178to179_bb4__23_i325_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i336_valid_out = 1'b1;
assign rnode_178to179_bb4__23_i325_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor36_i_stall_local;
wire [31:0] local_bb4_xor36_i;

assign local_bb4_xor36_i = (rnode_178to179_bb4__23_i325_2_NO_SHIFT_REG ^ rnode_178to179_bb4__22_i324_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i327_stall_local;
wire [31:0] local_bb4_and17_i327;

assign local_bb4_and17_i327 = ((rnode_178to180_bb4_shr16_i326_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_shr16_i326_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i326_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i326_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i326_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_shr16_i326_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i326_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i326_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_shr16_i326_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_shr16_i326_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_shr16_i326_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_shr16_i326_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_shr16_i326_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_shr16_i326_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((rnode_178to180_bb4_shr16_i326_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_180to182_bb4_shr16_i326_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_shr16_i326_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_shr16_i326_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_shr16_i326_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_shr16_i326_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_shr16_i326_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to180_bb4_shr16_i326_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_shr16_i326_0_NO_SHIFT_REG = rnode_180to182_bb4_shr16_i326_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_shr16_i326_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_shr16_i326_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and94_i_stall_local;
wire [31:0] local_bb4_and94_i;

assign local_bb4_and94_i = ((rnode_178to179_bb4_align_0_i355_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and96_i_stall_local;
wire [31:0] local_bb4_and96_i;

assign local_bb4_and96_i = ((rnode_178to179_bb4_align_0_i355_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and116_i_stall_local;
wire [31:0] local_bb4_and116_i;

assign local_bb4_and116_i = ((rnode_178to179_bb4_align_0_i355_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and131_i_stall_local;
wire [31:0] local_bb4_and131_i;

assign local_bb4_and131_i = ((rnode_178to179_bb4_align_0_i355_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and150_i_stall_local;
wire [31:0] local_bb4_and150_i;

assign local_bb4_and150_i = ((rnode_178to179_bb4_align_0_i355_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements a registered operation.
// 
wire SFC_3_VALID_193_194_0_inputs_ready;
 reg SFC_3_VALID_193_194_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_193_194_0_stall_in;
wire SFC_3_VALID_193_194_0_output_regs_ready;
 reg SFC_3_VALID_193_194_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_193_194_0_causedstall;

assign SFC_3_VALID_193_194_0_inputs_ready = 1'b1;
assign SFC_3_VALID_193_194_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_192_193_0_stall_in = 1'b0;
assign SFC_3_VALID_193_194_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_193_194_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_193_194_0_output_regs_ready)
		begin
			SFC_3_VALID_193_194_0_NO_SHIFT_REG <= SFC_3_VALID_192_193_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4_cmp34_0_valid_out_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp34_0_stall_in_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp34_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp34_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp34_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp34_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp34_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp34_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4_cmp34_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4_cmp34_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4_cmp34_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4_cmp34_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4_cmp34_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(rnode_239to242_bb4_cmp34_0_NO_SHIFT_REG),
	.data_out(rnode_242to243_bb4_cmp34_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4_cmp34_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4_cmp34_0_reg_243_fifo.DATA_WIDTH = 1;
defparam rnode_242to243_bb4_cmp34_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4_cmp34_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4_cmp34_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_239to242_bb4_cmp34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_cmp34_0_NO_SHIFT_REG = rnode_242to243_bb4_cmp34_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_cmp34_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_cmp34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i340_stall_local;
wire local_bb4_lnot33_not_i340;

assign local_bb4_lnot33_not_i340 = ((local_bb4_and21_i331 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or65_i_stall_local;
wire [31:0] local_bb4_or65_i;

assign local_bb4_or65_i = ((local_bb4_and21_i331 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_and20_i330_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i330_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and20_i330_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i330_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i330_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and20_i330_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i330_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and20_i330_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i330_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i330_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and20_i330_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_and20_i330_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_and20_i330_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_and20_i330_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_and20_i330_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_and20_i330_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i330 & 32'h7FFFFF)),
	.data_out(rnode_179to180_bb4_and20_i330_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_and20_i330_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_and20_i330_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_and20_i330_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_and20_i330_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_and20_i330_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i330_stall_in = 1'b0;
assign rnode_179to180_bb4_and20_i330_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and20_i330_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_and20_i330_0_NO_SHIFT_REG = rnode_179to180_bb4_and20_i330_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_and20_i330_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_and20_i330_1_NO_SHIFT_REG = rnode_179to180_bb4_and20_i330_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_and35_i336_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i336_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and35_i336_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i336_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and35_i336_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i336_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i336_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and35_i336_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_and35_i336_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_and35_i336_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_and35_i336_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_and35_i336_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_and35_i336_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i336 & 32'h80000000)),
	.data_out(rnode_179to180_bb4_and35_i336_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_and35_i336_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_and35_i336_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_and35_i336_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_and35_i336_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_and35_i336_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i336_stall_in = 1'b0;
assign rnode_179to180_bb4_and35_i336_0_NO_SHIFT_REG = rnode_179to180_bb4_and35_i336_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_and35_i336_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and35_i336_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp38_i_stall_local;
wire local_bb4_cmp38_i;

assign local_bb4_cmp38_i = ($signed(local_bb4_xor36_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor36_lobit_i_stall_local;
wire [31:0] local_bb4_xor36_lobit_i;

assign local_bb4_xor36_lobit_i = ($signed(local_bb4_xor36_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and37_lobit_i_stall_local;
wire [31:0] local_bb4_and37_lobit_i;

assign local_bb4_and37_lobit_i = (local_bb4_xor36_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i332_stall_local;
wire local_bb4_lnot_i332;

assign local_bb4_lnot_i332 = ((local_bb4_and17_i327 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i334_stall_local;
wire local_bb4_cmp25_i334;

assign local_bb4_cmp25_i334 = ((local_bb4_and17_i327 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp97_i_stall_local;
wire local_bb4_cmp97_i;

assign local_bb4_cmp97_i = ((local_bb4_and96_i & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp117_i_stall_local;
wire local_bb4_cmp117_i;

assign local_bb4_cmp117_i = ((local_bb4_and116_i & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp132_not_i_stall_local;
wire local_bb4_cmp132_not_i;

assign local_bb4_cmp132_not_i = ((local_bb4_and131_i & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i366_stall_local;
wire local_bb4_Pivot20_i366;

assign local_bb4_Pivot20_i366 = ((local_bb4_and150_i & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i367_stall_local;
wire local_bb4_SwitchLeaf_i367;

assign local_bb4_SwitchLeaf_i367 = ((local_bb4_and150_i & 32'h3) == 32'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_194_195_0_inputs_ready;
 reg SFC_3_VALID_194_195_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_194_195_0_stall_in;
wire SFC_3_VALID_194_195_0_output_regs_ready;
 reg SFC_3_VALID_194_195_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_194_195_0_causedstall;

assign SFC_3_VALID_194_195_0_inputs_ready = 1'b1;
assign SFC_3_VALID_194_195_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_193_194_0_stall_in = 1'b0;
assign SFC_3_VALID_194_195_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_194_195_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_194_195_0_output_regs_ready)
		begin
			SFC_3_VALID_194_195_0_NO_SHIFT_REG <= SFC_3_VALID_193_194_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shl66_i_stall_local;
wire [31:0] local_bb4_shl66_i;

assign local_bb4_shl66_i = ((local_bb4_or65_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i338_stall_local;
wire local_bb4_lnot30_i338;

assign local_bb4_lnot30_i338 = ((rnode_179to180_bb4_and20_i330_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i350_stall_local;
wire [31:0] local_bb4_or_i350;

assign local_bb4_or_i350 = ((rnode_179to180_bb4_and20_i330_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_and35_i336_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i336_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and35_i336_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i336_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and35_i336_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i336_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i336_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and35_i336_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_and35_i336_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_and35_i336_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_and35_i336_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_and35_i336_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_and35_i336_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((rnode_179to180_bb4_and35_i336_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_180to182_bb4_and35_i336_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_and35_i336_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_and35_i336_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_and35_i336_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_and35_i336_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_and35_i336_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_and35_i336_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and35_i336_0_NO_SHIFT_REG = rnode_180to182_bb4_and35_i336_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_and35_i336_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and35_i336_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i337_stall_local;
wire local_bb4_cmp25_not_i337;

assign local_bb4_cmp25_not_i337 = (local_bb4_cmp25_i334 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u38_stall_local;
wire local_bb4_var__u38;

assign local_bb4_var__u38 = (local_bb4_cmp25_i334 | rnode_178to180_bb4_cmp27_i335_2_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_3_VALID_195_196_0_inputs_ready;
 reg SFC_3_VALID_195_196_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_195_196_0_stall_in;
wire SFC_3_VALID_195_196_0_output_regs_ready;
 reg SFC_3_VALID_195_196_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_195_196_0_causedstall;

assign SFC_3_VALID_195_196_0_inputs_ready = 1'b1;
assign SFC_3_VALID_195_196_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_194_195_0_stall_in = 1'b0;
assign SFC_3_VALID_195_196_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_195_196_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_195_196_0_output_regs_ready)
		begin
			SFC_3_VALID_195_196_0_NO_SHIFT_REG <= SFC_3_VALID_194_195_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__28_i353_stall_local;
wire [31:0] local_bb4__28_i353;

assign local_bb4__28_i353 = (rnode_178to179_bb4_lnot23_i333_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl66_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i342_stall_local;
wire local_bb4_lnot30_not_i342;

assign local_bb4_lnot30_not_i342 = (local_bb4_lnot30_i338 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i351_stall_local;
wire [31:0] local_bb4_shl_i351;

assign local_bb4_shl_i351 = ((local_bb4_or_i350 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_and35_i336_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i336_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and35_i336_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i336_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and35_i336_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i336_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i336_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and35_i336_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_and35_i336_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_and35_i336_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_and35_i336_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_and35_i336_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_and35_i336_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in((rnode_180to182_bb4_and35_i336_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_182to183_bb4_and35_i336_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_and35_i336_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_and35_i336_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_and35_i336_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_and35_i336_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_and35_i336_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_and35_i336_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and35_i336_0_NO_SHIFT_REG = rnode_182to183_bb4_and35_i336_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_and35_i336_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and35_i336_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i339_stall_local;
wire local_bb4_or_cond_i339;

assign local_bb4_or_cond_i339 = (local_bb4_lnot30_i338 | local_bb4_cmp25_not_i337);

// This section implements a registered operation.
// 
wire SFC_3_VALID_196_197_0_inputs_ready;
 reg SFC_3_VALID_196_197_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_196_197_0_stall_in;
wire SFC_3_VALID_196_197_0_output_regs_ready;
 reg SFC_3_VALID_196_197_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_196_197_0_causedstall;

assign SFC_3_VALID_196_197_0_inputs_ready = 1'b1;
assign SFC_3_VALID_196_197_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_195_196_0_stall_in = 1'b0;
assign SFC_3_VALID_196_197_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_196_197_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_196_197_0_output_regs_ready)
		begin
			SFC_3_VALID_196_197_0_NO_SHIFT_REG <= SFC_3_VALID_195_196_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and73_i_stall_local;
wire [31:0] local_bb4_and73_i;

assign local_bb4_and73_i = ((local_bb4__28_i353 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and76_i_stall_local;
wire [31:0] local_bb4_and76_i;

assign local_bb4_and76_i = ((local_bb4__28_i353 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and79_i_stall_local;
wire [31:0] local_bb4_and79_i;

assign local_bb4_and79_i = ((local_bb4__28_i353 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr95_i_stall_local;
wire [31:0] local_bb4_shr95_i;

assign local_bb4_shr95_i = ((local_bb4__28_i353 & 32'h7FFFFF8) >> (local_bb4_and94_i & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and91_i_stall_local;
wire [31:0] local_bb4_and91_i;

assign local_bb4_and91_i = ((local_bb4__28_i353 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i357_stall_local;
wire [31:0] local_bb4_and88_i357;

assign local_bb4_and88_i357 = ((local_bb4__28_i353 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and85_i_stall_local;
wire [31:0] local_bb4_and85_i;

assign local_bb4_and85_i = ((local_bb4__28_i353 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u39_stall_local;
wire [31:0] local_bb4_var__u39;

assign local_bb4_var__u39 = ((local_bb4__28_i353 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i343_stall_local;
wire local_bb4_or_cond_not_i343;

assign local_bb4_or_cond_not_i343 = (local_bb4_cmp25_i334 & local_bb4_lnot30_not_i342);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i352_stall_local;
wire [31:0] local_bb4__27_i352;

assign local_bb4__27_i352 = (local_bb4_lnot_i332 ? 32'h0 : ((local_bb4_shl_i351 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i347_stall_local;
wire local_bb4_reduction_8_i347;

assign local_bb4_reduction_8_i347 = (rnode_178to180_bb4_cmp27_i335_1_NO_SHIFT_REG & local_bb4_or_cond_i339);

// This section implements a registered operation.
// 
wire SFC_3_VALID_197_198_0_inputs_ready;
 reg SFC_3_VALID_197_198_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_197_198_0_stall_in;
wire SFC_3_VALID_197_198_0_output_regs_ready;
 reg SFC_3_VALID_197_198_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_197_198_0_causedstall;

assign SFC_3_VALID_197_198_0_inputs_ready = 1'b1;
assign SFC_3_VALID_197_198_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_196_197_0_stall_in = 1'b0;
assign SFC_3_VALID_197_198_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_197_198_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_197_198_0_output_regs_ready)
		begin
			SFC_3_VALID_197_198_0_NO_SHIFT_REG <= SFC_3_VALID_196_197_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and73_tr_i_stall_local;
wire [7:0] local_bb4_and73_tr_i;
wire [31:0] local_bb4_and73_tr_i$ps;

assign local_bb4_and73_tr_i$ps = (local_bb4_and73_i & 32'hFFFFFF);
assign local_bb4_and73_tr_i = local_bb4_and73_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i356_stall_local;
wire local_bb4_cmp77_i356;

assign local_bb4_cmp77_i356 = ((local_bb4_and76_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp80_i_stall_local;
wire local_bb4_cmp80_i;

assign local_bb4_cmp80_i = ((local_bb4_and79_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and143_i_stall_local;
wire [31:0] local_bb4_and143_i;

assign local_bb4_and143_i = (local_bb4_shr95_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr151_i_stall_local;
wire [31:0] local_bb4_shr151_i;

assign local_bb4_shr151_i = (local_bb4_shr95_i >> (local_bb4_and150_i & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u40_stall_local;
wire [31:0] local_bb4_var__u40;

assign local_bb4_var__u40 = (local_bb4_shr95_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and147_i_stall_local;
wire [31:0] local_bb4_and147_i;

assign local_bb4_and147_i = (local_bb4_shr95_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp92_i_stall_local;
wire local_bb4_cmp92_i;

assign local_bb4_cmp92_i = ((local_bb4_and91_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp89_i_stall_local;
wire local_bb4_cmp89_i;

assign local_bb4_cmp89_i = ((local_bb4_and88_i357 & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp86_i_stall_local;
wire local_bb4_cmp86_i;

assign local_bb4_cmp86_i = ((local_bb4_and85_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u41_stall_local;
wire local_bb4_var__u41;

assign local_bb4_var__u41 = ((local_bb4_var__u39 & 32'hFFF8) != 32'h0);

// This section implements a registered operation.
// 
wire SFC_3_VALID_198_199_0_inputs_ready;
 reg SFC_3_VALID_198_199_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_198_199_0_stall_in;
wire SFC_3_VALID_198_199_0_output_regs_ready;
 reg SFC_3_VALID_198_199_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_198_199_0_causedstall;

assign SFC_3_VALID_198_199_0_inputs_ready = 1'b1;
assign SFC_3_VALID_198_199_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_197_198_0_stall_in = 1'b0;
assign SFC_3_VALID_198_199_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_198_199_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_198_199_0_output_regs_ready)
		begin
			SFC_3_VALID_198_199_0_NO_SHIFT_REG <= SFC_3_VALID_197_198_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_frombool75_i_stall_local;
wire [7:0] local_bb4_frombool75_i;

assign local_bb4_frombool75_i = (local_bb4_and73_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u42_stall_local;
wire [31:0] local_bb4_var__u42;

assign local_bb4_var__u42 = ((local_bb4_and147_i & 32'h3FFFFFFF) | local_bb4_shr95_i);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i361_stall_local;
wire local_bb4__31_v_i361;

assign local_bb4__31_v_i361 = (local_bb4_cmp97_i ? local_bb4_cmp80_i : local_bb4_cmp92_i);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i359_stall_local;
wire local_bb4__30_v_i359;

assign local_bb4__30_v_i359 = (local_bb4_cmp97_i ? local_bb4_cmp77_i356 : local_bb4_cmp89_i);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool110_i_stall_local;
wire [7:0] local_bb4_frombool110_i;

assign local_bb4_frombool110_i[7:1] = 7'h0;
assign local_bb4_frombool110_i[0] = local_bb4_cmp86_i;

// This section implements an unregistered operation.
// 
wire local_bb4_or108_i_stall_local;
wire [31:0] local_bb4_or108_i;

assign local_bb4_or108_i[31:1] = 31'h0;
assign local_bb4_or108_i[0] = local_bb4_var__u41;

// This section implements a registered operation.
// 
wire SFC_3_VALID_199_200_0_inputs_ready;
 reg SFC_3_VALID_199_200_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_199_200_0_stall_in;
wire SFC_3_VALID_199_200_0_output_regs_ready;
 reg SFC_3_VALID_199_200_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_199_200_0_causedstall;

assign SFC_3_VALID_199_200_0_inputs_ready = 1'b1;
assign SFC_3_VALID_199_200_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_198_199_0_stall_in = 1'b0;
assign SFC_3_VALID_199_200_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_199_200_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_199_200_0_output_regs_ready)
		begin
			SFC_3_VALID_199_200_0_NO_SHIFT_REG <= SFC_3_VALID_198_199_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or1606_i_stall_local;
wire [31:0] local_bb4_or1606_i;

assign local_bb4_or1606_i = (local_bb4_var__u42 | (local_bb4_and143_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i362_stall_local;
wire [7:0] local_bb4__31_i362;

assign local_bb4__31_i362[7:1] = 7'h0;
assign local_bb4__31_i362[0] = local_bb4__31_v_i361;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i360_stall_local;
wire [7:0] local_bb4__30_i360;

assign local_bb4__30_i360[7:1] = 7'h0;
assign local_bb4__30_i360[0] = local_bb4__30_v_i359;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i358_stall_local;
wire [7:0] local_bb4__29_i358;

assign local_bb4__29_i358 = (local_bb4_cmp97_i ? (local_bb4_frombool75_i & 8'h1) : (local_bb4_frombool110_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i363_stall_local;
wire [31:0] local_bb4__32_i363;

assign local_bb4__32_i363 = (local_bb4_cmp97_i ? 32'h0 : (local_bb4_or108_i & 32'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_200_201_0_inputs_ready;
 reg SFC_3_VALID_200_201_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_200_201_0_stall_in;
wire SFC_3_VALID_200_201_0_output_regs_ready;
 reg SFC_3_VALID_200_201_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_200_201_0_causedstall;

assign SFC_3_VALID_200_201_0_inputs_ready = 1'b1;
assign SFC_3_VALID_200_201_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_199_200_0_stall_in = 1'b0;
assign SFC_3_VALID_200_201_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_200_201_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_200_201_0_output_regs_ready)
		begin
			SFC_3_VALID_200_201_0_NO_SHIFT_REG <= SFC_3_VALID_199_200_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or163_i_stall_local;
wire [31:0] local_bb4_or163_i;

assign local_bb4_or163_i = (local_bb4_or1606_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1247_i_stall_local;
wire [7:0] local_bb4_or1247_i;

assign local_bb4_or1247_i = ((local_bb4__30_i360 & 8'h1) | (local_bb4__29_i358 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i365_stall_local;
wire [7:0] local_bb4__33_i365;

assign local_bb4__33_i365 = (local_bb4_cmp117_i ? (local_bb4__29_i358 & 8'h1) : (local_bb4__31_i362 & 8'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_201_202_0_inputs_ready;
 reg SFC_3_VALID_201_202_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_201_202_0_stall_in;
wire SFC_3_VALID_201_202_0_output_regs_ready;
 reg SFC_3_VALID_201_202_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_201_202_0_causedstall;

assign SFC_3_VALID_201_202_0_inputs_ready = 1'b1;
assign SFC_3_VALID_201_202_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_200_201_0_stall_in = 1'b0;
assign SFC_3_VALID_201_202_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_201_202_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_201_202_0_output_regs_ready)
		begin
			SFC_3_VALID_201_202_0_NO_SHIFT_REG <= SFC_3_VALID_200_201_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i368_stall_local;
wire [31:0] local_bb4__37_v_i368;

assign local_bb4__37_v_i368 = (local_bb4_Pivot20_i366 ? 32'h0 : (local_bb4_or163_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i364_stall_local;
wire [31:0] local_bb4_or124_i364;

assign local_bb4_or124_i364[31:8] = 24'h0;
assign local_bb4_or124_i364[7:0] = (local_bb4_or1247_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u43_stall_local;
wire [7:0] local_bb4_var__u43;

assign local_bb4_var__u43 = ((local_bb4__33_i365 & 8'h1) & 8'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_202_203_0_inputs_ready;
 reg SFC_3_VALID_202_203_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_202_203_0_stall_in;
wire SFC_3_VALID_202_203_0_output_regs_ready;
 reg SFC_3_VALID_202_203_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_202_203_0_causedstall;

assign SFC_3_VALID_202_203_0_inputs_ready = 1'b1;
assign SFC_3_VALID_202_203_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_201_202_0_stall_in = 1'b0;
assign SFC_3_VALID_202_203_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_202_203_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_202_203_0_output_regs_ready)
		begin
			SFC_3_VALID_202_203_0_NO_SHIFT_REG <= SFC_3_VALID_201_202_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i369_stall_local;
wire [31:0] local_bb4__39_v_i369;

assign local_bb4__39_v_i369 = (local_bb4_SwitchLeaf_i367 ? (local_bb4_var__u40 & 32'h1) : (local_bb4__37_v_i368 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or125_i_stall_local;
wire [31:0] local_bb4_or125_i;

assign local_bb4_or125_i = (local_bb4_cmp117_i ? 32'h0 : (local_bb4_or124_i364 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv136_i_stall_local;
wire [31:0] local_bb4_conv136_i;

assign local_bb4_conv136_i[31:8] = 24'h0;
assign local_bb4_conv136_i[7:0] = (local_bb4_var__u43 & 8'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_203_204_0_inputs_ready;
 reg SFC_3_VALID_203_204_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_203_204_0_stall_in;
wire SFC_3_VALID_203_204_0_output_regs_ready;
 reg SFC_3_VALID_203_204_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_203_204_0_causedstall;

assign SFC_3_VALID_203_204_0_inputs_ready = 1'b1;
assign SFC_3_VALID_203_204_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_202_203_0_stall_in = 1'b0;
assign SFC_3_VALID_203_204_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_203_204_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_203_204_0_output_regs_ready)
		begin
			SFC_3_VALID_203_204_0_NO_SHIFT_REG <= SFC_3_VALID_202_203_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i370_stall_local;
wire [31:0] local_bb4_reduction_3_i370;

assign local_bb4_reduction_3_i370 = ((local_bb4__32_i363 & 32'h1) | (local_bb4_or125_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or137_i_stall_local;
wire [31:0] local_bb4_or137_i;

assign local_bb4_or137_i = (local_bb4_cmp132_not_i ? (local_bb4_conv136_i & 32'h1) : 32'h0);

// This section implements a registered operation.
// 
wire SFC_3_VALID_204_205_0_inputs_ready;
 reg SFC_3_VALID_204_205_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_204_205_0_stall_in;
wire SFC_3_VALID_204_205_0_output_regs_ready;
 reg SFC_3_VALID_204_205_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_204_205_0_causedstall;

assign SFC_3_VALID_204_205_0_inputs_ready = 1'b1;
assign SFC_3_VALID_204_205_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_203_204_0_stall_in = 1'b0;
assign SFC_3_VALID_204_205_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_204_205_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_204_205_0_output_regs_ready)
		begin
			SFC_3_VALID_204_205_0_NO_SHIFT_REG <= SFC_3_VALID_203_204_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i372_stall_local;
wire [31:0] local_bb4_reduction_5_i372;

assign local_bb4_reduction_5_i372 = (local_bb4_shr151_i | (local_bb4_reduction_3_i370 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i371_stall_local;
wire [31:0] local_bb4_reduction_4_i371;

assign local_bb4_reduction_4_i371 = ((local_bb4_or137_i & 32'h1) | (local_bb4__39_v_i369 & 32'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_205_206_0_inputs_ready;
 reg SFC_3_VALID_205_206_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_205_206_0_stall_in;
wire SFC_3_VALID_205_206_0_output_regs_ready;
 reg SFC_3_VALID_205_206_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_205_206_0_causedstall;

assign SFC_3_VALID_205_206_0_inputs_ready = 1'b1;
assign SFC_3_VALID_205_206_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_204_205_0_stall_in = 1'b0;
assign SFC_3_VALID_205_206_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_205_206_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_205_206_0_output_regs_ready)
		begin
			SFC_3_VALID_205_206_0_NO_SHIFT_REG <= SFC_3_VALID_204_205_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i373_stall_local;
wire [31:0] local_bb4_reduction_6_i373;

assign local_bb4_reduction_6_i373 = ((local_bb4_reduction_4_i371 & 32'h1) | local_bb4_reduction_5_i372);

// This section implements a registered operation.
// 
wire SFC_3_VALID_206_207_0_inputs_ready;
 reg SFC_3_VALID_206_207_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_206_207_0_stall_in;
wire SFC_3_VALID_206_207_0_output_regs_ready;
 reg SFC_3_VALID_206_207_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_206_207_0_causedstall;

assign SFC_3_VALID_206_207_0_inputs_ready = 1'b1;
assign SFC_3_VALID_206_207_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_205_206_0_stall_in = 1'b0;
assign SFC_3_VALID_206_207_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_206_207_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_206_207_0_output_regs_ready)
		begin
			SFC_3_VALID_206_207_0_NO_SHIFT_REG <= SFC_3_VALID_205_206_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i340_valid_out;
wire local_bb4_lnot33_not_i340_stall_in;
wire local_bb4_cmp38_i_valid_out;
wire local_bb4_cmp38_i_stall_in;
wire local_bb4_and37_lobit_i_valid_out;
wire local_bb4_and37_lobit_i_stall_in;
wire local_bb4_xor189_i_valid_out;
wire local_bb4_xor189_i_stall_in;
wire local_bb4_xor189_i_inputs_ready;
wire local_bb4_xor189_i_stall_local;
wire [31:0] local_bb4_xor189_i;

assign local_bb4_xor189_i_inputs_ready = (rnode_178to179_bb4__22_i324_0_valid_out_0_NO_SHIFT_REG & rnode_178to179_bb4_lnot23_i333_0_valid_out_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i355_0_valid_out_0_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i355_0_valid_out_4_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i355_0_valid_out_1_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i355_0_valid_out_2_NO_SHIFT_REG & rnode_178to179_bb4_align_0_i355_0_valid_out_3_NO_SHIFT_REG & rnode_178to179_bb4__23_i325_0_valid_out_2_NO_SHIFT_REG & rnode_178to179_bb4__22_i324_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor189_i = (local_bb4_reduction_6_i373 ^ local_bb4_xor36_lobit_i);
assign local_bb4_lnot33_not_i340_valid_out = 1'b1;
assign local_bb4_cmp38_i_valid_out = 1'b1;
assign local_bb4_and37_lobit_i_valid_out = 1'b1;
assign local_bb4_xor189_i_valid_out = 1'b1;
assign rnode_178to179_bb4__22_i324_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_lnot23_i333_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i355_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i355_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i355_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i355_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4_align_0_i355_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__23_i325_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb4__22_i324_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_207_208_0_inputs_ready;
 reg SFC_3_VALID_207_208_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_207_208_0_stall_in;
wire SFC_3_VALID_207_208_0_output_regs_ready;
 reg SFC_3_VALID_207_208_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_207_208_0_causedstall;

assign SFC_3_VALID_207_208_0_inputs_ready = 1'b1;
assign SFC_3_VALID_207_208_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_206_207_0_stall_in = 1'b0;
assign SFC_3_VALID_207_208_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_207_208_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_207_208_0_output_regs_ready)
		begin
			SFC_3_VALID_207_208_0_NO_SHIFT_REG <= SFC_3_VALID_206_207_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_lnot33_not_i340_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i340_0_stall_in_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i340_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i340_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i340_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i340_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i340_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_lnot33_not_i340_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_lnot33_not_i340_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_lnot33_not_i340_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_lnot33_not_i340_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_lnot33_not_i340_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_lnot33_not_i340_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i340),
	.data_out(rnode_179to180_bb4_lnot33_not_i340_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_lnot33_not_i340_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_lnot33_not_i340_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb4_lnot33_not_i340_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_lnot33_not_i340_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_lnot33_not_i340_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i340_stall_in = 1'b0;
assign rnode_179to180_bb4_lnot33_not_i340_0_NO_SHIFT_REG = rnode_179to180_bb4_lnot33_not_i340_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_lnot33_not_i340_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_lnot33_not_i340_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_cmp38_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_cmp38_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_cmp38_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_cmp38_i_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_cmp38_i_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_cmp38_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_cmp38_i),
	.data_out(rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_cmp38_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_cmp38_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp38_i_stall_in = 1'b0;
assign rnode_179to180_bb4_cmp38_i_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp38_i_0_NO_SHIFT_REG = rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp38_i_1_NO_SHIFT_REG = rnode_179to180_bb4_cmp38_i_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and37_lobit_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_and37_lobit_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_and37_lobit_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_and37_lobit_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_and37_lobit_i_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_and37_lobit_i_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_and37_lobit_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in((local_bb4_and37_lobit_i & 32'h1)),
	.data_out(rnode_179to180_bb4_and37_lobit_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_and37_lobit_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_and37_lobit_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and37_lobit_i_stall_in = 1'b0;
assign rnode_179to180_bb4_and37_lobit_i_0_NO_SHIFT_REG = rnode_179to180_bb4_and37_lobit_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_and37_lobit_i_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb4_xor189_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_xor189_i_0_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb4_xor189_i_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb4_xor189_i_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb4_xor189_i_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb4_xor189_i_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb4_xor189_i_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb4_xor189_i_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb4_xor189_i_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb4_xor189_i),
	.data_out(rnode_179to180_bb4_xor189_i_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb4_xor189_i_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb4_xor189_i_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor189_i_stall_in = 1'b0;
assign rnode_179to180_bb4_xor189_i_0_NO_SHIFT_REG = rnode_179to180_bb4_xor189_i_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb4_xor189_i_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_xor189_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_208_209_0_inputs_ready;
 reg SFC_3_VALID_208_209_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_208_209_0_stall_in;
wire SFC_3_VALID_208_209_0_output_regs_ready;
 reg SFC_3_VALID_208_209_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_208_209_0_causedstall;

assign SFC_3_VALID_208_209_0_inputs_ready = 1'b1;
assign SFC_3_VALID_208_209_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_207_208_0_stall_in = 1'b0;
assign SFC_3_VALID_208_209_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_208_209_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_208_209_0_output_regs_ready)
		begin
			SFC_3_VALID_208_209_0_NO_SHIFT_REG <= SFC_3_VALID_207_208_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i341_stall_local;
wire local_bb4_brmerge_not_i341;

assign local_bb4_brmerge_not_i341 = (rnode_178to180_bb4_cmp27_i335_0_NO_SHIFT_REG & rnode_179to180_bb4_lnot33_not_i340_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_2_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_cmp38_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_cmp38_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_cmp38_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_cmp38_i_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_cmp38_i_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_cmp38_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_179to180_bb4_cmp38_i_1_NO_SHIFT_REG),
	.data_out(rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_cmp38_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_cmp38_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp38_i_0_NO_SHIFT_REG = rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp38_i_1_NO_SHIFT_REG = rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb4_cmp38_i_2_NO_SHIFT_REG = rnode_180to182_bb4_cmp38_i_0_reg_182_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i374_stall_local;
wire [31:0] local_bb4_add_i374;

assign local_bb4_add_i374 = ((local_bb4__27_i352 & 32'h7FFFFF8) | (rnode_179to180_bb4_and37_lobit_i_0_NO_SHIFT_REG & 32'h1));

// This section implements a registered operation.
// 
wire SFC_3_VALID_209_210_0_inputs_ready;
 reg SFC_3_VALID_209_210_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_209_210_0_stall_in;
wire SFC_3_VALID_209_210_0_output_regs_ready;
 reg SFC_3_VALID_209_210_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_209_210_0_causedstall;

assign SFC_3_VALID_209_210_0_inputs_ready = 1'b1;
assign SFC_3_VALID_209_210_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_208_209_0_stall_in = 1'b0;
assign SFC_3_VALID_209_210_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_209_210_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_209_210_0_output_regs_ready)
		begin
			SFC_3_VALID_209_210_0_NO_SHIFT_REG <= SFC_3_VALID_208_209_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__24_i344_stall_local;
wire local_bb4__24_i344;

assign local_bb4__24_i344 = (local_bb4_or_cond_not_i343 | local_bb4_brmerge_not_i341);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i345_stall_local;
wire local_bb4_brmerge_not_not_i345;

assign local_bb4_brmerge_not_not_i345 = (local_bb4_brmerge_not_i341 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp38_i_stall_local;
wire local_bb4_not_cmp38_i;

assign local_bb4_not_cmp38_i = (rnode_180to182_bb4_cmp38_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add193_i_stall_local;
wire [31:0] local_bb4_add193_i;

assign local_bb4_add193_i = ((local_bb4_add_i374 & 32'h7FFFFF9) + rnode_179to180_bb4_xor189_i_0_NO_SHIFT_REG);

// This section implements a registered operation.
// 
wire SFC_3_VALID_210_211_0_inputs_ready;
 reg SFC_3_VALID_210_211_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_210_211_0_stall_in;
wire SFC_3_VALID_210_211_0_output_regs_ready;
 reg SFC_3_VALID_210_211_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_210_211_0_causedstall;

assign SFC_3_VALID_210_211_0_inputs_ready = 1'b1;
assign SFC_3_VALID_210_211_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_209_210_0_stall_in = 1'b0;
assign SFC_3_VALID_210_211_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_210_211_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_210_211_0_output_regs_ready)
		begin
			SFC_3_VALID_210_211_0_NO_SHIFT_REG <= SFC_3_VALID_209_210_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i346_stall_local;
wire local_bb4_reduction_7_i346;

assign local_bb4_reduction_7_i346 = (local_bb4_cmp25_i334 & local_bb4_brmerge_not_not_i345);

// This section implements a registered operation.
// 
wire SFC_3_VALID_211_212_0_inputs_ready;
 reg SFC_3_VALID_211_212_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_211_212_0_stall_in;
wire SFC_3_VALID_211_212_0_output_regs_ready;
 reg SFC_3_VALID_211_212_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_211_212_0_causedstall;

assign SFC_3_VALID_211_212_0_inputs_ready = 1'b1;
assign SFC_3_VALID_211_212_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_210_211_0_stall_in = 1'b0;
assign SFC_3_VALID_211_212_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_211_212_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_211_212_0_output_regs_ready)
		begin
			SFC_3_VALID_211_212_0_NO_SHIFT_REG <= SFC_3_VALID_210_211_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i348_stall_local;
wire local_bb4_reduction_9_i348;

assign local_bb4_reduction_9_i348 = (local_bb4_reduction_7_i346 & local_bb4_reduction_8_i347);

// This section implements a registered operation.
// 
wire SFC_3_VALID_212_213_0_inputs_ready;
 reg SFC_3_VALID_212_213_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_212_213_0_stall_in;
wire SFC_3_VALID_212_213_0_output_regs_ready;
 reg SFC_3_VALID_212_213_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_212_213_0_causedstall;

assign SFC_3_VALID_212_213_0_inputs_ready = 1'b1;
assign SFC_3_VALID_212_213_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_211_212_0_stall_in = 1'b0;
assign SFC_3_VALID_212_213_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_212_213_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_212_213_0_output_regs_ready)
		begin
			SFC_3_VALID_212_213_0_NO_SHIFT_REG <= SFC_3_VALID_211_212_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and17_i327_valid_out_2;
wire local_bb4_and17_i327_stall_in_2;
wire local_bb4_var__u38_valid_out;
wire local_bb4_var__u38_stall_in;
wire local_bb4_add193_i_valid_out;
wire local_bb4_add193_i_stall_in;
wire local_bb4__26_i349_valid_out;
wire local_bb4__26_i349_stall_in;
wire local_bb4__26_i349_inputs_ready;
wire local_bb4__26_i349_stall_local;
wire local_bb4__26_i349;

assign local_bb4__26_i349_inputs_ready = (rnode_178to180_bb4_shr16_i326_0_valid_out_0_NO_SHIFT_REG & rnode_178to180_bb4_cmp27_i335_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb4_and37_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_179to180_bb4_xor189_i_0_valid_out_NO_SHIFT_REG & rnode_179to180_bb4_and20_i330_0_valid_out_0_NO_SHIFT_REG & rnode_178to180_bb4_cmp27_i335_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb4_lnot33_not_i340_0_valid_out_NO_SHIFT_REG & rnode_178to180_bb4_cmp27_i335_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb4_and20_i330_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i349 = (local_bb4_reduction_9_i348 ? rnode_179to180_bb4_cmp38_i_0_NO_SHIFT_REG : local_bb4__24_i344);
assign local_bb4_and17_i327_valid_out_2 = 1'b1;
assign local_bb4_var__u38_valid_out = 1'b1;
assign local_bb4_add193_i_valid_out = 1'b1;
assign local_bb4__26_i349_valid_out = 1'b1;
assign rnode_178to180_bb4_shr16_i326_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i335_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and37_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_xor189_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and20_i330_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i335_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_lnot33_not_i340_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to180_bb4_cmp27_i335_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_and20_i330_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_213_214_0_inputs_ready;
 reg SFC_3_VALID_213_214_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_213_214_0_stall_in;
wire SFC_3_VALID_213_214_0_output_regs_ready;
 reg SFC_3_VALID_213_214_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_213_214_0_causedstall;

assign SFC_3_VALID_213_214_0_inputs_ready = 1'b1;
assign SFC_3_VALID_213_214_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_212_213_0_stall_in = 1'b0;
assign SFC_3_VALID_213_214_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_213_214_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_213_214_0_output_regs_ready)
		begin
			SFC_3_VALID_213_214_0_NO_SHIFT_REG <= SFC_3_VALID_212_213_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb4_and17_i327_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i327_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and17_i327_0_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i327_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb4_and17_i327_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i327_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i327_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb4_and17_i327_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb4_and17_i327_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb4_and17_i327_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb4_and17_i327_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb4_and17_i327_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb4_and17_i327_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i327 & 32'hFF)),
	.data_out(rnode_180to182_bb4_and17_i327_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb4_and17_i327_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb4_and17_i327_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb4_and17_i327_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb4_and17_i327_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb4_and17_i327_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i327_stall_in_2 = 1'b0;
assign rnode_180to182_bb4_and17_i327_0_NO_SHIFT_REG = rnode_180to182_bb4_and17_i327_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb4_and17_i327_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and17_i327_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_var__u38_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u38_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u38_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u38_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u38_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u38_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u38_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_var__u38_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_var__u38_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_var__u38_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_var__u38_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_var__u38_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_var__u38_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4_var__u38),
	.data_out(rnode_180to181_bb4_var__u38_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_var__u38_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_var__u38_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb4_var__u38_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_var__u38_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_var__u38_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u38_stall_in = 1'b0;
assign rnode_180to181_bb4_var__u38_0_NO_SHIFT_REG = rnode_180to181_bb4_var__u38_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_var__u38_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_var__u38_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_1_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_2_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_3_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4_add193_i_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4_add193_i_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4_add193_i_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4_add193_i_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4_add193_i_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4_add193_i_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4_add193_i),
	.data_out(rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4_add193_i_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4_add193_i_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add193_i_stall_in = 1'b0;
assign rnode_180to181_bb4_add193_i_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_0_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_1_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_2_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_add193_i_3_NO_SHIFT_REG = rnode_180to181_bb4_add193_i_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb4__26_i349_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i349_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i349_0_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i349_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i349_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i349_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i349_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb4__26_i349_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb4__26_i349_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb4__26_i349_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb4__26_i349_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb4__26_i349_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb4__26_i349_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb4__26_i349),
	.data_out(rnode_180to181_bb4__26_i349_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb4__26_i349_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb4__26_i349_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb4__26_i349_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb4__26_i349_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb4__26_i349_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i349_stall_in = 1'b0;
assign rnode_180to181_bb4__26_i349_0_NO_SHIFT_REG = rnode_180to181_bb4__26_i349_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb4__26_i349_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb4__26_i349_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_214_215_0_inputs_ready;
 reg SFC_3_VALID_214_215_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_214_215_0_stall_in;
wire SFC_3_VALID_214_215_0_output_regs_ready;
 reg SFC_3_VALID_214_215_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_214_215_0_causedstall;

assign SFC_3_VALID_214_215_0_inputs_ready = 1'b1;
assign SFC_3_VALID_214_215_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_213_214_0_stall_in = 1'b0;
assign SFC_3_VALID_214_215_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_214_215_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_214_215_0_output_regs_ready)
		begin
			SFC_3_VALID_214_215_0_NO_SHIFT_REG <= SFC_3_VALID_213_214_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_var__u38_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u38_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u38_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u38_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u38_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u38_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u38_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_var__u38_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_var__u38_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_var__u38_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_var__u38_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_var__u38_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_var__u38_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb4_var__u38_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb4_var__u38_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_var__u38_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_var__u38_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb4_var__u38_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_var__u38_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_var__u38_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4_var__u38_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_var__u38_0_NO_SHIFT_REG = rnode_181to182_bb4_var__u38_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_var__u38_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_var__u38_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and194_i_valid_out;
wire local_bb4_and194_i_stall_in;
wire local_bb4_and194_i_inputs_ready;
wire local_bb4_and194_i_stall_local;
wire [31:0] local_bb4_and194_i;

assign local_bb4_and194_i_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and194_i = (rnode_180to181_bb4_add193_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and194_i_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and196_i_valid_out;
wire local_bb4_and196_i_stall_in;
wire local_bb4_and196_i_inputs_ready;
wire local_bb4_and196_i_stall_local;
wire [31:0] local_bb4_and196_i;

assign local_bb4_and196_i_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and196_i = (rnode_180to181_bb4_add193_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and196_i_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and199_i_valid_out;
wire local_bb4_and199_i_stall_in;
wire local_bb4_and199_i_inputs_ready;
wire local_bb4_and199_i_stall_local;
wire [31:0] local_bb4_and199_i;

assign local_bb4_and199_i_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and199_i = (rnode_180to181_bb4_add193_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and199_i_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and202_i_stall_local;
wire [31:0] local_bb4_and202_i;

assign local_bb4_and202_i = (rnode_180to181_bb4_add193_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_181to183_bb4__26_i349_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i349_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i349_0_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i349_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i349_0_reg_183_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i349_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i349_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_181to183_bb4__26_i349_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_181to183_bb4__26_i349_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to183_bb4__26_i349_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to183_bb4__26_i349_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_181to183_bb4__26_i349_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_181to183_bb4__26_i349_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb4__26_i349_0_NO_SHIFT_REG),
	.data_out(rnode_181to183_bb4__26_i349_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_181to183_bb4__26_i349_0_reg_183_fifo.DEPTH = 2;
defparam rnode_181to183_bb4__26_i349_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_181to183_bb4__26_i349_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to183_bb4__26_i349_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_181to183_bb4__26_i349_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb4__26_i349_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to183_bb4__26_i349_0_NO_SHIFT_REG = rnode_181to183_bb4__26_i349_0_reg_183_NO_SHIFT_REG;
assign rnode_181to183_bb4__26_i349_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_181to183_bb4__26_i349_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_215_216_0_inputs_ready;
 reg SFC_3_VALID_215_216_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_215_216_0_stall_in;
wire SFC_3_VALID_215_216_0_output_regs_ready;
 reg SFC_3_VALID_215_216_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_215_216_0_causedstall;

assign SFC_3_VALID_215_216_0_inputs_ready = 1'b1;
assign SFC_3_VALID_215_216_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_214_215_0_stall_in = 1'b0;
assign SFC_3_VALID_215_216_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_215_216_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_215_216_0_output_regs_ready)
		begin
			SFC_3_VALID_215_216_0_NO_SHIFT_REG <= SFC_3_VALID_214_215_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_var__u38_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u38_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u38_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u38_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u38_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u38_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u38_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_var__u38_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_var__u38_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_var__u38_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_var__u38_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_var__u38_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_var__u38_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb4_var__u38_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb4_var__u38_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_var__u38_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_var__u38_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4_var__u38_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_var__u38_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_var__u38_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_var__u38_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u38_0_NO_SHIFT_REG = rnode_182to183_bb4_var__u38_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_var__u38_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u38_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and194_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and194_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and194_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and194_i_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and194_i_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and194_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and194_i & 32'hFFFFFFF)),
	.data_out(rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and194_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and194_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and194_i_stall_in = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and194_i_0_NO_SHIFT_REG = rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and194_i_1_NO_SHIFT_REG = rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4_and194_i_2_NO_SHIFT_REG = rnode_181to182_bb4_and194_i_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and196_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and196_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and196_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and196_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and196_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and196_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and196_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and196_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and196_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and196_i & 32'h1F)),
	.data_out(rnode_181to182_bb4_and196_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and196_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and196_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and196_i_stall_in = 1'b0;
assign rnode_181to182_bb4_and196_i_0_NO_SHIFT_REG = rnode_181to182_bb4_and196_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and196_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and196_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4_and199_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and199_i_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4_and199_i_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4_and199_i_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4_and199_i_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4_and199_i_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4_and199_i_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4_and199_i_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4_and199_i_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4_and199_i & 32'h1)),
	.data_out(rnode_181to182_bb4_and199_i_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4_and199_i_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4_and199_i_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and199_i_stall_in = 1'b0;
assign rnode_181to182_bb4_and199_i_0_NO_SHIFT_REG = rnode_181to182_bb4_and199_i_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4_and199_i_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and199_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i375_stall_local;
wire [31:0] local_bb4_shr_i_i375;

assign local_bb4_shr_i_i375 = ((local_bb4_and202_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4__26_i349_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__26_i349_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4__26_i349_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4__26_i349_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4__26_i349_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4__26_i349_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4__26_i349_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_181to183_bb4__26_i349_0_NO_SHIFT_REG),
	.data_out(rnode_183to184_bb4__26_i349_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4__26_i349_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4__26_i349_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4__26_i349_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4__26_i349_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4__26_i349_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to183_bb4__26_i349_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i349_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i349_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__26_i349_0_NO_SHIFT_REG = rnode_183to184_bb4__26_i349_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__26_i349_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__26_i349_1_NO_SHIFT_REG = rnode_183to184_bb4__26_i349_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__26_i349_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__26_i349_2_NO_SHIFT_REG = rnode_183to184_bb4__26_i349_0_reg_184_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_216_217_0_inputs_ready;
 reg SFC_3_VALID_216_217_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_216_217_0_stall_in;
wire SFC_3_VALID_216_217_0_output_regs_ready;
 reg SFC_3_VALID_216_217_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_216_217_0_causedstall;

assign SFC_3_VALID_216_217_0_inputs_ready = 1'b1;
assign SFC_3_VALID_216_217_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_215_216_0_stall_in = 1'b0;
assign SFC_3_VALID_216_217_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_216_217_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_216_217_0_output_regs_ready)
		begin
			SFC_3_VALID_216_217_0_NO_SHIFT_REG <= SFC_3_VALID_215_216_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr217_i_stall_local;
wire [31:0] local_bb4_shr217_i;

assign local_bb4_shr217_i = ((rnode_181to182_bb4_and194_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i389_stall_local;
wire [31:0] local_bb4__pre_i389;

assign local_bb4__pre_i389 = ((rnode_181to182_bb4_and196_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i376_stall_local;
wire [31:0] local_bb4_or_i_i376;

assign local_bb4_or_i_i376 = ((local_bb4_shr_i_i375 & 32'h3FFFFFF) | (local_bb4_and202_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond293_i_stall_local;
wire [31:0] local_bb4_cond293_i;

assign local_bb4_cond293_i = (rnode_183to184_bb4__26_i349_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u44_stall_local;
wire [31:0] local_bb4_var__u44;

assign local_bb4_var__u44[31:1] = 31'h0;
assign local_bb4_var__u44[0] = rnode_183to184_bb4__26_i349_2_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_217_218_0_inputs_ready;
 reg SFC_3_VALID_217_218_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_217_218_0_stall_in;
wire SFC_3_VALID_217_218_0_output_regs_ready;
 reg SFC_3_VALID_217_218_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_217_218_0_causedstall;

assign SFC_3_VALID_217_218_0_inputs_ready = 1'b1;
assign SFC_3_VALID_217_218_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_216_217_0_stall_in = 1'b0;
assign SFC_3_VALID_217_218_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_217_218_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_217_218_0_output_regs_ready)
		begin
			SFC_3_VALID_217_218_0_NO_SHIFT_REG <= SFC_3_VALID_216_217_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or220_i_stall_local;
wire [31:0] local_bb4_or220_i;

assign local_bb4_or220_i = ((local_bb4_shr217_i & 32'h7FFFFFF) | (rnode_181to182_bb4_and199_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool214_i_stall_local;
wire local_bb4_tobool214_i;

assign local_bb4_tobool214_i = ((local_bb4__pre_i389 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i377_stall_local;
wire [31:0] local_bb4_shr1_i_i377;

assign local_bb4_shr1_i_i377 = ((local_bb4_or_i_i376 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i406_stall_local;
wire [31:0] local_bb4_lnot_ext_i406;

assign local_bb4_lnot_ext_i406 = ((local_bb4_var__u44 & 32'h1) ^ 32'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_218_219_0_inputs_ready;
 reg SFC_3_VALID_218_219_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_218_219_0_stall_in;
wire SFC_3_VALID_218_219_0_output_regs_ready;
 reg SFC_3_VALID_218_219_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_218_219_0_causedstall;

assign SFC_3_VALID_218_219_0_inputs_ready = 1'b1;
assign SFC_3_VALID_218_219_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_217_218_0_stall_in = 1'b0;
assign SFC_3_VALID_218_219_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_218_219_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_218_219_0_output_regs_ready)
		begin
			SFC_3_VALID_218_219_0_NO_SHIFT_REG <= SFC_3_VALID_217_218_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i390_stall_local;
wire local_bb4__40_demorgan_i390;

assign local_bb4__40_demorgan_i390 = (rnode_180to182_bb4_cmp38_i_0_NO_SHIFT_REG | local_bb4_tobool214_i);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i391_stall_local;
wire local_bb4__42_i391;

assign local_bb4__42_i391 = (local_bb4_tobool214_i & local_bb4_not_cmp38_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i378_stall_local;
wire [31:0] local_bb4_or2_i_i378;

assign local_bb4_or2_i_i378 = ((local_bb4_shr1_i_i377 & 32'h1FFFFFF) | (local_bb4_or_i_i376 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_219_220_0_inputs_ready;
 reg SFC_3_VALID_219_220_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_219_220_0_stall_in;
wire SFC_3_VALID_219_220_0_output_regs_ready;
 reg SFC_3_VALID_219_220_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_219_220_0_causedstall;

assign SFC_3_VALID_219_220_0_inputs_ready = 1'b1;
assign SFC_3_VALID_219_220_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_218_219_0_stall_in = 1'b0;
assign SFC_3_VALID_219_220_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_219_220_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_219_220_0_output_regs_ready)
		begin
			SFC_3_VALID_219_220_0_NO_SHIFT_REG <= SFC_3_VALID_218_219_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__43_i392_stall_local;
wire [31:0] local_bb4__43_i392;

assign local_bb4__43_i392 = (local_bb4__42_i391 ? 32'h0 : (local_bb4__pre_i389 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i379_stall_local;
wire [31:0] local_bb4_shr3_i_i379;

assign local_bb4_shr3_i_i379 = ((local_bb4_or2_i_i378 & 32'h7FFFFFF) >> 32'h4);

// This section implements a registered operation.
// 
wire SFC_3_VALID_220_221_0_inputs_ready;
 reg SFC_3_VALID_220_221_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_220_221_0_stall_in;
wire SFC_3_VALID_220_221_0_output_regs_ready;
 reg SFC_3_VALID_220_221_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_220_221_0_causedstall;

assign SFC_3_VALID_220_221_0_inputs_ready = 1'b1;
assign SFC_3_VALID_220_221_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_219_220_0_stall_in = 1'b0;
assign SFC_3_VALID_220_221_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_220_221_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_220_221_0_output_regs_ready)
		begin
			SFC_3_VALID_220_221_0_NO_SHIFT_REG <= SFC_3_VALID_219_220_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i380_stall_local;
wire [31:0] local_bb4_or4_i_i380;

assign local_bb4_or4_i_i380 = ((local_bb4_shr3_i_i379 & 32'h7FFFFF) | (local_bb4_or2_i_i378 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_221_222_0_inputs_ready;
 reg SFC_3_VALID_221_222_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_221_222_0_stall_in;
wire SFC_3_VALID_221_222_0_output_regs_ready;
 reg SFC_3_VALID_221_222_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_221_222_0_causedstall;

assign SFC_3_VALID_221_222_0_inputs_ready = 1'b1;
assign SFC_3_VALID_221_222_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_220_221_0_stall_in = 1'b0;
assign SFC_3_VALID_221_222_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_221_222_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_221_222_0_output_regs_ready)
		begin
			SFC_3_VALID_221_222_0_NO_SHIFT_REG <= SFC_3_VALID_220_221_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i381_stall_local;
wire [31:0] local_bb4_shr5_i_i381;

assign local_bb4_shr5_i_i381 = ((local_bb4_or4_i_i380 & 32'h7FFFFFF) >> 32'h8);

// This section implements a registered operation.
// 
wire SFC_3_VALID_222_223_0_inputs_ready;
 reg SFC_3_VALID_222_223_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_222_223_0_stall_in;
wire SFC_3_VALID_222_223_0_output_regs_ready;
 reg SFC_3_VALID_222_223_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_222_223_0_causedstall;

assign SFC_3_VALID_222_223_0_inputs_ready = 1'b1;
assign SFC_3_VALID_222_223_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_221_222_0_stall_in = 1'b0;
assign SFC_3_VALID_222_223_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_222_223_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_222_223_0_output_regs_ready)
		begin
			SFC_3_VALID_222_223_0_NO_SHIFT_REG <= SFC_3_VALID_221_222_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i382_stall_local;
wire [31:0] local_bb4_or6_i_i382;

assign local_bb4_or6_i_i382 = ((local_bb4_shr5_i_i381 & 32'h7FFFF) | (local_bb4_or4_i_i380 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_223_224_0_inputs_ready;
 reg SFC_3_VALID_223_224_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_223_224_0_stall_in;
wire SFC_3_VALID_223_224_0_output_regs_ready;
 reg SFC_3_VALID_223_224_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_223_224_0_causedstall;

assign SFC_3_VALID_223_224_0_inputs_ready = 1'b1;
assign SFC_3_VALID_223_224_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_222_223_0_stall_in = 1'b0;
assign SFC_3_VALID_223_224_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_223_224_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_223_224_0_output_regs_ready)
		begin
			SFC_3_VALID_223_224_0_NO_SHIFT_REG <= SFC_3_VALID_222_223_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i383_stall_local;
wire [31:0] local_bb4_shr7_i_i383;

assign local_bb4_shr7_i_i383 = ((local_bb4_or6_i_i382 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i384_stall_local;
wire [31:0] local_bb4_or6_masked_i_i384;

assign local_bb4_or6_masked_i_i384 = ((local_bb4_or6_i_i382 & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_224_225_0_inputs_ready;
 reg SFC_3_VALID_224_225_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_224_225_0_stall_in;
wire SFC_3_VALID_224_225_0_output_regs_ready;
 reg SFC_3_VALID_224_225_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_224_225_0_causedstall;

assign SFC_3_VALID_224_225_0_inputs_ready = 1'b1;
assign SFC_3_VALID_224_225_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_223_224_0_stall_in = 1'b0;
assign SFC_3_VALID_224_225_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_224_225_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_224_225_0_output_regs_ready)
		begin
			SFC_3_VALID_224_225_0_NO_SHIFT_REG <= SFC_3_VALID_223_224_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i385_stall_local;
wire [31:0] local_bb4_neg_i_i385;

assign local_bb4_neg_i_i385 = ((local_bb4_or6_masked_i_i384 & 32'h7FFFFFF) | (local_bb4_shr7_i_i383 & 32'h7FF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_225_226_0_inputs_ready;
 reg SFC_3_VALID_225_226_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_225_226_0_stall_in;
wire SFC_3_VALID_225_226_0_output_regs_ready;
 reg SFC_3_VALID_225_226_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_225_226_0_causedstall;

assign SFC_3_VALID_225_226_0_inputs_ready = 1'b1;
assign SFC_3_VALID_225_226_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_224_225_0_stall_in = 1'b0;
assign SFC_3_VALID_225_226_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_225_226_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_225_226_0_output_regs_ready)
		begin
			SFC_3_VALID_225_226_0_NO_SHIFT_REG <= SFC_3_VALID_224_225_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i386_stall_local;
wire [31:0] local_bb4_and_i_i386;

assign local_bb4_and_i_i386 = ((local_bb4_neg_i_i385 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_226_227_0_inputs_ready;
 reg SFC_3_VALID_226_227_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_226_227_0_stall_in;
wire SFC_3_VALID_226_227_0_output_regs_ready;
 reg SFC_3_VALID_226_227_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_226_227_0_causedstall;

assign SFC_3_VALID_226_227_0_inputs_ready = 1'b1;
assign SFC_3_VALID_226_227_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_225_226_0_stall_in = 1'b0;
assign SFC_3_VALID_226_227_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_226_227_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_226_227_0_output_regs_ready)
		begin
			SFC_3_VALID_226_227_0_NO_SHIFT_REG <= SFC_3_VALID_225_226_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i386_valid_out;
wire local_bb4__and_i_i386_stall_in;
wire local_bb4__and_i_i386_inputs_ready;
wire local_bb4__and_i_i386_stall_local;
wire [31:0] local_bb4__and_i_i386;

thirtysix_six_comp local_bb4__and_i_i386_popcnt_instance (
	.data((local_bb4_and_i_i386 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i386)
);


assign local_bb4__and_i_i386_inputs_ready = rnode_180to181_bb4_add193_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i386_valid_out = 1'b1;
assign rnode_180to181_bb4_add193_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_227_228_0_inputs_ready;
 reg SFC_3_VALID_227_228_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_227_228_0_stall_in;
wire SFC_3_VALID_227_228_0_output_regs_ready;
 reg SFC_3_VALID_227_228_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_227_228_0_causedstall;

assign SFC_3_VALID_227_228_0_inputs_ready = 1'b1;
assign SFC_3_VALID_227_228_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_226_227_0_stall_in = 1'b0;
assign SFC_3_VALID_227_228_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_227_228_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_227_228_0_output_regs_ready)
		begin
			SFC_3_VALID_227_228_0_NO_SHIFT_REG <= SFC_3_VALID_226_227_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb4__and_i_i386_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i386_0_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i386_1_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i386_2_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb4__and_i_i386_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb4__and_i_i386_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb4__and_i_i386_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb4__and_i_i386_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb4__and_i_i386_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb4__and_i_i386_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb4__and_i_i386_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i386 & 32'h3F)),
	.data_out(rnode_181to182_bb4__and_i_i386_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb4__and_i_i386_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb4__and_i_i386_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb4__and_i_i386_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb4__and_i_i386_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb4__and_i_i386_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i386_stall_in = 1'b0;
assign rnode_181to182_bb4__and_i_i386_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i386_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4__and_i_i386_0_NO_SHIFT_REG = rnode_181to182_bb4__and_i_i386_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4__and_i_i386_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4__and_i_i386_1_NO_SHIFT_REG = rnode_181to182_bb4__and_i_i386_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb4__and_i_i386_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb4__and_i_i386_2_NO_SHIFT_REG = rnode_181to182_bb4__and_i_i386_0_reg_182_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_228_229_0_inputs_ready;
 reg SFC_3_VALID_228_229_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_228_229_0_stall_in;
wire SFC_3_VALID_228_229_0_output_regs_ready;
 reg SFC_3_VALID_228_229_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_228_229_0_causedstall;

assign SFC_3_VALID_228_229_0_inputs_ready = 1'b1;
assign SFC_3_VALID_228_229_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_227_228_0_stall_in = 1'b0;
assign SFC_3_VALID_228_229_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_228_229_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_228_229_0_output_regs_ready)
		begin
			SFC_3_VALID_228_229_0_NO_SHIFT_REG <= SFC_3_VALID_227_228_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i387_stall_local;
wire [31:0] local_bb4_and9_i_i387;

assign local_bb4_and9_i_i387 = ((rnode_181to182_bb4__and_i_i386_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and204_i_stall_local;
wire [31:0] local_bb4_and204_i;

assign local_bb4_and204_i = ((rnode_181to182_bb4__and_i_i386_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and207_i_stall_local;
wire [31:0] local_bb4_and207_i;

assign local_bb4_and207_i = ((rnode_181to182_bb4__and_i_i386_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements a registered operation.
// 
wire SFC_3_VALID_229_230_0_inputs_ready;
 reg SFC_3_VALID_229_230_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_229_230_0_stall_in_0;
 reg SFC_3_VALID_229_230_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_229_230_0_stall_in_1;
wire SFC_3_VALID_229_230_0_output_regs_ready;
 reg SFC_3_VALID_229_230_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_229_230_0_causedstall;

assign SFC_3_VALID_229_230_0_inputs_ready = 1'b1;
assign SFC_3_VALID_229_230_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_228_229_0_stall_in = 1'b0;
assign SFC_3_VALID_229_230_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_229_230_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_229_230_0_output_regs_ready)
		begin
			SFC_3_VALID_229_230_0_NO_SHIFT_REG <= SFC_3_VALID_228_229_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_sub240_i_stall_local;
wire [31:0] local_bb4_sub240_i;

assign local_bb4_sub240_i = (32'h0 - (local_bb4_and9_i_i387 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl205_i_stall_local;
wire [31:0] local_bb4_shl205_i;

assign local_bb4_shl205_i = ((rnode_181to182_bb4_and194_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and204_i & 32'h18));

// This section implements a registered operation.
// 
wire SFC_3_VALID_230_231_0_inputs_ready;
 reg SFC_3_VALID_230_231_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_230_231_0_stall_in;
wire SFC_3_VALID_230_231_0_output_regs_ready;
 reg SFC_3_VALID_230_231_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_230_231_0_causedstall;

assign SFC_3_VALID_230_231_0_inputs_ready = 1'b1;
assign SFC_3_VALID_230_231_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_229_230_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_230_231_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_230_231_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_230_231_0_output_regs_ready)
		begin
			SFC_3_VALID_230_231_0_NO_SHIFT_REG <= SFC_3_VALID_229_230_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_sum_321_pop9_c1_ene5_valid_out;
wire local_bb4_sum_321_pop9_c1_ene5_stall_in;
wire local_bb4_sum_321_pop9_c1_ene5_inputs_ready;
wire local_bb4_sum_321_pop9_c1_ene5_stall_local;
wire [31:0] local_bb4_sum_321_pop9_c1_ene5;
wire local_bb4_sum_321_pop9_c1_ene5_fu_valid_out;
wire local_bb4_sum_321_pop9_c1_ene5_fu_stall_out;

acl_pop local_bb4_sum_321_pop9_c1_ene5_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_229to230_bb4_c1_ene4_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_229to230_bb4_c1_ene5_0_NO_SHIFT_REG),
	.stall_out(local_bb4_sum_321_pop9_c1_ene5_fu_stall_out),
	.valid_in(SFC_3_VALID_229_230_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sum_321_pop9_c1_ene5_fu_valid_out),
	.stall_in(local_bb4_sum_321_pop9_c1_ene5_stall_local),
	.data_out(local_bb4_sum_321_pop9_c1_ene5),
	.feedback_in(feedback_data_in_9),
	.feedback_valid_in(feedback_valid_in_9),
	.feedback_stall_out(feedback_stall_out_9)
);

defparam local_bb4_sum_321_pop9_c1_ene5_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_sum_321_pop9_c1_ene5_feedback.DATA_WIDTH = 32;
defparam local_bb4_sum_321_pop9_c1_ene5_feedback.STYLE = "REGULAR";

assign local_bb4_sum_321_pop9_c1_ene5_inputs_ready = (SFC_3_VALID_229_230_0_valid_out_1_NO_SHIFT_REG & rnode_229to230_bb4_c1_ene4_0_valid_out_0_NO_SHIFT_REG & rnode_229to230_bb4_c1_ene5_0_valid_out_NO_SHIFT_REG);
assign local_bb4_sum_321_pop9_c1_ene5_stall_local = 1'b0;
assign local_bb4_sum_321_pop9_c1_ene5_valid_out = 1'b1;
assign SFC_3_VALID_229_230_0_stall_in_1 = 1'b0;
assign rnode_229to230_bb4_c1_ene4_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cond245_i_stall_local;
wire [31:0] local_bb4_cond245_i;

assign local_bb4_cond245_i = (rnode_180to182_bb4_cmp38_i_2_NO_SHIFT_REG ? local_bb4_sub240_i : (local_bb4__43_i392 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i388_stall_local;
wire [31:0] local_bb4_and206_i388;

assign local_bb4_and206_i388 = (local_bb4_shl205_i & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_231_232_0_inputs_ready;
 reg SFC_3_VALID_231_232_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_231_232_0_stall_in;
wire SFC_3_VALID_231_232_0_output_regs_ready;
 reg SFC_3_VALID_231_232_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_231_232_0_causedstall;

assign SFC_3_VALID_231_232_0_inputs_ready = 1'b1;
assign SFC_3_VALID_231_232_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_230_231_0_stall_in = 1'b0;
assign SFC_3_VALID_231_232_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_231_232_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_231_232_0_output_regs_ready)
		begin
			SFC_3_VALID_231_232_0_NO_SHIFT_REG <= SFC_3_VALID_230_231_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_sum_321_pop9_c1_ene5_1_NO_SHIFT_REG;
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_valid_out_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_in_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_in_0_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_valid_out_0_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in(local_bb4_sum_321_pop9_c1_ene5),
	.data_out(rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_fifo.DATA_WIDTH = 32;
defparam rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_sum_321_pop9_c1_ene5_stall_in = 1'b0;
assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_in_0_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG = rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_1_NO_SHIFT_REG = rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_reg_231_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add246_i_stall_local;
wire [31:0] local_bb4_add246_i;

assign local_bb4_add246_i = (local_bb4_cond245_i + (rnode_180to182_bb4_and17_i327_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i397_stall_local;
wire [31:0] local_bb4_fold_i397;

assign local_bb4_fold_i397 = (local_bb4_cond245_i + (rnode_180to182_bb4_shr16_i326_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl208_i_stall_local;
wire [31:0] local_bb4_shl208_i;

assign local_bb4_shl208_i = ((local_bb4_and206_i388 & 32'h7FFFFFF) << (local_bb4_and207_i & 32'h7));

// This section implements a registered operation.
// 
wire SFC_3_VALID_232_233_0_inputs_ready;
 reg SFC_3_VALID_232_233_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_232_233_0_stall_in;
wire SFC_3_VALID_232_233_0_output_regs_ready;
 reg SFC_3_VALID_232_233_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_232_233_0_causedstall;

assign SFC_3_VALID_232_233_0_inputs_ready = 1'b1;
assign SFC_3_VALID_232_233_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_231_232_0_stall_in = 1'b0;
assign SFC_3_VALID_232_233_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_232_233_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_232_233_0_output_regs_ready)
		begin
			SFC_3_VALID_232_233_0_NO_SHIFT_REG <= SFC_3_VALID_231_232_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u45_stall_local;
wire [31:0] local_bb4_var__u45;

assign local_bb4_var__u45 = rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_valid_out_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_232_NO_SHIFT_REG;

acl_data_fifo rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_232_NO_SHIFT_REG),
	.valid_out(rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_valid_out_reg_232_NO_SHIFT_REG),
	.stall_out(rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_232_NO_SHIFT_REG),
	.data_in(rnode_230to231_bb4_sum_321_pop9_c1_ene5_1_NO_SHIFT_REG),
	.data_out(rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_NO_SHIFT_REG)
);

defparam rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_fifo.DEPTH = 1;
defparam rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_fifo.DATA_WIDTH = 32;
defparam rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_fifo.IMPL = "shift_reg";

assign rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG = rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_reg_232_NO_SHIFT_REG;
assign rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_232_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and251_i_stall_local;
wire [31:0] local_bb4_and251_i;

assign local_bb4_and251_i = (local_bb4_fold_i397 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i402_stall_local;
wire [31:0] local_bb4_and270_i402;

assign local_bb4_and270_i402 = (local_bb4_fold_i397 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and209_i_stall_local;
wire [31:0] local_bb4_and209_i;

assign local_bb4_and209_i = (local_bb4_shl208_i & 32'h7FFFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_233_234_0_inputs_ready;
 reg SFC_3_VALID_233_234_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_233_234_0_stall_in;
wire SFC_3_VALID_233_234_0_output_regs_ready;
 reg SFC_3_VALID_233_234_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_233_234_0_causedstall;

assign SFC_3_VALID_233_234_0_inputs_ready = 1'b1;
assign SFC_3_VALID_233_234_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_232_233_0_stall_in = 1'b0;
assign SFC_3_VALID_233_234_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_233_234_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_233_234_0_output_regs_ready)
		begin
			SFC_3_VALID_233_234_0_NO_SHIFT_REG <= SFC_3_VALID_232_233_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and2_i2_stall_local;
wire [31:0] local_bb4_and2_i2;

assign local_bb4_and2_i2 = (local_bb4_var__u45 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i_stall_local;
wire [31:0] local_bb4_and12_i;

assign local_bb4_and12_i = (local_bb4_var__u45 & 32'hFFFF);

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_NO_SHIFT_REG;
 logic rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_fifo.DEPTH = 5;
defparam rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4_sum_321_pop9_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG = rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_reg_237_NO_SHIFT_REG;
assign rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__44_i393_stall_local;
wire [31:0] local_bb4__44_i393;

assign local_bb4__44_i393 = (local_bb4__40_demorgan_i390 ? (local_bb4_and209_i & 32'h7FFFFFF) : (local_bb4_or220_i & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire SFC_3_VALID_234_235_0_inputs_ready;
 reg SFC_3_VALID_234_235_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_234_235_0_stall_in_0;
 reg SFC_3_VALID_234_235_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_234_235_0_stall_in_1;
wire SFC_3_VALID_234_235_0_output_regs_ready;
 reg SFC_3_VALID_234_235_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_234_235_0_causedstall;

assign SFC_3_VALID_234_235_0_inputs_ready = 1'b1;
assign SFC_3_VALID_234_235_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_233_234_0_stall_in = 1'b0;
assign SFC_3_VALID_234_235_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_234_235_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_234_235_0_output_regs_ready)
		begin
			SFC_3_VALID_234_235_0_NO_SHIFT_REG <= SFC_3_VALID_233_234_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_stall_local;
wire [31:0] local_bb4_shr3_i;

assign local_bb4_shr3_i = ((local_bb4_and2_i2 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_fifo.DATA_WIDTH = 32;
defparam rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_232to237_bb4_sum_321_pop9_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG = rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and251_i_valid_out;
wire local_bb4_and251_i_stall_in;
wire local_bb4_and270_i402_valid_out;
wire local_bb4_and270_i402_stall_in;
wire local_bb4_add246_i_valid_out;
wire local_bb4_add246_i_stall_in;
wire local_bb4__45_i394_valid_out;
wire local_bb4__45_i394_stall_in;
wire local_bb4_not_cmp38_i_valid_out_1;
wire local_bb4_not_cmp38_i_stall_in_1;
wire local_bb4__45_i394_inputs_ready;
wire local_bb4__45_i394_stall_local;
wire [31:0] local_bb4__45_i394;

assign local_bb4__45_i394_inputs_ready = (rnode_180to182_bb4_shr16_i326_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb4_and17_i327_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb4_cmp38_i_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb4_cmp38_i_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb4_and194_i_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb4_cmp38_i_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_and196_i_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_and194_i_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4_and199_i_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb4_and194_i_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb4__and_i_i386_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb4__and_i_i386_0_valid_out_2_NO_SHIFT_REG & rnode_181to182_bb4__and_i_i386_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i394 = (local_bb4__42_i391 ? (rnode_181to182_bb4_and194_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i393 & 32'h7FFFFFF));
assign local_bb4_and251_i_valid_out = 1'b1;
assign local_bb4_and270_i402_valid_out = 1'b1;
assign local_bb4_add246_i_valid_out = 1'b1;
assign local_bb4__45_i394_valid_out = 1'b1;
assign local_bb4_not_cmp38_i_valid_out_1 = 1'b1;
assign rnode_180to182_bb4_shr16_i326_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_and17_i327_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb4_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and196_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and199_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4_and194_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i386_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i386_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb4__and_i_i386_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_235_236_0_inputs_ready;
 reg SFC_3_VALID_235_236_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_235_236_0_stall_in;
wire SFC_3_VALID_235_236_0_output_regs_ready;
 reg SFC_3_VALID_235_236_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_235_236_0_causedstall;

assign SFC_3_VALID_235_236_0_inputs_ready = 1'b1;
assign SFC_3_VALID_235_236_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_234_235_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_235_236_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_235_236_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_235_236_0_output_regs_ready)
		begin
			SFC_3_VALID_235_236_0_NO_SHIFT_REG <= SFC_3_VALID_234_235_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_t_322_pop8_c1_ene3_valid_out;
wire local_bb4_t_322_pop8_c1_ene3_stall_in;
wire local_bb4_t_322_pop8_c1_ene3_inputs_ready;
wire local_bb4_t_322_pop8_c1_ene3_stall_local;
wire [31:0] local_bb4_t_322_pop8_c1_ene3;
wire local_bb4_t_322_pop8_c1_ene3_fu_valid_out;
wire local_bb4_t_322_pop8_c1_ene3_fu_stall_out;

acl_pop local_bb4_t_322_pop8_c1_ene3_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_234to235_bb4_c1_ene4_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_234to235_bb4_c1_ene3_0_NO_SHIFT_REG),
	.stall_out(local_bb4_t_322_pop8_c1_ene3_fu_stall_out),
	.valid_in(SFC_3_VALID_234_235_0_NO_SHIFT_REG),
	.valid_out(local_bb4_t_322_pop8_c1_ene3_fu_valid_out),
	.stall_in(local_bb4_t_322_pop8_c1_ene3_stall_local),
	.data_out(local_bb4_t_322_pop8_c1_ene3),
	.feedback_in(feedback_data_in_8),
	.feedback_valid_in(feedback_valid_in_8),
	.feedback_stall_out(feedback_stall_out_8)
);

defparam local_bb4_t_322_pop8_c1_ene3_feedback.COALESCE_DISTANCE = 1;
defparam local_bb4_t_322_pop8_c1_ene3_feedback.DATA_WIDTH = 32;
defparam local_bb4_t_322_pop8_c1_ene3_feedback.STYLE = "REGULAR";

assign local_bb4_t_322_pop8_c1_ene3_inputs_ready = (SFC_3_VALID_234_235_0_valid_out_1_NO_SHIFT_REG & rnode_234to235_bb4_c1_ene3_0_valid_out_NO_SHIFT_REG & rnode_234to235_bb4_c1_ene4_0_valid_out_NO_SHIFT_REG);
assign local_bb4_t_322_pop8_c1_ene3_stall_local = 1'b0;
assign local_bb4_t_322_pop8_c1_ene3_valid_out = 1'b1;
assign SFC_3_VALID_234_235_0_stall_in_1 = 1'b0;
assign rnode_234to235_bb4_c1_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_c1_ene4_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_and251_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and251_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_and251_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_and251_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_and251_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_and251_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_and251_i_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_and251_i_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_and251_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in((local_bb4_and251_i & 32'hFF)),
	.data_out(rnode_182to183_bb4_and251_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_and251_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_and251_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and251_i_stall_in = 1'b0;
assign rnode_182to183_bb4_and251_i_0_NO_SHIFT_REG = rnode_182to183_bb4_and251_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_and251_i_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and251_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_182to184_bb4_and270_i402_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i402_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and270_i402_0_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i402_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to184_bb4_and270_i402_0_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i402_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i402_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_182to184_bb4_and270_i402_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_182to184_bb4_and270_i402_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to184_bb4_and270_i402_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to184_bb4_and270_i402_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_182to184_bb4_and270_i402_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_182to184_bb4_and270_i402_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_and270_i402 & 32'hFF800000)),
	.data_out(rnode_182to184_bb4_and270_i402_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_182to184_bb4_and270_i402_0_reg_184_fifo.DEPTH = 2;
defparam rnode_182to184_bb4_and270_i402_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_182to184_bb4_and270_i402_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to184_bb4_and270_i402_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_182to184_bb4_and270_i402_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and270_i402_stall_in = 1'b0;
assign rnode_182to184_bb4_and270_i402_0_NO_SHIFT_REG = rnode_182to184_bb4_and270_i402_0_reg_184_NO_SHIFT_REG;
assign rnode_182to184_bb4_and270_i402_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_182to184_bb4_and270_i402_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add246_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add246_i_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_add246_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_add246_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_add246_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_add246_i_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_add246_i_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_add246_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_add246_i),
	.data_out(rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_add246_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_add246_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add246_i_stall_in = 1'b0;
assign rnode_182to183_bb4_add246_i_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add246_i_0_NO_SHIFT_REG = rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4_add246_i_1_NO_SHIFT_REG = rnode_182to183_bb4_add246_i_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4__45_i394_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i394_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i394_1_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i394_2_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb4__45_i394_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4__45_i394_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4__45_i394_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4__45_i394_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4__45_i394_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4__45_i394_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4__45_i394_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in((local_bb4__45_i394 & 32'hFFFFFFF)),
	.data_out(rnode_182to183_bb4__45_i394_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4__45_i394_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4__45_i394_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb4__45_i394_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4__45_i394_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4__45_i394_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i394_stall_in = 1'b0;
assign rnode_182to183_bb4__45_i394_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4__45_i394_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__45_i394_0_NO_SHIFT_REG = rnode_182to183_bb4__45_i394_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4__45_i394_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__45_i394_1_NO_SHIFT_REG = rnode_182to183_bb4__45_i394_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4__45_i394_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb4__45_i394_2_NO_SHIFT_REG = rnode_182to183_bb4__45_i394_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb4_not_cmp38_i_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb4_not_cmp38_i_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb4_not_cmp38_i_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb4_not_cmp38_i_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb4_not_cmp38_i_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp38_i),
	.data_out(rnode_182to183_bb4_not_cmp38_i_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb4_not_cmp38_i_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb4_not_cmp38_i_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp38_i_stall_in_1 = 1'b0;
assign rnode_182to183_bb4_not_cmp38_i_0_NO_SHIFT_REG = rnode_182to183_bb4_not_cmp38_i_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb4_not_cmp38_i_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_236_237_0_inputs_ready;
 reg SFC_3_VALID_236_237_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_236_237_0_stall_in;
wire SFC_3_VALID_236_237_0_output_regs_ready;
 reg SFC_3_VALID_236_237_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_236_237_0_causedstall;

assign SFC_3_VALID_236_237_0_inputs_ready = 1'b1;
assign SFC_3_VALID_236_237_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_235_236_0_stall_in = 1'b0;
assign SFC_3_VALID_236_237_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_236_237_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_236_237_0_output_regs_ready)
		begin
			SFC_3_VALID_236_237_0_NO_SHIFT_REG <= SFC_3_VALID_235_236_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_t_322_pop8_c1_ene3_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_valid_out_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_in_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_in_0_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_235to236_bb4_t_322_pop8_c1_ene3_0_valid_out_0_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in(local_bb4_t_322_pop8_c1_ene3),
	.data_out(rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_fifo.DEPTH = 1;
defparam rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_t_322_pop8_c1_ene3_stall_in = 1'b0;
assign rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_in_0_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_t_322_pop8_c1_ene3_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG = rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_t_322_pop8_c1_ene3_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_t_322_pop8_c1_ene3_1_NO_SHIFT_REG = rnode_235to236_bb4_t_322_pop8_c1_ene3_0_reg_236_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i399_stall_local;
wire local_bb4_notrhs_i399;

assign local_bb4_notrhs_i399 = ((rnode_182to183_bb4_and251_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl274_i_stall_local;
wire [31:0] local_bb4_shl274_i;

assign local_bb4_shl274_i = ((rnode_182to184_bb4_and270_i402_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and248_i_stall_local;
wire [31:0] local_bb4_and248_i;

assign local_bb4_and248_i = (rnode_182to183_bb4_add246_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp259_i_stall_local;
wire local_bb4_cmp259_i;

assign local_bb4_cmp259_i = ($signed(rnode_182to183_bb4_add246_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and226_i_stall_local;
wire [31:0] local_bb4_and226_i;

assign local_bb4_and226_i = ((rnode_182to183_bb4__45_i394_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and271_i_stall_local;
wire [31:0] local_bb4_and271_i;

assign local_bb4_and271_i = ((rnode_182to183_bb4__45_i394_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr272_i_valid_out;
wire local_bb4_shr272_i_stall_in;
wire local_bb4_shr272_i_inputs_ready;
wire local_bb4_shr272_i_stall_local;
wire [31:0] local_bb4_shr272_i;

assign local_bb4_shr272_i_inputs_ready = rnode_182to183_bb4__45_i394_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr272_i = ((rnode_182to183_bb4__45_i394_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr272_i_valid_out = 1'b1;
assign rnode_182to183_bb4__45_i394_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_237_238_0_inputs_ready;
 reg SFC_3_VALID_237_238_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_237_238_0_stall_in;
wire SFC_3_VALID_237_238_0_output_regs_ready;
 reg SFC_3_VALID_237_238_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_237_238_0_causedstall;

assign SFC_3_VALID_237_238_0_inputs_ready = 1'b1;
assign SFC_3_VALID_237_238_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_236_237_0_stall_in = 1'b0;
assign SFC_3_VALID_237_238_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_237_238_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_237_238_0_output_regs_ready)
		begin
			SFC_3_VALID_237_238_0_NO_SHIFT_REG <= SFC_3_VALID_236_237_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_var__u46_stall_local;
wire [31:0] local_bb4_var__u46;

assign local_bb4_var__u46 = rnode_235to236_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_t_322_pop8_c1_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_236to237_bb4_t_322_pop8_c1_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_t_322_pop8_c1_ene3_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_t_322_pop8_c1_ene3_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(rnode_235to236_bb4_t_322_pop8_c1_ene3_1_NO_SHIFT_REG),
	.data_out(rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG = rnode_236to237_bb4_t_322_pop8_c1_ene3_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_t_322_pop8_c1_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i398_stall_local;
wire local_bb4_notlhs_i398;

assign local_bb4_notlhs_i398 = ((local_bb4_and248_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp227_i_stall_local;
wire local_bb4_cmp227_i;

assign local_bb4_cmp227_i = ((local_bb4_and226_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp297_i_stall_local;
wire local_bb4_cmp297_i;

assign local_bb4_cmp297_i = ((local_bb4_and271_i & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp297_i_valid_out;
wire local_bb4_cmp297_i_stall_in;
wire local_bb4_cmp300_i_valid_out;
wire local_bb4_cmp300_i_stall_in;
wire local_bb4_cmp300_i_inputs_ready;
wire local_bb4_cmp300_i_stall_local;
wire local_bb4_cmp300_i;

assign local_bb4_cmp300_i_inputs_ready = rnode_182to183_bb4__45_i394_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp300_i = ((local_bb4_and271_i & 32'h7) == 32'h4);
assign local_bb4_cmp297_i_valid_out = 1'b1;
assign local_bb4_cmp300_i_valid_out = 1'b1;
assign rnode_182to183_bb4__45_i394_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_shr272_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_shr272_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_shr272_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_shr272_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_shr272_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_shr272_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_shr272_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_shr272_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_shr272_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_shr272_i & 32'h1FFFFFF)),
	.data_out(rnode_183to184_bb4_shr272_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_shr272_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_shr272_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr272_i_stall_in = 1'b0;
assign rnode_183to184_bb4_shr272_i_0_NO_SHIFT_REG = rnode_183to184_bb4_shr272_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_shr272_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_shr272_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_3_VALID_238_239_0_inputs_ready;
 reg SFC_3_VALID_238_239_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_238_239_0_stall_in_0;
 reg SFC_3_VALID_238_239_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_238_239_0_stall_in_1;
wire SFC_3_VALID_238_239_0_output_regs_ready;
 reg SFC_3_VALID_238_239_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_238_239_0_causedstall;

assign SFC_3_VALID_238_239_0_inputs_ready = 1'b1;
assign SFC_3_VALID_238_239_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_237_238_0_stall_in = 1'b0;
assign SFC_3_VALID_238_239_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_238_239_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_238_239_0_output_regs_ready)
		begin
			SFC_3_VALID_238_239_0_NO_SHIFT_REG <= SFC_3_VALID_237_238_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and2_i13_stall_local;
wire [31:0] local_bb4_and2_i13;

assign local_bb4_and2_i13 = (local_bb4_var__u46 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and12_i18_stall_local;
wire [31:0] local_bb4_and12_i18;

assign local_bb4_and12_i18 = (local_bb4_var__u46 & 32'hFFFF);

// Register node:
//  * latency = 5
//  * capacity = 5
 logic rnode_237to242_bb4_t_322_pop8_c1_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_237to242_bb4_t_322_pop8_c1_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_237to242_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_NO_SHIFT_REG;
 logic rnode_237to242_bb4_t_322_pop8_c1_ene3_0_valid_out_reg_242_NO_SHIFT_REG;
 logic rnode_237to242_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_242_NO_SHIFT_REG;
 logic rnode_237to242_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to242_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_237to242_bb4_t_322_pop8_c1_ene3_0_valid_out_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_237to242_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in(rnode_236to237_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_fifo.DEPTH = 5;
defparam rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_fifo.DATA_WIDTH = 32;
defparam rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4_t_322_pop8_c1_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to242_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG = rnode_237to242_bb4_t_322_pop8_c1_ene3_0_reg_242_NO_SHIFT_REG;
assign rnode_237to242_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_237to242_bb4_t_322_pop8_c1_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i400_stall_local;
wire local_bb4_not__46_i400;

assign local_bb4_not__46_i400 = (local_bb4_notrhs_i399 | local_bb4_notlhs_i398);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp227_not_i_stall_local;
wire local_bb4_cmp227_not_i;

assign local_bb4_cmp227_not_i = (local_bb4_cmp227_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp297_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_cmp297_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_cmp297_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_cmp297_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_cmp297_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_cmp297_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4_cmp297_i),
	.data_out(rnode_183to184_bb4_cmp297_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_cmp297_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_cmp297_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp297_i_stall_in = 1'b0;
assign rnode_183to184_bb4_cmp297_i_0_NO_SHIFT_REG = rnode_183to184_bb4_cmp297_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_cmp297_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_cmp300_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_cmp300_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_cmp300_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_cmp300_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_cmp300_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_cmp300_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4_cmp300_i),
	.data_out(rnode_183to184_bb4_cmp300_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_cmp300_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_cmp300_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp300_i_stall_in = 1'b0;
assign rnode_183to184_bb4_cmp300_i_0_NO_SHIFT_REG = rnode_183to184_bb4_cmp300_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_cmp300_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and273_i_stall_local;
wire [31:0] local_bb4_and273_i;

assign local_bb4_and273_i = ((rnode_183to184_bb4_shr272_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements a registered operation.
// 
wire SFC_3_VALID_239_240_0_inputs_ready;
 reg SFC_3_VALID_239_240_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_239_240_0_stall_in;
wire SFC_3_VALID_239_240_0_output_regs_ready;
 reg SFC_3_VALID_239_240_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_239_240_0_causedstall;

assign SFC_3_VALID_239_240_0_inputs_ready = 1'b1;
assign SFC_3_VALID_239_240_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_238_239_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_239_240_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_239_240_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_239_240_0_output_regs_ready)
		begin
			SFC_3_VALID_239_240_0_NO_SHIFT_REG <= SFC_3_VALID_238_239_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i14_stall_local;
wire [31:0] local_bb4_shr3_i14;

assign local_bb4_shr3_i14 = ((local_bb4_and2_i13 & 32'hFFFF) & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4_t_322_pop8_c1_ene3_0_valid_out_NO_SHIFT_REG;
 logic rnode_242to243_bb4_t_322_pop8_c1_ene3_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_242to243_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_t_322_pop8_c1_ene3_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4_t_322_pop8_c1_ene3_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4_t_322_pop8_c1_ene3_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(rnode_237to242_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG),
	.data_out(rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_fifo.DATA_WIDTH = 32;
defparam rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_237to242_bb4_t_322_pop8_c1_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG = rnode_242to243_bb4_t_322_pop8_c1_ene3_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_t_322_pop8_c1_ene3_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_t_322_pop8_c1_ene3_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__47_i401_stall_local;
wire local_bb4__47_i401;

assign local_bb4__47_i401 = (local_bb4_cmp227_i | local_bb4_not__46_i400);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i395_stall_local;
wire local_bb4_brmerge12_i395;

assign local_bb4_brmerge12_i395 = (local_bb4_cmp227_not_i | rnode_182to183_bb4_not_cmp38_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot263__i_stall_local;
wire local_bb4_lnot263__i;

assign local_bb4_lnot263__i = (local_bb4_cmp259_i & local_bb4_cmp227_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29749_i_stall_local;
wire [31:0] local_bb4_cmp29749_i;

assign local_bb4_cmp29749_i[31:1] = 31'h0;
assign local_bb4_cmp29749_i[0] = rnode_183to184_bb4_cmp297_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv301_i_stall_local;
wire [31:0] local_bb4_conv301_i;

assign local_bb4_conv301_i[31:1] = 31'h0;
assign local_bb4_conv301_i[0] = rnode_183to184_bb4_cmp300_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i403_stall_local;
wire [31:0] local_bb4_or275_i403;

assign local_bb4_or275_i403 = ((local_bb4_and273_i & 32'h7FFFFF) | (local_bb4_shl274_i & 32'h7F800000));

// This section implements a registered operation.
// 
wire SFC_3_VALID_240_241_0_inputs_ready;
 reg SFC_3_VALID_240_241_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_240_241_0_stall_in;
wire SFC_3_VALID_240_241_0_output_regs_ready;
 reg SFC_3_VALID_240_241_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_240_241_0_causedstall;

assign SFC_3_VALID_240_241_0_inputs_ready = 1'b1;
assign SFC_3_VALID_240_241_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_239_240_0_stall_in = 1'b0;
assign SFC_3_VALID_240_241_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_240_241_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_240_241_0_output_regs_ready)
		begin
			SFC_3_VALID_240_241_0_NO_SHIFT_REG <= SFC_3_VALID_239_240_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i396_stall_local;
wire [31:0] local_bb4_resultSign_0_i396;

assign local_bb4_resultSign_0_i396 = (local_bb4_brmerge12_i395 ? (rnode_182to183_bb4_and35_i336_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i396_valid_out;
wire local_bb4_resultSign_0_i396_stall_in;
wire local_bb4__47_i401_valid_out;
wire local_bb4__47_i401_stall_in;
wire local_bb4_or2672_i_valid_out;
wire local_bb4_or2672_i_stall_in;
wire local_bb4_or2672_i_inputs_ready;
wire local_bb4_or2672_i_stall_local;
wire local_bb4_or2672_i;

assign local_bb4_or2672_i_inputs_ready = (rnode_182to183_bb4_and35_i336_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb4_not_cmp38_i_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb4_add246_i_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb4_and251_i_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb4__45_i394_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb4_add246_i_0_valid_out_1_NO_SHIFT_REG & rnode_182to183_bb4_var__u38_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2672_i = (rnode_182to183_bb4_var__u38_0_NO_SHIFT_REG | local_bb4_lnot263__i);
assign local_bb4_resultSign_0_i396_valid_out = 1'b1;
assign local_bb4__47_i401_valid_out = 1'b1;
assign local_bb4_or2672_i_valid_out = 1'b1;
assign rnode_182to183_bb4_and35_i336_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_not_cmp38_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add246_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_and251_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4__45_i394_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_add246_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb4_var__u38_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_3_VALID_241_242_0_inputs_ready;
 reg SFC_3_VALID_241_242_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_241_242_0_stall_in;
wire SFC_3_VALID_241_242_0_output_regs_ready;
 reg SFC_3_VALID_241_242_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_241_242_0_causedstall;

assign SFC_3_VALID_241_242_0_inputs_ready = 1'b1;
assign SFC_3_VALID_241_242_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_240_241_0_stall_in = 1'b0;
assign SFC_3_VALID_241_242_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_241_242_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_241_242_0_output_regs_ready)
		begin
			SFC_3_VALID_241_242_0_NO_SHIFT_REG <= SFC_3_VALID_240_241_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_resultSign_0_i396_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i396_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_resultSign_0_i396_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i396_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb4_resultSign_0_i396_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i396_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i396_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_resultSign_0_i396_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_resultSign_0_i396_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_resultSign_0_i396_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_resultSign_0_i396_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_resultSign_0_i396_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_resultSign_0_i396_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i396 & 32'h80000000)),
	.data_out(rnode_183to184_bb4_resultSign_0_i396_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_resultSign_0_i396_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_resultSign_0_i396_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb4_resultSign_0_i396_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_resultSign_0_i396_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_resultSign_0_i396_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i396_stall_in = 1'b0;
assign rnode_183to184_bb4_resultSign_0_i396_0_NO_SHIFT_REG = rnode_183to184_bb4_resultSign_0_i396_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_resultSign_0_i396_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_resultSign_0_i396_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4__47_i401_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4__47_i401_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4__47_i401_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4__47_i401_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4__47_i401_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4__47_i401_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4__47_i401_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4__47_i401),
	.data_out(rnode_183to184_bb4__47_i401_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4__47_i401_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4__47_i401_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4__47_i401_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4__47_i401_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4__47_i401_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i401_stall_in = 1'b0;
assign rnode_183to184_bb4__47_i401_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__47_i401_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__47_i401_0_NO_SHIFT_REG = rnode_183to184_bb4__47_i401_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4__47_i401_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4__47_i401_1_NO_SHIFT_REG = rnode_183to184_bb4__47_i401_0_reg_184_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_1_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_2_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_valid_out_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_in_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb4_or2672_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb4_or2672_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb4_or2672_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb4_or2672_i_0_stall_in_0_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb4_or2672_i_0_valid_out_0_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb4_or2672_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb4_or2672_i),
	.data_out(rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.DATA_WIDTH = 1;
defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb4_or2672_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb4_or2672_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2672_i_stall_in = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_0_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_or2672_i_0_NO_SHIFT_REG = rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_or2672_i_1_NO_SHIFT_REG = rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_183to184_bb4_or2672_i_2_NO_SHIFT_REG = rnode_183to184_bb4_or2672_i_0_reg_184_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_242_243_0_inputs_ready;
 reg SFC_3_VALID_242_243_0_valid_out_NO_SHIFT_REG;
wire SFC_3_VALID_242_243_0_stall_in;
wire SFC_3_VALID_242_243_0_output_regs_ready;
 reg SFC_3_VALID_242_243_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_242_243_0_causedstall;

assign SFC_3_VALID_242_243_0_inputs_ready = 1'b1;
assign SFC_3_VALID_242_243_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_241_242_0_stall_in = 1'b0;
assign SFC_3_VALID_242_243_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_242_243_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_242_243_0_output_regs_ready)
		begin
			SFC_3_VALID_242_243_0_NO_SHIFT_REG <= SFC_3_VALID_241_242_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_or276_i_stall_local;
wire [31:0] local_bb4_or276_i;

assign local_bb4_or276_i = ((local_bb4_or275_i403 & 32'h7FFFFFFF) | (rnode_183to184_bb4_resultSign_0_i396_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u47_stall_local;
wire [31:0] local_bb4_var__u47;

assign local_bb4_var__u47[31:1] = 31'h0;
assign local_bb4_var__u47[0] = rnode_183to184_bb4__47_i401_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2814_i_stall_local;
wire local_bb4_or2814_i;

assign local_bb4_or2814_i = (rnode_183to184_bb4__47_i401_0_NO_SHIFT_REG | rnode_183to184_bb4_or2672_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2885_i_stall_local;
wire local_bb4_or2885_i;

assign local_bb4_or2885_i = (rnode_183to184_bb4_or2672_i_1_NO_SHIFT_REG | rnode_183to184_bb4__26_i349_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u48_stall_local;
wire [31:0] local_bb4_var__u48;

assign local_bb4_var__u48[31:1] = 31'h0;
assign local_bb4_var__u48[0] = rnode_183to184_bb4_or2672_i_2_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire SFC_3_VALID_243_244_0_inputs_ready;
 reg SFC_3_VALID_243_244_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_243_244_0_stall_in_0;
 reg SFC_3_VALID_243_244_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_243_244_0_stall_in_1;
wire SFC_3_VALID_243_244_0_output_regs_ready;
 reg SFC_3_VALID_243_244_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_243_244_0_causedstall;

assign SFC_3_VALID_243_244_0_inputs_ready = 1'b1;
assign SFC_3_VALID_243_244_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_242_243_0_stall_in = 1'b0;
assign SFC_3_VALID_243_244_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_243_244_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_243_244_0_output_regs_ready)
		begin
			SFC_3_VALID_243_244_0_NO_SHIFT_REG <= SFC_3_VALID_242_243_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext315_i_stall_local;
wire [31:0] local_bb4_lnot_ext315_i;

assign local_bb4_lnot_ext315_i = ((local_bb4_var__u47 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond283_i_stall_local;
wire [31:0] local_bb4_cond283_i;

assign local_bb4_cond283_i = (local_bb4_or2814_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond290_i_stall_local;
wire [31:0] local_bb4_cond290_i;

assign local_bb4_cond290_i = (local_bb4_or2885_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext311_i_stall_local;
wire [31:0] local_bb4_lnot_ext311_i;

assign local_bb4_lnot_ext311_i = ((local_bb4_var__u48 & 32'h1) ^ 32'h1);

// This section implements a registered operation.
// 
wire SFC_3_VALID_244_245_0_inputs_ready;
 reg SFC_3_VALID_244_245_0_valid_out_0_NO_SHIFT_REG;
wire SFC_3_VALID_244_245_0_stall_in_0;
 reg SFC_3_VALID_244_245_0_valid_out_1_NO_SHIFT_REG;
wire SFC_3_VALID_244_245_0_stall_in_1;
 reg SFC_3_VALID_244_245_0_valid_out_2_NO_SHIFT_REG;
wire SFC_3_VALID_244_245_0_stall_in_2;
wire SFC_3_VALID_244_245_0_output_regs_ready;
 reg SFC_3_VALID_244_245_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_3_VALID_244_245_0_causedstall;

assign SFC_3_VALID_244_245_0_inputs_ready = 1'b1;
assign SFC_3_VALID_244_245_0_output_regs_ready = 1'b1;
assign SFC_3_VALID_243_244_0_stall_in_0 = 1'b0;
assign SFC_3_VALID_244_245_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_3_VALID_244_245_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_3_VALID_244_245_0_output_regs_ready)
		begin
			SFC_3_VALID_244_245_0_NO_SHIFT_REG <= SFC_3_VALID_243_244_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and294_i_stall_local;
wire [31:0] local_bb4_and294_i;

assign local_bb4_and294_i = ((local_bb4_cond283_i | 32'h80000000) & local_bb4_or276_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i404_stall_local;
wire [31:0] local_bb4_or295_i404;

assign local_bb4_or295_i404 = ((local_bb4_cond290_i & 32'h7F800000) | (local_bb4_cond293_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i407_stall_local;
wire [31:0] local_bb4_reduction_0_i407;

assign local_bb4_reduction_0_i407 = ((local_bb4_lnot_ext311_i & 32'h1) & (local_bb4_lnot_ext_i406 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and303_i_stall_local;
wire [31:0] local_bb4_and303_i;

assign local_bb4_and303_i = ((local_bb4_conv301_i & 32'h1) & local_bb4_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or296_i_stall_local;
wire [31:0] local_bb4_or296_i;

assign local_bb4_or296_i = ((local_bb4_or295_i404 & 32'h7FC00000) | local_bb4_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i405_stall_local;
wire [31:0] local_bb4_lor_ext_i405;

assign local_bb4_lor_ext_i405 = ((local_bb4_cmp29749_i & 32'h1) | (local_bb4_and303_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i408_stall_local;
wire [31:0] local_bb4_reduction_1_i408;

assign local_bb4_reduction_1_i408 = ((local_bb4_lnot_ext315_i & 32'h1) & (local_bb4_lor_ext_i405 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i409_stall_local;
wire [31:0] local_bb4_reduction_2_i409;

assign local_bb4_reduction_2_i409 = ((local_bb4_reduction_0_i407 & 32'h1) & (local_bb4_reduction_1_i408 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_add321_i_stall_local;
wire [31:0] local_bb4_add321_i;

assign local_bb4_add321_i = ((local_bb4_reduction_2_i409 & 32'h1) + local_bb4_or296_i);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u49_valid_out;
wire local_bb4_var__u49_stall_in;
wire local_bb4_var__u49_inputs_ready;
wire local_bb4_var__u49_stall_local;
wire [31:0] local_bb4_var__u49;

assign local_bb4_var__u49_inputs_ready = (rnode_182to184_bb4_and270_i402_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_resultSign_0_i396_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_or2672_i_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4__26_i349_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4__26_i349_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4__47_i401_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4_or2672_i_0_valid_out_0_NO_SHIFT_REG & rnode_183to184_bb4__26_i349_0_valid_out_2_NO_SHIFT_REG & rnode_183to184_bb4_or2672_i_0_valid_out_2_NO_SHIFT_REG & rnode_183to184_bb4_shr272_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4__47_i401_0_valid_out_1_NO_SHIFT_REG & rnode_183to184_bb4_cmp297_i_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb4_cmp300_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_var__u49 = local_bb4_add321_i;
assign local_bb4_var__u49_valid_out = 1'b1;
assign rnode_182to184_bb4_and270_i402_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_resultSign_0_i396_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i349_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i349_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__47_i401_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__26_i349_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_or2672_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_shr272_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4__47_i401_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp297_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb4_cmp300_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_call_i13__inputs_ready;
 reg local_bb4_call_i13__valid_out_NO_SHIFT_REG;
wire local_bb4_call_i13__stall_in;
wire local_bb4_call_i13__output_regs_ready;
wire [31:0] local_bb4_call_i13_;
 reg local_bb4_call_i13__valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_1_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_2_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_3_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_4_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_5_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_6_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_7_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_8_NO_SHIFT_REG;
 reg local_bb4_call_i13__valid_pipe_9_NO_SHIFT_REG;
wire local_bb4_call_i13__causedstall;

acl_fp_sqrt_s5 fp_module_local_bb4_call_i13_ (
	.clock(clock),
	.dataa(local_bb4_var__u49),
	.enable(local_bb4_call_i13__output_regs_ready),
	.result(local_bb4_call_i13_)
);


assign local_bb4_call_i13__inputs_ready = 1'b1;
assign local_bb4_call_i13__output_regs_ready = 1'b1;
assign local_bb4_var__u49_stall_in = 1'b0;
assign local_bb4_call_i13__causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_call_i13__valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i13__valid_pipe_9_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_call_i13__output_regs_ready)
		begin
			local_bb4_call_i13__valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_call_i13__valid_pipe_1_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_0_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_2_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_1_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_3_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_2_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_4_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_3_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_5_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_4_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_6_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_5_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_7_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_6_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_8_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_7_NO_SHIFT_REG;
			local_bb4_call_i13__valid_pipe_9_NO_SHIFT_REG <= local_bb4_call_i13__valid_pipe_8_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_call_i13__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_call_i13__output_regs_ready)
		begin
			local_bb4_call_i13__valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_call_i13__stall_in))
			begin
				local_bb4_call_i13__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_astype_i_i14_stall_local;
wire [31:0] local_bb4_astype_i_i14;

assign local_bb4_astype_i_i14 = local_bb4_call_i13_;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i15_stall_local;
wire [31:0] local_bb4_and_i_i15;

assign local_bb4_and_i_i15 = (local_bb4_astype_i_i14 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4__op_stall_local;
wire [31:0] local_bb4__op;

assign local_bb4__op = (local_bb4_astype_i_i14 ^ 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i_i16_stall_local;
wire local_bb4_cmp_i_i16;

assign local_bb4_cmp_i_i16 = ((local_bb4_and_i_i15 & 32'h7F800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u50_stall_local;
wire [31:0] local_bb4_var__u50;

assign local_bb4_var__u50 = local_bb4__op;

// This section implements an unregistered operation.
// 
wire local_bb4_cast_after_negation_valid_out;
wire local_bb4_cast_after_negation_stall_in;
wire local_bb4_cast_after_negation_inputs_ready;
wire local_bb4_cast_after_negation_stall_local;
wire [31:0] local_bb4_cast_after_negation;

assign local_bb4_cast_after_negation_inputs_ready = local_bb4_call_i13__valid_out_NO_SHIFT_REG;
assign local_bb4_cast_after_negation = (local_bb4_cmp_i_i16 ? 32'h80000000 : local_bb4_var__u50);
assign local_bb4_cast_after_negation_valid_out = 1'b1;
assign local_bb4_call_i13__stall_in = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_div_inputs_ready;
 reg local_bb4_div_valid_out_NO_SHIFT_REG;
wire local_bb4_div_stall_in;
wire local_bb4_div_output_regs_ready;
wire [31:0] local_bb4_div;
 reg local_bb4_div_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb4_div_valid_pipe_12_NO_SHIFT_REG;
wire local_bb4_div_causedstall;

acl_fp_div_s5 fp_module_local_bb4_div (
	.clock(clock),
	.dataa(local_bb4_cast_after_negation),
	.datab(input_wii_mul48),
	.enable(local_bb4_div_output_regs_ready),
	.result(local_bb4_div)
);


assign local_bb4_div_inputs_ready = 1'b1;
assign local_bb4_div_output_regs_ready = 1'b1;
assign local_bb4_cast_after_negation_stall_in = 1'b0;
assign local_bb4_div_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_div_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb4_div_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_div_output_regs_ready)
		begin
			local_bb4_div_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_div_valid_pipe_1_NO_SHIFT_REG <= local_bb4_div_valid_pipe_0_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_2_NO_SHIFT_REG <= local_bb4_div_valid_pipe_1_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_3_NO_SHIFT_REG <= local_bb4_div_valid_pipe_2_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_4_NO_SHIFT_REG <= local_bb4_div_valid_pipe_3_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_5_NO_SHIFT_REG <= local_bb4_div_valid_pipe_4_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_6_NO_SHIFT_REG <= local_bb4_div_valid_pipe_5_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_7_NO_SHIFT_REG <= local_bb4_div_valid_pipe_6_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_8_NO_SHIFT_REG <= local_bb4_div_valid_pipe_7_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_9_NO_SHIFT_REG <= local_bb4_div_valid_pipe_8_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_10_NO_SHIFT_REG <= local_bb4_div_valid_pipe_9_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_11_NO_SHIFT_REG <= local_bb4_div_valid_pipe_10_NO_SHIFT_REG;
			local_bb4_div_valid_pipe_12_NO_SHIFT_REG <= local_bb4_div_valid_pipe_11_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_div_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_div_output_regs_ready)
		begin
			local_bb4_div_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_div_stall_in))
			begin
				local_bb4_div_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb4_call_i_div_inputs_ready;
 reg local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG;
wire local_bb4_call_i_div_stall_in_0;
 reg local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG;
wire local_bb4_call_i_div_stall_in_1;
wire local_bb4_call_i_div_output_regs_ready;
wire [31:0] local_bb4_call_i_div;
 reg local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG;
 reg local_bb4_call_i_div_valid_pipe_14_NO_SHIFT_REG;
wire local_bb4_call_i_div_causedstall;

acl_fp_exp_s5 fp_module_local_bb4_call_i_div (
	.clock(clock),
	.dataa(local_bb4_div),
	.enable(local_bb4_call_i_div_output_regs_ready),
	.result(local_bb4_call_i_div)
);


assign local_bb4_call_i_div_inputs_ready = 1'b1;
assign local_bb4_call_i_div_output_regs_ready = 1'b1;
assign local_bb4_div_stall_in = 1'b0;
assign local_bb4_call_i_div_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_pipe_14_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_call_i_div_output_regs_ready)
		begin
			local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_0_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_1_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_2_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_3_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_4_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_5_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_6_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_7_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_8_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_9_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_10_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_11_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_12_NO_SHIFT_REG;
			local_bb4_call_i_div_valid_pipe_14_NO_SHIFT_REG <= local_bb4_call_i_div_valid_pipe_13_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_call_i_div_output_regs_ready)
		begin
			local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_call_i_div_stall_in_0))
			begin
				local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_call_i_div_stall_in_1))
			begin
				local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_astype_i_i_stall_local;
wire [31:0] local_bb4_astype_i_i;

assign local_bb4_astype_i_i = local_bb4_call_i_div;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u51_stall_local;
wire [31:0] local_bb4_var__u51;

assign local_bb4_var__u51 = local_bb4_call_i_div;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i_stall_local;
wire [31:0] local_bb4_and_i_i;

assign local_bb4_and_i_i = (local_bb4_astype_i_i & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i_i_stall_local;
wire local_bb4_cmp_i_i;

assign local_bb4_cmp_i_i = ((local_bb4_and_i_i & 32'h7F800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u52_stall_local;
wire [31:0] local_bb4_var__u52;

assign local_bb4_var__u52 = (local_bb4_cmp_i_i ? 32'h0 : local_bb4_var__u51);

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i222_stall_local;
wire [31:0] local_bb4_shr2_i222;

assign local_bb4_shr2_i222 = (local_bb4_var__u52 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i224_stall_local;
wire [31:0] local_bb4_xor_i224;

assign local_bb4_xor_i224 = (local_bb4_var__u52 ^ local_bb4_var__u36);

// This section implements an unregistered operation.
// 
wire local_bb4_and6_i227_stall_local;
wire [31:0] local_bb4_and6_i227;

assign local_bb4_and6_i227 = (local_bb4_var__u52 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and3_i223_stall_local;
wire [31:0] local_bb4_and3_i223;

assign local_bb4_and3_i223 = ((local_bb4_shr2_i222 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_i233_stall_local;
wire local_bb4_lnot17_i233;

assign local_bb4_lnot17_i233 = ((local_bb4_and6_i227 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u53_stall_local;
wire [31:0] local_bb4_var__u53;

assign local_bb4_var__u53 = ((local_bb4_and6_i227 & 32'h7FFFFF) | (local_bb4_and_i221 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_or47_i255_stall_local;
wire [31:0] local_bb4_or47_i255;

assign local_bb4_or47_i255 = ((local_bb4_and6_i227 & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot8_i229_stall_local;
wire local_bb4_lnot8_i229;

assign local_bb4_lnot8_i229 = ((local_bb4_and3_i223 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_i231_stall_local;
wire local_bb4_cmp11_i231;

assign local_bb4_cmp11_i231 = ((local_bb4_and3_i223 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u54_stall_local;
wire [31:0] local_bb4_var__u54;

assign local_bb4_var__u54 = ((local_bb4_and3_i223 & 32'hFF) | (local_bb4_and6_i227 & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i265_stall_local;
wire [31:0] local_bb4_add_i265;

assign local_bb4_add_i265 = ((local_bb4_and3_i223 & 32'hFF) + (local_bb4_and_i221 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_not_i237_stall_local;
wire local_bb4_lnot17_not_i237;

assign local_bb4_lnot17_not_i237 = (local_bb4_lnot17_i233 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u55_stall_local;
wire local_bb4_var__u55;

assign local_bb4_var__u55 = ((local_bb4_var__u53 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_conv1_i_i257_stall_local;
wire [63:0] local_bb4_conv1_i_i257;

assign local_bb4_conv1_i_i257[63:32] = 32'h0;
assign local_bb4_conv1_i_i257[31:0] = ((local_bb4_or47_i255 & 32'hFFFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_not_i238_stall_local;
wire local_bb4_cmp11_not_i238;

assign local_bb4_cmp11_not_i238 = (local_bb4_cmp11_i231 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u56_stall_local;
wire local_bb4_var__u56;

assign local_bb4_var__u56 = ((local_bb4_var__u54 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge3_i239_stall_local;
wire local_bb4_brmerge3_i239;

assign local_bb4_brmerge3_i239 = (local_bb4_var__u56 | local_bb4_cmp11_not_i238);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_i241_stall_local;
wire local_bb4__mux_mux_i241;

assign local_bb4__mux_mux_i241 = (local_bb4_var__u56 | local_bb4_cmp11_i231);

// This section implements an unregistered operation.
// 
wire local_bb4__not_i243_stall_local;
wire local_bb4__not_i243;

assign local_bb4__not_i243 = (local_bb4_var__u56 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge5_i240_stall_local;
wire local_bb4_brmerge5_i240;

assign local_bb4_brmerge5_i240 = (local_bb4_brmerge3_i239 | local_bb4_lnot17_not_i237);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i244_stall_local;
wire local_bb4_reduction_3_i244;

assign local_bb4_reduction_3_i244 = (local_bb4_cmp11_i231 & local_bb4__not_i243);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_mux_i242_stall_local;
wire local_bb4__mux_mux_mux_i242;

assign local_bb4__mux_mux_mux_i242 = (local_bb4_brmerge5_i240 & local_bb4__mux_mux_i241);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i245_stall_local;
wire local_bb4_reduction_5_i245;

assign local_bb4_reduction_5_i245 = (local_bb4_lnot14_i232 & local_bb4_reduction_3_i244);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i224_valid_out;
wire local_bb4_xor_i224_stall_in;
wire local_bb4_lnot14_i232_valid_out_1;
wire local_bb4_lnot14_i232_stall_in_1;
wire local_bb4_lnot_i228_valid_out;
wire local_bb4_lnot_i228_stall_in;
wire local_bb4_cmp_i230_valid_out;
wire local_bb4_cmp_i230_stall_in;
wire local_bb4_add_i265_valid_out;
wire local_bb4_add_i265_stall_in;
wire local_bb4_conv_i_i256_valid_out;
wire local_bb4_conv_i_i256_stall_in;
wire local_bb4_reduction_6_i246_valid_out;
wire local_bb4_reduction_6_i246_stall_in;
wire local_bb4_lnot17_i233_valid_out_1;
wire local_bb4_lnot17_i233_stall_in_1;
wire local_bb4_lnot8_i229_valid_out;
wire local_bb4_lnot8_i229_stall_in;
wire local_bb4_cmp11_i231_valid_out_3;
wire local_bb4_cmp11_i231_stall_in_3;
wire local_bb4_conv1_i_i257_valid_out;
wire local_bb4_conv1_i_i257_stall_in;
wire local_bb4__mux_mux_mux_i242_valid_out;
wire local_bb4__mux_mux_mux_i242_stall_in;
wire local_bb4_reduction_6_i246_inputs_ready;
wire local_bb4_reduction_6_i246_stall_local;
wire local_bb4_reduction_6_i246;

assign local_bb4_reduction_6_i246_inputs_ready = (rnode_224to225_bb4_c1_ene2_0_valid_out_NO_SHIFT_REG & local_bb4_call_i_div_valid_out_1_NO_SHIFT_REG & local_bb4_call_i_div_valid_out_0_NO_SHIFT_REG);
assign local_bb4_reduction_6_i246 = (local_bb4_var__u55 & local_bb4_reduction_5_i245);
assign local_bb4_xor_i224_valid_out = 1'b1;
assign local_bb4_lnot14_i232_valid_out_1 = 1'b1;
assign local_bb4_lnot_i228_valid_out = 1'b1;
assign local_bb4_cmp_i230_valid_out = 1'b1;
assign local_bb4_add_i265_valid_out = 1'b1;
assign local_bb4_conv_i_i256_valid_out = 1'b1;
assign local_bb4_reduction_6_i246_valid_out = 1'b1;
assign local_bb4_lnot17_i233_valid_out_1 = 1'b1;
assign local_bb4_lnot8_i229_valid_out = 1'b1;
assign local_bb4_cmp11_i231_valid_out_3 = 1'b1;
assign local_bb4_conv1_i_i257_valid_out = 1'b1;
assign local_bb4__mux_mux_mux_i242_valid_out = 1'b1;
assign rnode_224to225_bb4_c1_ene2_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_call_i_div_stall_in_1 = 1'b0;
assign local_bb4_call_i_div_stall_in_0 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_225to226_bb4_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_225to226_bb4_xor_i224_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_xor_i224_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_225to226_bb4_xor_i224_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_xor_i224_0_valid_out_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_xor_i224_0_stall_in_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_xor_i224_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_xor_i224_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_xor_i224_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_xor_i224_0_stall_in_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_xor_i224_0_valid_out_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_xor_i224_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i224),
	.data_out(rnode_225to226_bb4_xor_i224_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_xor_i224_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_xor_i224_0_reg_226_fifo.DATA_WIDTH = 32;
defparam rnode_225to226_bb4_xor_i224_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_xor_i224_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_xor_i224_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i224_stall_in = 1'b0;
assign rnode_225to226_bb4_xor_i224_0_NO_SHIFT_REG = rnode_225to226_bb4_xor_i224_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_xor_i224_0_stall_in_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_lnot14_i232_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_valid_out_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_stall_in_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot14_i232_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_lnot14_i232_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_lnot14_i232_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_lnot14_i232_0_stall_in_0_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_lnot14_i232_0_valid_out_0_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_lnot14_i232_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_lnot14_i232),
	.data_out(rnode_225to226_bb4_lnot14_i232_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_lnot14_i232_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_lnot14_i232_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4_lnot14_i232_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_lnot14_i232_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_lnot14_i232_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot14_i232_stall_in_1 = 1'b0;
assign rnode_225to226_bb4_lnot14_i232_0_stall_in_0_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot14_i232_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_lnot14_i232_0_NO_SHIFT_REG = rnode_225to226_bb4_lnot14_i232_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_lnot14_i232_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_lnot14_i232_1_NO_SHIFT_REG = rnode_225to226_bb4_lnot14_i232_0_reg_226_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_lnot_i228_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_valid_out_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_stall_in_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot_i228_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_lnot_i228_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_lnot_i228_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_lnot_i228_0_stall_in_0_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_lnot_i228_0_valid_out_0_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_lnot_i228_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_lnot_i228),
	.data_out(rnode_225to226_bb4_lnot_i228_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_lnot_i228_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_lnot_i228_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4_lnot_i228_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_lnot_i228_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_lnot_i228_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot_i228_stall_in = 1'b0;
assign rnode_225to226_bb4_lnot_i228_0_stall_in_0_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot_i228_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_lnot_i228_0_NO_SHIFT_REG = rnode_225to226_bb4_lnot_i228_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_lnot_i228_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_lnot_i228_1_NO_SHIFT_REG = rnode_225to226_bb4_lnot_i228_0_reg_226_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_cmp_i230_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_2_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_3_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_valid_out_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_stall_in_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp_i230_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_cmp_i230_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_cmp_i230_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_cmp_i230_0_stall_in_0_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_cmp_i230_0_valid_out_0_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_cmp_i230_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_cmp_i230),
	.data_out(rnode_225to226_bb4_cmp_i230_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_cmp_i230_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_cmp_i230_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4_cmp_i230_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_cmp_i230_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_cmp_i230_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp_i230_stall_in = 1'b0;
assign rnode_225to226_bb4_cmp_i230_0_stall_in_0_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp_i230_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_cmp_i230_0_NO_SHIFT_REG = rnode_225to226_bb4_cmp_i230_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_cmp_i230_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_cmp_i230_1_NO_SHIFT_REG = rnode_225to226_bb4_cmp_i230_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_cmp_i230_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_cmp_i230_2_NO_SHIFT_REG = rnode_225to226_bb4_cmp_i230_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_cmp_i230_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_cmp_i230_3_NO_SHIFT_REG = rnode_225to226_bb4_cmp_i230_0_reg_226_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_add_i265_0_valid_out_NO_SHIFT_REG;
 logic rnode_225to226_bb4_add_i265_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_225to226_bb4_add_i265_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_add_i265_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_225to226_bb4_add_i265_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_add_i265_0_valid_out_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_add_i265_0_stall_in_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_add_i265_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_add_i265_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_add_i265_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_add_i265_0_stall_in_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_add_i265_0_valid_out_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_add_i265_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in((local_bb4_add_i265 & 32'h1FF)),
	.data_out(rnode_225to226_bb4_add_i265_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_add_i265_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_add_i265_0_reg_226_fifo.DATA_WIDTH = 32;
defparam rnode_225to226_bb4_add_i265_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_add_i265_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_add_i265_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add_i265_stall_in = 1'b0;
assign rnode_225to226_bb4_add_i265_0_NO_SHIFT_REG = rnode_225to226_bb4_add_i265_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_add_i265_0_stall_in_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_add_i265_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_reduction_6_i246_0_valid_out_NO_SHIFT_REG;
 logic rnode_225to226_bb4_reduction_6_i246_0_stall_in_NO_SHIFT_REG;
 logic rnode_225to226_bb4_reduction_6_i246_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_reduction_6_i246_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4_reduction_6_i246_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_reduction_6_i246_0_valid_out_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_reduction_6_i246_0_stall_in_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_reduction_6_i246_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_reduction_6_i246_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_reduction_6_i246_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_reduction_6_i246_0_stall_in_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_reduction_6_i246_0_valid_out_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_reduction_6_i246_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_6_i246),
	.data_out(rnode_225to226_bb4_reduction_6_i246_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_reduction_6_i246_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_reduction_6_i246_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4_reduction_6_i246_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_reduction_6_i246_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_reduction_6_i246_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_6_i246_stall_in = 1'b0;
assign rnode_225to226_bb4_reduction_6_i246_0_NO_SHIFT_REG = rnode_225to226_bb4_reduction_6_i246_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_reduction_6_i246_0_stall_in_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_reduction_6_i246_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_lnot17_i233_0_valid_out_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot17_i233_0_stall_in_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot17_i233_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot17_i233_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot17_i233_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot17_i233_0_valid_out_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot17_i233_0_stall_in_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot17_i233_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_lnot17_i233_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_lnot17_i233_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_lnot17_i233_0_stall_in_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_lnot17_i233_0_valid_out_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_lnot17_i233_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_lnot17_i233),
	.data_out(rnode_225to226_bb4_lnot17_i233_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_lnot17_i233_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_lnot17_i233_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4_lnot17_i233_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_lnot17_i233_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_lnot17_i233_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot17_i233_stall_in_1 = 1'b0;
assign rnode_225to226_bb4_lnot17_i233_0_NO_SHIFT_REG = rnode_225to226_bb4_lnot17_i233_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_lnot17_i233_0_stall_in_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot17_i233_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_lnot8_i229_0_valid_out_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot8_i229_0_stall_in_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot8_i229_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot8_i229_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot8_i229_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot8_i229_0_valid_out_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot8_i229_0_stall_in_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_lnot8_i229_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_lnot8_i229_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_lnot8_i229_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_lnot8_i229_0_stall_in_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_lnot8_i229_0_valid_out_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_lnot8_i229_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_lnot8_i229),
	.data_out(rnode_225to226_bb4_lnot8_i229_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_lnot8_i229_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_lnot8_i229_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4_lnot8_i229_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_lnot8_i229_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_lnot8_i229_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot8_i229_stall_in = 1'b0;
assign rnode_225to226_bb4_lnot8_i229_0_NO_SHIFT_REG = rnode_225to226_bb4_lnot8_i229_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_lnot8_i229_0_stall_in_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot8_i229_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4_cmp11_i231_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_1_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_2_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_valid_out_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_stall_in_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4_cmp11_i231_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4_cmp11_i231_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4_cmp11_i231_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4_cmp11_i231_0_stall_in_0_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4_cmp11_i231_0_valid_out_0_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4_cmp11_i231_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4_cmp11_i231),
	.data_out(rnode_225to226_bb4_cmp11_i231_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4_cmp11_i231_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4_cmp11_i231_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4_cmp11_i231_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4_cmp11_i231_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4_cmp11_i231_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp11_i231_stall_in_3 = 1'b0;
assign rnode_225to226_bb4_cmp11_i231_0_stall_in_0_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp11_i231_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_cmp11_i231_0_NO_SHIFT_REG = rnode_225to226_bb4_cmp11_i231_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_cmp11_i231_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_cmp11_i231_1_NO_SHIFT_REG = rnode_225to226_bb4_cmp11_i231_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4_cmp11_i231_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_cmp11_i231_2_NO_SHIFT_REG = rnode_225to226_bb4_cmp11_i231_0_reg_226_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_mul_i_i258_inputs_ready;
 reg local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG;
wire local_bb4_mul_i_i258_stall_in_0;
 reg local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i258_stall_in_1;
wire local_bb4_mul_i_i258_output_regs_ready;
wire [63:0] local_bb4_mul_i_i258;
 reg local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul_i_i258_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i258_causedstall;

acl_int_mult int_module_local_bb4_mul_i_i258 (
	.clock(clock),
	.dataa(((local_bb4_conv1_i_i257 & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb4_conv_i_i256 & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb4_mul_i_i258_output_regs_ready),
	.result(local_bb4_mul_i_i258)
);

defparam int_module_local_bb4_mul_i_i258.INPUT1_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i258.INPUT2_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i258.OUTPUT_WIDTH = 64;
defparam int_module_local_bb4_mul_i_i258.LATENCY = 3;
defparam int_module_local_bb4_mul_i_i258.SIGNED = 0;

assign local_bb4_mul_i_i258_inputs_ready = 1'b1;
assign local_bb4_mul_i_i258_output_regs_ready = 1'b1;
assign local_bb4_conv1_i_i257_stall_in = 1'b0;
assign local_bb4_conv_i_i256_stall_in = 1'b0;
assign local_bb4_mul_i_i258_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i258_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i258_output_regs_ready)
		begin
			local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i258_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul_i_i258_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i258_output_regs_ready)
		begin
			local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul_i_i258_stall_in_0))
			begin
				local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_mul_i_i258_stall_in_1))
			begin
				local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_valid_out_NO_SHIFT_REG;
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_stall_in_NO_SHIFT_REG;
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_NO_SHIFT_REG;
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_inputs_ready_NO_SHIFT_REG;
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_valid_out_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_stall_in_reg_226_NO_SHIFT_REG;
 logic rnode_225to226_bb4__mux_mux_mux_i242_0_stall_out_reg_226_NO_SHIFT_REG;

acl_data_fifo rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_225to226_bb4__mux_mux_mux_i242_0_stall_in_reg_226_NO_SHIFT_REG),
	.valid_out(rnode_225to226_bb4__mux_mux_mux_i242_0_valid_out_reg_226_NO_SHIFT_REG),
	.stall_out(rnode_225to226_bb4__mux_mux_mux_i242_0_stall_out_reg_226_NO_SHIFT_REG),
	.data_in(local_bb4__mux_mux_mux_i242),
	.data_out(rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_NO_SHIFT_REG)
);

defparam rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_fifo.DEPTH = 1;
defparam rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_fifo.DATA_WIDTH = 1;
defparam rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_fifo.IMPL = "shift_reg";

assign rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__mux_mux_mux_i242_stall_in = 1'b0;
assign rnode_225to226_bb4__mux_mux_mux_i242_0_NO_SHIFT_REG = rnode_225to226_bb4__mux_mux_mux_i242_0_reg_226_NO_SHIFT_REG;
assign rnode_225to226_bb4__mux_mux_mux_i242_0_stall_in_reg_226_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4__mux_mux_mux_i242_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_226to229_bb4_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_226to229_bb4_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_226to229_bb4_xor_i224_0_NO_SHIFT_REG;
 logic rnode_226to229_bb4_xor_i224_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_226to229_bb4_xor_i224_0_reg_229_NO_SHIFT_REG;
 logic rnode_226to229_bb4_xor_i224_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_226to229_bb4_xor_i224_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_226to229_bb4_xor_i224_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_226to229_bb4_xor_i224_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_226to229_bb4_xor_i224_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_226to229_bb4_xor_i224_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_226to229_bb4_xor_i224_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_226to229_bb4_xor_i224_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in(rnode_225to226_bb4_xor_i224_0_NO_SHIFT_REG),
	.data_out(rnode_226to229_bb4_xor_i224_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_226to229_bb4_xor_i224_0_reg_229_fifo.DEPTH = 3;
defparam rnode_226to229_bb4_xor_i224_0_reg_229_fifo.DATA_WIDTH = 32;
defparam rnode_226to229_bb4_xor_i224_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_226to229_bb4_xor_i224_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_226to229_bb4_xor_i224_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_226to229_bb4_xor_i224_0_NO_SHIFT_REG = rnode_226to229_bb4_xor_i224_0_reg_229_NO_SHIFT_REG;
assign rnode_226to229_bb4_xor_i224_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_226to229_bb4_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_not_i251_stall_local;
wire local_bb4_lnot14_not_i251;

assign local_bb4_lnot14_not_i251 = (rnode_225to226_bb4_lnot14_i232_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_226to227_bb4_add_i265_0_valid_out_NO_SHIFT_REG;
 logic rnode_226to227_bb4_add_i265_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_226to227_bb4_add_i265_0_NO_SHIFT_REG;
 logic rnode_226to227_bb4_add_i265_0_reg_227_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_226to227_bb4_add_i265_0_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_add_i265_0_valid_out_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_add_i265_0_stall_in_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_add_i265_0_stall_out_reg_227_NO_SHIFT_REG;

acl_data_fifo rnode_226to227_bb4_add_i265_0_reg_227_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_226to227_bb4_add_i265_0_reg_227_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_226to227_bb4_add_i265_0_stall_in_reg_227_NO_SHIFT_REG),
	.valid_out(rnode_226to227_bb4_add_i265_0_valid_out_reg_227_NO_SHIFT_REG),
	.stall_out(rnode_226to227_bb4_add_i265_0_stall_out_reg_227_NO_SHIFT_REG),
	.data_in((rnode_225to226_bb4_add_i265_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_226to227_bb4_add_i265_0_reg_227_NO_SHIFT_REG)
);

defparam rnode_226to227_bb4_add_i265_0_reg_227_fifo.DEPTH = 1;
defparam rnode_226to227_bb4_add_i265_0_reg_227_fifo.DATA_WIDTH = 32;
defparam rnode_226to227_bb4_add_i265_0_reg_227_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_226to227_bb4_add_i265_0_reg_227_fifo.IMPL = "shift_reg";

assign rnode_226to227_bb4_add_i265_0_reg_227_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_225to226_bb4_add_i265_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_226to227_bb4_add_i265_0_NO_SHIFT_REG = rnode_226to227_bb4_add_i265_0_reg_227_NO_SHIFT_REG;
assign rnode_226to227_bb4_add_i265_0_stall_in_reg_227_NO_SHIFT_REG = 1'b0;
assign rnode_226to227_bb4_add_i265_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i283_valid_out;
wire local_bb4_reduction_0_i283_stall_in;
wire local_bb4_reduction_0_i283_inputs_ready;
wire local_bb4_reduction_0_i283_stall_local;
wire local_bb4_reduction_0_i283;

assign local_bb4_reduction_0_i283_inputs_ready = (rnode_225to226_bb4_lnot_i228_0_valid_out_1_NO_SHIFT_REG & rnode_225to226_bb4_lnot8_i229_0_valid_out_NO_SHIFT_REG);
assign local_bb4_reduction_0_i283 = (rnode_225to226_bb4_lnot_i228_1_NO_SHIFT_REG | rnode_225to226_bb4_lnot8_i229_0_NO_SHIFT_REG);
assign local_bb4_reduction_0_i283_valid_out = 1'b1;
assign rnode_225to226_bb4_lnot_i228_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot8_i229_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge8_demorgan_i234_stall_local;
wire local_bb4_brmerge8_demorgan_i234;

assign local_bb4_brmerge8_demorgan_i234 = (rnode_225to226_bb4_cmp11_i231_0_NO_SHIFT_REG & rnode_225to226_bb4_lnot17_i233_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u57_valid_out;
wire local_bb4_var__u57_stall_in;
wire local_bb4_var__u57_inputs_ready;
wire local_bb4_var__u57_stall_local;
wire local_bb4_var__u57;

assign local_bb4_var__u57_inputs_ready = (rnode_225to226_bb4_cmp_i230_0_valid_out_3_NO_SHIFT_REG & rnode_225to226_bb4_cmp11_i231_0_valid_out_2_NO_SHIFT_REG);
assign local_bb4_var__u57 = (rnode_225to226_bb4_cmp_i230_3_NO_SHIFT_REG | rnode_225to226_bb4_cmp11_i231_2_NO_SHIFT_REG);
assign local_bb4_var__u57_valid_out = 1'b1;
assign rnode_225to226_bb4_cmp_i230_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp11_i231_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_conv3_i_i259_stall_local;
wire [31:0] local_bb4_conv3_i_i259;
wire [63:0] local_bb4_conv3_i_i259$ps;

assign local_bb4_conv3_i_i259$ps = (local_bb4_mul_i_i258 & 64'hFFFFFFFFFFFF);
assign local_bb4_conv3_i_i259 = local_bb4_conv3_i_i259$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u58_stall_local;
wire [63:0] local_bb4_var__u58;

assign local_bb4_var__u58 = ((local_bb4_mul_i_i258 & 64'hFFFFFFFFFFFF) >> 64'h18);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_xor_i224_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4_xor_i224_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_xor_i224_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_xor_i224_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_xor_i224_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_xor_i224_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_xor_i224_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_xor_i224_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_xor_i224_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_xor_i224_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_xor_i224_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_xor_i224_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_xor_i224_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(rnode_226to229_bb4_xor_i224_0_NO_SHIFT_REG),
	.data_out(rnode_229to230_bb4_xor_i224_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_xor_i224_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_xor_i224_0_reg_230_fifo.DATA_WIDTH = 32;
defparam rnode_229to230_bb4_xor_i224_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_xor_i224_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_xor_i224_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_226to229_bb4_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_xor_i224_0_NO_SHIFT_REG = rnode_229to230_bb4_xor_i224_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_xor_i224_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_xor_i224_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__28_i252_stall_local;
wire local_bb4__28_i252;

assign local_bb4__28_i252 = (rnode_225to226_bb4_cmp_i230_2_NO_SHIFT_REG & local_bb4_lnot14_not_i251);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_227to228_bb4_add_i265_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_227to228_bb4_add_i265_0_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_227to228_bb4_add_i265_1_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_227to228_bb4_add_i265_2_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_reg_228_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_227to228_bb4_add_i265_0_reg_228_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_valid_out_0_reg_228_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_stall_in_0_reg_228_NO_SHIFT_REG;
 logic rnode_227to228_bb4_add_i265_0_stall_out_reg_228_NO_SHIFT_REG;

acl_data_fifo rnode_227to228_bb4_add_i265_0_reg_228_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_227to228_bb4_add_i265_0_reg_228_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_227to228_bb4_add_i265_0_stall_in_0_reg_228_NO_SHIFT_REG),
	.valid_out(rnode_227to228_bb4_add_i265_0_valid_out_0_reg_228_NO_SHIFT_REG),
	.stall_out(rnode_227to228_bb4_add_i265_0_stall_out_reg_228_NO_SHIFT_REG),
	.data_in((rnode_226to227_bb4_add_i265_0_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_227to228_bb4_add_i265_0_reg_228_NO_SHIFT_REG)
);

defparam rnode_227to228_bb4_add_i265_0_reg_228_fifo.DEPTH = 1;
defparam rnode_227to228_bb4_add_i265_0_reg_228_fifo.DATA_WIDTH = 32;
defparam rnode_227to228_bb4_add_i265_0_reg_228_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_227to228_bb4_add_i265_0_reg_228_fifo.IMPL = "shift_reg";

assign rnode_227to228_bb4_add_i265_0_reg_228_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_226to227_bb4_add_i265_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_227to228_bb4_add_i265_0_stall_in_0_reg_228_NO_SHIFT_REG = 1'b0;
assign rnode_227to228_bb4_add_i265_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_227to228_bb4_add_i265_0_NO_SHIFT_REG = rnode_227to228_bb4_add_i265_0_reg_228_NO_SHIFT_REG;
assign rnode_227to228_bb4_add_i265_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_227to228_bb4_add_i265_1_NO_SHIFT_REG = rnode_227to228_bb4_add_i265_0_reg_228_NO_SHIFT_REG;
assign rnode_227to228_bb4_add_i265_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_227to228_bb4_add_i265_2_NO_SHIFT_REG = rnode_227to228_bb4_add_i265_0_reg_228_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_226to227_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_226to227_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_226to227_bb4_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_226to227_bb4_reduction_0_i283_0_reg_227_inputs_ready_NO_SHIFT_REG;
 logic rnode_226to227_bb4_reduction_0_i283_0_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_reduction_0_i283_0_valid_out_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_reduction_0_i283_0_stall_in_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_reduction_0_i283_0_stall_out_reg_227_NO_SHIFT_REG;

acl_data_fifo rnode_226to227_bb4_reduction_0_i283_0_reg_227_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_226to227_bb4_reduction_0_i283_0_reg_227_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_226to227_bb4_reduction_0_i283_0_stall_in_reg_227_NO_SHIFT_REG),
	.valid_out(rnode_226to227_bb4_reduction_0_i283_0_valid_out_reg_227_NO_SHIFT_REG),
	.stall_out(rnode_226to227_bb4_reduction_0_i283_0_stall_out_reg_227_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_0_i283),
	.data_out(rnode_226to227_bb4_reduction_0_i283_0_reg_227_NO_SHIFT_REG)
);

defparam rnode_226to227_bb4_reduction_0_i283_0_reg_227_fifo.DEPTH = 1;
defparam rnode_226to227_bb4_reduction_0_i283_0_reg_227_fifo.DATA_WIDTH = 1;
defparam rnode_226to227_bb4_reduction_0_i283_0_reg_227_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_226to227_bb4_reduction_0_i283_0_reg_227_fifo.IMPL = "shift_reg";

assign rnode_226to227_bb4_reduction_0_i283_0_reg_227_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_0_i283_stall_in = 1'b0;
assign rnode_226to227_bb4_reduction_0_i283_0_NO_SHIFT_REG = rnode_226to227_bb4_reduction_0_i283_0_reg_227_NO_SHIFT_REG;
assign rnode_226to227_bb4_reduction_0_i283_0_stall_in_reg_227_NO_SHIFT_REG = 1'b0;
assign rnode_226to227_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge10_demorgan_i235_stall_local;
wire local_bb4_brmerge10_demorgan_i235;

assign local_bb4_brmerge10_demorgan_i235 = (local_bb4_brmerge8_demorgan_i234 & rnode_225to226_bb4_lnot_i228_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__mux9_mux_i236_stall_local;
wire local_bb4__mux9_mux_i236;

assign local_bb4__mux9_mux_i236 = (local_bb4_brmerge8_demorgan_i234 ^ rnode_225to226_bb4_cmp11_i231_1_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_226to227_bb4_var__u57_0_valid_out_NO_SHIFT_REG;
 logic rnode_226to227_bb4_var__u57_0_stall_in_NO_SHIFT_REG;
 logic rnode_226to227_bb4_var__u57_0_NO_SHIFT_REG;
 logic rnode_226to227_bb4_var__u57_0_reg_227_inputs_ready_NO_SHIFT_REG;
 logic rnode_226to227_bb4_var__u57_0_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_var__u57_0_valid_out_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_var__u57_0_stall_in_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4_var__u57_0_stall_out_reg_227_NO_SHIFT_REG;

acl_data_fifo rnode_226to227_bb4_var__u57_0_reg_227_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_226to227_bb4_var__u57_0_reg_227_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_226to227_bb4_var__u57_0_stall_in_reg_227_NO_SHIFT_REG),
	.valid_out(rnode_226to227_bb4_var__u57_0_valid_out_reg_227_NO_SHIFT_REG),
	.stall_out(rnode_226to227_bb4_var__u57_0_stall_out_reg_227_NO_SHIFT_REG),
	.data_in(local_bb4_var__u57),
	.data_out(rnode_226to227_bb4_var__u57_0_reg_227_NO_SHIFT_REG)
);

defparam rnode_226to227_bb4_var__u57_0_reg_227_fifo.DEPTH = 1;
defparam rnode_226to227_bb4_var__u57_0_reg_227_fifo.DATA_WIDTH = 1;
defparam rnode_226to227_bb4_var__u57_0_reg_227_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_226to227_bb4_var__u57_0_reg_227_fifo.IMPL = "shift_reg";

assign rnode_226to227_bb4_var__u57_0_reg_227_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u57_stall_in = 1'b0;
assign rnode_226to227_bb4_var__u57_0_NO_SHIFT_REG = rnode_226to227_bb4_var__u57_0_reg_227_NO_SHIFT_REG;
assign rnode_226to227_bb4_var__u57_0_stall_in_reg_227_NO_SHIFT_REG = 1'b0;
assign rnode_226to227_bb4_var__u57_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i16_i262_stall_local;
wire [31:0] local_bb4_shr_i16_i262;

assign local_bb4_shr_i16_i262 = (local_bb4_conv3_i_i259 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i18_i264_stall_local;
wire [31:0] local_bb4_shl1_i18_i264;

assign local_bb4_shl1_i18_i264 = (local_bb4_conv3_i_i259 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u59_stall_local;
wire [31:0] local_bb4_var__u59;

assign local_bb4_var__u59 = (local_bb4_conv3_i_i259 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i_i272_stall_local;
wire [31:0] local_bb4_shl1_i_i272;

assign local_bb4_shl1_i_i272 = (local_bb4_conv3_i_i259 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb4__tr_i260_stall_local;
wire [31:0] local_bb4__tr_i260;
wire [63:0] local_bb4__tr_i260$ps;

assign local_bb4__tr_i260$ps = (local_bb4_var__u58 & 64'hFFFFFF);
assign local_bb4__tr_i260 = local_bb4__tr_i260$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_and4_i225_stall_local;
wire [31:0] local_bb4_and4_i225;

assign local_bb4_and4_i225 = (rnode_229to230_bb4_xor_i224_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_inc_i268_stall_local;
wire [31:0] local_bb4_inc_i268;

assign local_bb4_inc_i268 = ((rnode_227to228_bb4_add_i265_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp50_not_i273_stall_local;
wire local_bb4_cmp50_not_i273;

assign local_bb4_cmp50_not_i273 = ((rnode_227to228_bb4_add_i265_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_227to229_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_227to229_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_227to229_bb4_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_227to229_bb4_reduction_0_i283_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic rnode_227to229_bb4_reduction_0_i283_0_reg_229_NO_SHIFT_REG;
 logic rnode_227to229_bb4_reduction_0_i283_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_227to229_bb4_reduction_0_i283_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_227to229_bb4_reduction_0_i283_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_227to229_bb4_reduction_0_i283_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_227to229_bb4_reduction_0_i283_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_227to229_bb4_reduction_0_i283_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_227to229_bb4_reduction_0_i283_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_227to229_bb4_reduction_0_i283_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in(rnode_226to227_bb4_reduction_0_i283_0_NO_SHIFT_REG),
	.data_out(rnode_227to229_bb4_reduction_0_i283_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_227to229_bb4_reduction_0_i283_0_reg_229_fifo.DEPTH = 2;
defparam rnode_227to229_bb4_reduction_0_i283_0_reg_229_fifo.DATA_WIDTH = 1;
defparam rnode_227to229_bb4_reduction_0_i283_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_227to229_bb4_reduction_0_i283_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_227to229_bb4_reduction_0_i283_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_226to227_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_227to229_bb4_reduction_0_i283_0_NO_SHIFT_REG = rnode_227to229_bb4_reduction_0_i283_0_reg_229_NO_SHIFT_REG;
assign rnode_227to229_bb4_reduction_0_i283_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_227to229_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__24_i247_stall_local;
wire local_bb4__24_i247;

assign local_bb4__24_i247 = (rnode_225to226_bb4_cmp_i230_0_NO_SHIFT_REG ? rnode_225to226_bb4_reduction_6_i246_0_NO_SHIFT_REG : local_bb4_brmerge10_demorgan_i235);

// This section implements an unregistered operation.
// 
wire local_bb4__26_demorgan_i249_stall_local;
wire local_bb4__26_demorgan_i249;

assign local_bb4__26_demorgan_i249 = (rnode_225to226_bb4_cmp_i230_1_NO_SHIFT_REG | local_bb4_brmerge10_demorgan_i235);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_227to228_bb4_var__u57_0_valid_out_NO_SHIFT_REG;
 logic rnode_227to228_bb4_var__u57_0_stall_in_NO_SHIFT_REG;
 logic rnode_227to228_bb4_var__u57_0_NO_SHIFT_REG;
 logic rnode_227to228_bb4_var__u57_0_reg_228_inputs_ready_NO_SHIFT_REG;
 logic rnode_227to228_bb4_var__u57_0_reg_228_NO_SHIFT_REG;
 logic rnode_227to228_bb4_var__u57_0_valid_out_reg_228_NO_SHIFT_REG;
 logic rnode_227to228_bb4_var__u57_0_stall_in_reg_228_NO_SHIFT_REG;
 logic rnode_227to228_bb4_var__u57_0_stall_out_reg_228_NO_SHIFT_REG;

acl_data_fifo rnode_227to228_bb4_var__u57_0_reg_228_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_227to228_bb4_var__u57_0_reg_228_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_227to228_bb4_var__u57_0_stall_in_reg_228_NO_SHIFT_REG),
	.valid_out(rnode_227to228_bb4_var__u57_0_valid_out_reg_228_NO_SHIFT_REG),
	.stall_out(rnode_227to228_bb4_var__u57_0_stall_out_reg_228_NO_SHIFT_REG),
	.data_in(rnode_226to227_bb4_var__u57_0_NO_SHIFT_REG),
	.data_out(rnode_227to228_bb4_var__u57_0_reg_228_NO_SHIFT_REG)
);

defparam rnode_227to228_bb4_var__u57_0_reg_228_fifo.DEPTH = 1;
defparam rnode_227to228_bb4_var__u57_0_reg_228_fifo.DATA_WIDTH = 1;
defparam rnode_227to228_bb4_var__u57_0_reg_228_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_227to228_bb4_var__u57_0_reg_228_fifo.IMPL = "shift_reg";

assign rnode_227to228_bb4_var__u57_0_reg_228_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_226to227_bb4_var__u57_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_227to228_bb4_var__u57_0_NO_SHIFT_REG = rnode_227to228_bb4_var__u57_0_reg_228_NO_SHIFT_REG;
assign rnode_227to228_bb4_var__u57_0_stall_in_reg_228_NO_SHIFT_REG = 1'b0;
assign rnode_227to228_bb4_var__u57_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i270_stall_local;
wire [31:0] local_bb4_shr_i_i270;

assign local_bb4_shr_i_i270 = ((local_bb4_var__u59 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i15_i261_stall_local;
wire [31:0] local_bb4_shl_i15_i261;

assign local_bb4_shl_i15_i261 = ((local_bb4__tr_i260 & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb4_and48_i266_stall_local;
wire [31:0] local_bb4_and48_i266;

assign local_bb4_and48_i266 = ((local_bb4__tr_i260 & 32'hFFFFFF) & 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG;
 logic rnode_229to230_bb4_reduction_0_i283_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_reduction_0_i283_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic rnode_229to230_bb4_reduction_0_i283_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_reduction_0_i283_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_reduction_0_i283_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_reduction_0_i283_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_reduction_0_i283_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_reduction_0_i283_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_reduction_0_i283_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_reduction_0_i283_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_reduction_0_i283_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(rnode_227to229_bb4_reduction_0_i283_0_NO_SHIFT_REG),
	.data_out(rnode_229to230_bb4_reduction_0_i283_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_reduction_0_i283_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_reduction_0_i283_0_reg_230_fifo.DATA_WIDTH = 1;
defparam rnode_229to230_bb4_reduction_0_i283_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_reduction_0_i283_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_reduction_0_i283_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_227to229_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_reduction_0_i283_0_NO_SHIFT_REG = rnode_229to230_bb4_reduction_0_i283_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_reduction_0_i283_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__25_i248_stall_local;
wire local_bb4__25_i248;

assign local_bb4__25_i248 = (local_bb4__24_i247 ? rnode_225to226_bb4_lnot14_i232_0_NO_SHIFT_REG : rnode_225to226_bb4__mux_mux_mux_i242_0_NO_SHIFT_REG);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_228to229_bb4_var__u57_0_valid_out_NO_SHIFT_REG;
 logic rnode_228to229_bb4_var__u57_0_stall_in_NO_SHIFT_REG;
 logic rnode_228to229_bb4_var__u57_0_NO_SHIFT_REG;
 logic rnode_228to229_bb4_var__u57_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic rnode_228to229_bb4_var__u57_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_var__u57_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_var__u57_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_var__u57_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_228to229_bb4_var__u57_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_228to229_bb4_var__u57_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_228to229_bb4_var__u57_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_228to229_bb4_var__u57_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_228to229_bb4_var__u57_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in(rnode_227to228_bb4_var__u57_0_NO_SHIFT_REG),
	.data_out(rnode_228to229_bb4_var__u57_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_228to229_bb4_var__u57_0_reg_229_fifo.DEPTH = 1;
defparam rnode_228to229_bb4_var__u57_0_reg_229_fifo.DATA_WIDTH = 1;
defparam rnode_228to229_bb4_var__u57_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_228to229_bb4_var__u57_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_228to229_bb4_var__u57_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_227to228_bb4_var__u57_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4_var__u57_0_NO_SHIFT_REG = rnode_228to229_bb4_var__u57_0_reg_229_NO_SHIFT_REG;
assign rnode_228to229_bb4_var__u57_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4_var__u57_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_i17_i263_stall_local;
wire [31:0] local_bb4_or_i17_i263;

assign local_bb4_or_i17_i263 = ((local_bb4_shl_i15_i261 & 32'hFFFF00) | (local_bb4_shr_i16_i262 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool49_i267_stall_local;
wire local_bb4_tobool49_i267;

assign local_bb4_tobool49_i267 = ((local_bb4_and48_i266 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i250_stall_local;
wire local_bb4__27_i250;

assign local_bb4__27_i250 = (local_bb4__26_demorgan_i249 ? local_bb4__25_i248 : local_bb4__mux9_mux_i236);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_i269_stall_local;
wire [31:0] local_bb4_shl_i_i269;

assign local_bb4_shl_i_i269 = ((local_bb4_or_i17_i263 & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__31_i274_stall_local;
wire local_bb4__31_i274;

assign local_bb4__31_i274 = (local_bb4_tobool49_i267 & local_bb4_cmp50_not_i273);

// This section implements an unregistered operation.
// 
wire local_bb4__29_i253_valid_out;
wire local_bb4__29_i253_stall_in;
wire local_bb4__29_i253_inputs_ready;
wire local_bb4__29_i253_stall_local;
wire local_bb4__29_i253;

assign local_bb4__29_i253_inputs_ready = (rnode_225to226_bb4_lnot14_i232_0_valid_out_0_NO_SHIFT_REG & rnode_225to226_bb4__mux_mux_mux_i242_0_valid_out_NO_SHIFT_REG & rnode_225to226_bb4_lnot_i228_0_valid_out_0_NO_SHIFT_REG & rnode_225to226_bb4_cmp_i230_0_valid_out_0_NO_SHIFT_REG & rnode_225to226_bb4_reduction_6_i246_0_valid_out_NO_SHIFT_REG & rnode_225to226_bb4_cmp_i230_0_valid_out_1_NO_SHIFT_REG & rnode_225to226_bb4_lnot14_i232_0_valid_out_1_NO_SHIFT_REG & rnode_225to226_bb4_cmp_i230_0_valid_out_2_NO_SHIFT_REG & rnode_225to226_bb4_cmp11_i231_0_valid_out_0_NO_SHIFT_REG & rnode_225to226_bb4_lnot17_i233_0_valid_out_NO_SHIFT_REG & rnode_225to226_bb4_cmp11_i231_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4__29_i253 = (local_bb4__28_i252 | local_bb4__27_i250);
assign local_bb4__29_i253_valid_out = 1'b1;
assign rnode_225to226_bb4_lnot14_i232_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4__mux_mux_mux_i242_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot_i228_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp_i230_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_reduction_6_i246_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp_i230_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot14_i232_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp_i230_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp11_i231_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_lnot17_i233_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_225to226_bb4_cmp11_i231_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i271_stall_local;
wire [31:0] local_bb4_or_i_i271;

assign local_bb4_or_i_i271 = ((local_bb4_shl_i_i269 & 32'h1FFFFFE) | (local_bb4_shr_i_i270 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i275_stall_local;
wire [31:0] local_bb4__32_i275;

assign local_bb4__32_i275 = (local_bb4__31_i274 ? (local_bb4_shl1_i_i272 & 32'hFFFFFE00) : (local_bb4_shl1_i18_i264 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__36_i279_stall_local;
wire [31:0] local_bb4__36_i279;

assign local_bb4__36_i279 = (local_bb4__31_i274 ? (rnode_227to228_bb4_add_i265_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_226to227_bb4__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_226to227_bb4__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_226to227_bb4__29_i253_0_NO_SHIFT_REG;
 logic rnode_226to227_bb4__29_i253_0_reg_227_inputs_ready_NO_SHIFT_REG;
 logic rnode_226to227_bb4__29_i253_0_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4__29_i253_0_valid_out_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4__29_i253_0_stall_in_reg_227_NO_SHIFT_REG;
 logic rnode_226to227_bb4__29_i253_0_stall_out_reg_227_NO_SHIFT_REG;

acl_data_fifo rnode_226to227_bb4__29_i253_0_reg_227_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_226to227_bb4__29_i253_0_reg_227_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_226to227_bb4__29_i253_0_stall_in_reg_227_NO_SHIFT_REG),
	.valid_out(rnode_226to227_bb4__29_i253_0_valid_out_reg_227_NO_SHIFT_REG),
	.stall_out(rnode_226to227_bb4__29_i253_0_stall_out_reg_227_NO_SHIFT_REG),
	.data_in(local_bb4__29_i253),
	.data_out(rnode_226to227_bb4__29_i253_0_reg_227_NO_SHIFT_REG)
);

defparam rnode_226to227_bb4__29_i253_0_reg_227_fifo.DEPTH = 1;
defparam rnode_226to227_bb4__29_i253_0_reg_227_fifo.DATA_WIDTH = 1;
defparam rnode_226to227_bb4__29_i253_0_reg_227_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_226to227_bb4__29_i253_0_reg_227_fifo.IMPL = "shift_reg";

assign rnode_226to227_bb4__29_i253_0_reg_227_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__29_i253_stall_in = 1'b0;
assign rnode_226to227_bb4__29_i253_0_NO_SHIFT_REG = rnode_226to227_bb4__29_i253_0_reg_227_NO_SHIFT_REG;
assign rnode_226to227_bb4__29_i253_0_stall_in_reg_227_NO_SHIFT_REG = 1'b0;
assign rnode_226to227_bb4__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__34_i277_stall_local;
wire [31:0] local_bb4__34_i277;

assign local_bb4__34_i277 = (local_bb4__31_i274 ? (local_bb4_or_i_i271 & 32'h1FFFFFF) : (local_bb4_or_i17_i263 & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i276_stall_local;
wire [31:0] local_bb4__33_i276;

assign local_bb4__33_i276 = (local_bb4_tobool49_i267 ? (local_bb4__32_i275 & 32'hFFFFFF00) : (local_bb4_shl1_i18_i264 & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__37_i280_stall_local;
wire [31:0] local_bb4__37_i280;

assign local_bb4__37_i280 = (local_bb4_tobool49_i267 ? (local_bb4__36_i279 & 32'h1FF) : (local_bb4_inc_i268 & 32'h3FF));

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_227to229_bb4__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_227to229_bb4__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_227to229_bb4__29_i253_0_NO_SHIFT_REG;
 logic rnode_227to229_bb4__29_i253_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic rnode_227to229_bb4__29_i253_0_reg_229_NO_SHIFT_REG;
 logic rnode_227to229_bb4__29_i253_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_227to229_bb4__29_i253_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_227to229_bb4__29_i253_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_227to229_bb4__29_i253_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_227to229_bb4__29_i253_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_227to229_bb4__29_i253_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_227to229_bb4__29_i253_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_227to229_bb4__29_i253_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in(rnode_226to227_bb4__29_i253_0_NO_SHIFT_REG),
	.data_out(rnode_227to229_bb4__29_i253_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_227to229_bb4__29_i253_0_reg_229_fifo.DEPTH = 2;
defparam rnode_227to229_bb4__29_i253_0_reg_229_fifo.DATA_WIDTH = 1;
defparam rnode_227to229_bb4__29_i253_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_227to229_bb4__29_i253_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_227to229_bb4__29_i253_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_226to227_bb4__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_227to229_bb4__29_i253_0_NO_SHIFT_REG = rnode_227to229_bb4__29_i253_0_reg_229_NO_SHIFT_REG;
assign rnode_227to229_bb4__29_i253_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_227to229_bb4__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__35_i278_stall_local;
wire [31:0] local_bb4__35_i278;

assign local_bb4__35_i278 = (local_bb4_tobool49_i267 ? (local_bb4__34_i277 & 32'h1FFFFFF) : (local_bb4_or_i17_i263 & 32'hFFFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4__29_i253_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4__29_i253_0_stall_in_NO_SHIFT_REG;
 logic rnode_229to230_bb4__29_i253_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4__29_i253_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic rnode_229to230_bb4__29_i253_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4__29_i253_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4__29_i253_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4__29_i253_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4__29_i253_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4__29_i253_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4__29_i253_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4__29_i253_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4__29_i253_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(rnode_227to229_bb4__29_i253_0_NO_SHIFT_REG),
	.data_out(rnode_229to230_bb4__29_i253_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4__29_i253_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4__29_i253_0_reg_230_fifo.DATA_WIDTH = 1;
defparam rnode_229to230_bb4__29_i253_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4__29_i253_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4__29_i253_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_227to229_bb4__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4__29_i253_0_NO_SHIFT_REG = rnode_229to230_bb4__29_i253_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4__29_i253_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4__29_i253_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i286_stall_local;
wire [31:0] local_bb4_and75_i286;

assign local_bb4_and75_i286 = ((local_bb4__35_i278 & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i276_valid_out;
wire local_bb4__33_i276_stall_in;
wire local_bb4__37_i280_valid_out;
wire local_bb4__37_i280_stall_in;
wire local_bb4_and75_i286_valid_out;
wire local_bb4_and75_i286_stall_in;
wire local_bb4_and83_i292_valid_out;
wire local_bb4_and83_i292_stall_in;
wire local_bb4_and83_i292_inputs_ready;
wire local_bb4_and83_i292_stall_local;
wire [31:0] local_bb4_and83_i292;

assign local_bb4_and83_i292_inputs_ready = (local_bb4_mul_i_i258_valid_out_0_NO_SHIFT_REG & local_bb4_mul_i_i258_valid_out_1_NO_SHIFT_REG & rnode_227to228_bb4_add_i265_0_valid_out_1_NO_SHIFT_REG & rnode_227to228_bb4_add_i265_0_valid_out_0_NO_SHIFT_REG & rnode_227to228_bb4_add_i265_0_valid_out_2_NO_SHIFT_REG);
assign local_bb4_and83_i292 = ((local_bb4__35_i278 & 32'h1FFFFFF) & 32'h1);
assign local_bb4__33_i276_valid_out = 1'b1;
assign local_bb4__37_i280_valid_out = 1'b1;
assign local_bb4_and75_i286_valid_out = 1'b1;
assign local_bb4_and83_i292_valid_out = 1'b1;
assign local_bb4_mul_i_i258_stall_in_0 = 1'b0;
assign local_bb4_mul_i_i258_stall_in_1 = 1'b0;
assign rnode_227to228_bb4_add_i265_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_227to228_bb4_add_i265_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_227to228_bb4_add_i265_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_228to229_bb4__33_i276_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_228to229_bb4__33_i276_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__33_i276_0_NO_SHIFT_REG;
 logic rnode_228to229_bb4__33_i276_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_228to229_bb4__33_i276_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__33_i276_1_NO_SHIFT_REG;
 logic rnode_228to229_bb4__33_i276_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__33_i276_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4__33_i276_0_valid_out_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4__33_i276_0_stall_in_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4__33_i276_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_228to229_bb4__33_i276_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_228to229_bb4__33_i276_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_228to229_bb4__33_i276_0_stall_in_0_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_228to229_bb4__33_i276_0_valid_out_0_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_228to229_bb4__33_i276_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in((local_bb4__33_i276 & 32'hFFFFFF00)),
	.data_out(rnode_228to229_bb4__33_i276_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_228to229_bb4__33_i276_0_reg_229_fifo.DEPTH = 1;
defparam rnode_228to229_bb4__33_i276_0_reg_229_fifo.DATA_WIDTH = 32;
defparam rnode_228to229_bb4__33_i276_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_228to229_bb4__33_i276_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_228to229_bb4__33_i276_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__33_i276_stall_in = 1'b0;
assign rnode_228to229_bb4__33_i276_0_stall_in_0_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4__33_i276_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_228to229_bb4__33_i276_0_NO_SHIFT_REG = rnode_228to229_bb4__33_i276_0_reg_229_NO_SHIFT_REG;
assign rnode_228to229_bb4__33_i276_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_228to229_bb4__33_i276_1_NO_SHIFT_REG = rnode_228to229_bb4__33_i276_0_reg_229_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_228to229_bb4__37_i280_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__37_i280_0_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__37_i280_1_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__37_i280_2_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__37_i280_3_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4__37_i280_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_valid_out_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_stall_in_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4__37_i280_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_228to229_bb4__37_i280_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_228to229_bb4__37_i280_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_228to229_bb4__37_i280_0_stall_in_0_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_228to229_bb4__37_i280_0_valid_out_0_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_228to229_bb4__37_i280_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in((local_bb4__37_i280 & 32'h3FF)),
	.data_out(rnode_228to229_bb4__37_i280_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_228to229_bb4__37_i280_0_reg_229_fifo.DEPTH = 1;
defparam rnode_228to229_bb4__37_i280_0_reg_229_fifo.DATA_WIDTH = 32;
defparam rnode_228to229_bb4__37_i280_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_228to229_bb4__37_i280_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_228to229_bb4__37_i280_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__37_i280_stall_in = 1'b0;
assign rnode_228to229_bb4__37_i280_0_stall_in_0_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4__37_i280_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_228to229_bb4__37_i280_0_NO_SHIFT_REG = rnode_228to229_bb4__37_i280_0_reg_229_NO_SHIFT_REG;
assign rnode_228to229_bb4__37_i280_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_228to229_bb4__37_i280_1_NO_SHIFT_REG = rnode_228to229_bb4__37_i280_0_reg_229_NO_SHIFT_REG;
assign rnode_228to229_bb4__37_i280_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_228to229_bb4__37_i280_2_NO_SHIFT_REG = rnode_228to229_bb4__37_i280_0_reg_229_NO_SHIFT_REG;
assign rnode_228to229_bb4__37_i280_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_228to229_bb4__37_i280_3_NO_SHIFT_REG = rnode_228to229_bb4__37_i280_0_reg_229_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_228to229_bb4_and75_i286_0_valid_out_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and75_i286_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4_and75_i286_0_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and75_i286_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4_and75_i286_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and75_i286_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and75_i286_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and75_i286_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_228to229_bb4_and75_i286_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_228to229_bb4_and75_i286_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_228to229_bb4_and75_i286_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_228to229_bb4_and75_i286_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_228to229_bb4_and75_i286_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in((local_bb4_and75_i286 & 32'h7FFFFF)),
	.data_out(rnode_228to229_bb4_and75_i286_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_228to229_bb4_and75_i286_0_reg_229_fifo.DEPTH = 1;
defparam rnode_228to229_bb4_and75_i286_0_reg_229_fifo.DATA_WIDTH = 32;
defparam rnode_228to229_bb4_and75_i286_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_228to229_bb4_and75_i286_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_228to229_bb4_and75_i286_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and75_i286_stall_in = 1'b0;
assign rnode_228to229_bb4_and75_i286_0_NO_SHIFT_REG = rnode_228to229_bb4_and75_i286_0_reg_229_NO_SHIFT_REG;
assign rnode_228to229_bb4_and75_i286_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4_and75_i286_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_228to229_bb4_and83_i292_0_valid_out_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and83_i292_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4_and83_i292_0_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and83_i292_0_reg_229_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_228to229_bb4_and83_i292_0_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and83_i292_0_valid_out_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and83_i292_0_stall_in_reg_229_NO_SHIFT_REG;
 logic rnode_228to229_bb4_and83_i292_0_stall_out_reg_229_NO_SHIFT_REG;

acl_data_fifo rnode_228to229_bb4_and83_i292_0_reg_229_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_228to229_bb4_and83_i292_0_reg_229_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_228to229_bb4_and83_i292_0_stall_in_reg_229_NO_SHIFT_REG),
	.valid_out(rnode_228to229_bb4_and83_i292_0_valid_out_reg_229_NO_SHIFT_REG),
	.stall_out(rnode_228to229_bb4_and83_i292_0_stall_out_reg_229_NO_SHIFT_REG),
	.data_in((local_bb4_and83_i292 & 32'h1)),
	.data_out(rnode_228to229_bb4_and83_i292_0_reg_229_NO_SHIFT_REG)
);

defparam rnode_228to229_bb4_and83_i292_0_reg_229_fifo.DEPTH = 1;
defparam rnode_228to229_bb4_and83_i292_0_reg_229_fifo.DATA_WIDTH = 32;
defparam rnode_228to229_bb4_and83_i292_0_reg_229_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_228to229_bb4_and83_i292_0_reg_229_fifo.IMPL = "shift_reg";

assign rnode_228to229_bb4_and83_i292_0_reg_229_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and83_i292_stall_in = 1'b0;
assign rnode_228to229_bb4_and83_i292_0_NO_SHIFT_REG = rnode_228to229_bb4_and83_i292_0_reg_229_NO_SHIFT_REG;
assign rnode_228to229_bb4_and83_i292_0_stall_in_reg_229_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4_and83_i292_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i291_stall_local;
wire local_bb4_cmp77_i291;

assign local_bb4_cmp77_i291 = ((rnode_228to229_bb4__33_i276_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u60_stall_local;
wire local_bb4_var__u60;

assign local_bb4_var__u60 = ($signed((rnode_228to229_bb4__33_i276_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp53_i281_stall_local;
wire local_bb4_cmp53_i281;

assign local_bb4_cmp53_i281 = ((rnode_228to229_bb4__37_i280_0_NO_SHIFT_REG & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp68_i285_valid_out;
wire local_bb4_cmp68_i285_stall_in;
wire local_bb4_cmp68_i285_inputs_ready;
wire local_bb4_cmp68_i285_stall_local;
wire local_bb4_cmp68_i285;

assign local_bb4_cmp68_i285_inputs_ready = rnode_228to229_bb4__37_i280_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp68_i285 = ((rnode_228to229_bb4__37_i280_1_NO_SHIFT_REG & 32'h3FF) < 32'h80);
assign local_bb4_cmp68_i285_valid_out = 1'b1;
assign rnode_228to229_bb4__37_i280_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i287_stall_local;
wire [31:0] local_bb4_sub_i287;

assign local_bb4_sub_i287 = ((rnode_228to229_bb4__37_i280_2_NO_SHIFT_REG & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp71_not_i302_valid_out;
wire local_bb4_cmp71_not_i302_stall_in;
wire local_bb4_cmp71_not_i302_inputs_ready;
wire local_bb4_cmp71_not_i302_stall_local;
wire local_bb4_cmp71_not_i302;

assign local_bb4_cmp71_not_i302_inputs_ready = rnode_228to229_bb4__37_i280_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4_cmp71_not_i302 = ((rnode_228to229_bb4__37_i280_3_NO_SHIFT_REG & 32'h3FF) != 32'h7F);
assign local_bb4_cmp71_not_i302_valid_out = 1'b1;
assign rnode_228to229_bb4__37_i280_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool84_i293_stall_local;
wire local_bb4_tobool84_i293;

assign local_bb4_tobool84_i293 = ((rnode_228to229_bb4_and83_i292_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or581_i282_valid_out;
wire local_bb4_or581_i282_stall_in;
wire local_bb4_or581_i282_inputs_ready;
wire local_bb4_or581_i282_stall_local;
wire local_bb4_or581_i282;

assign local_bb4_or581_i282_inputs_ready = (rnode_228to229_bb4_var__u57_0_valid_out_NO_SHIFT_REG & rnode_228to229_bb4__37_i280_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_or581_i282 = (rnode_228to229_bb4_var__u57_0_NO_SHIFT_REG | local_bb4_cmp53_i281);
assign local_bb4_or581_i282_valid_out = 1'b1;
assign rnode_228to229_bb4_var__u57_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4__37_i280_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_cmp68_i285_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp68_i285_0_stall_in_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp68_i285_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp68_i285_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp68_i285_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp68_i285_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp68_i285_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp68_i285_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_cmp68_i285_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_cmp68_i285_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_cmp68_i285_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_cmp68_i285_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_cmp68_i285_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(local_bb4_cmp68_i285),
	.data_out(rnode_229to230_bb4_cmp68_i285_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_cmp68_i285_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_cmp68_i285_0_reg_230_fifo.DATA_WIDTH = 1;
defparam rnode_229to230_bb4_cmp68_i285_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_cmp68_i285_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_cmp68_i285_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp68_i285_stall_in = 1'b0;
assign rnode_229to230_bb4_cmp68_i285_0_NO_SHIFT_REG = rnode_229to230_bb4_cmp68_i285_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_cmp68_i285_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_cmp68_i285_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and74_i288_stall_local;
wire [31:0] local_bb4_and74_i288;

assign local_bb4_and74_i288 = ((local_bb4_sub_i287 & 32'hFF800000) + 32'h40800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_cmp71_not_i302_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp71_not_i302_0_stall_in_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp71_not_i302_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp71_not_i302_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp71_not_i302_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp71_not_i302_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp71_not_i302_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_cmp71_not_i302_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_cmp71_not_i302_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_cmp71_not_i302_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_cmp71_not_i302_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_cmp71_not_i302_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_cmp71_not_i302_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(local_bb4_cmp71_not_i302),
	.data_out(rnode_229to230_bb4_cmp71_not_i302_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_cmp71_not_i302_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_cmp71_not_i302_0_reg_230_fifo.DATA_WIDTH = 1;
defparam rnode_229to230_bb4_cmp71_not_i302_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_cmp71_not_i302_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_cmp71_not_i302_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp71_not_i302_stall_in = 1'b0;
assign rnode_229to230_bb4_cmp71_not_i302_0_NO_SHIFT_REG = rnode_229to230_bb4_cmp71_not_i302_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_cmp71_not_i302_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_cmp71_not_i302_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__39_i294_stall_local;
wire local_bb4__39_i294;

assign local_bb4__39_i294 = (local_bb4_tobool84_i293 & local_bb4_var__u60);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_or581_i282_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_1_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_valid_out_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_stall_in_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or581_i282_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_or581_i282_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_or581_i282_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_or581_i282_0_stall_in_0_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_or581_i282_0_valid_out_0_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_or581_i282_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(local_bb4_or581_i282),
	.data_out(rnode_229to230_bb4_or581_i282_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_or581_i282_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_or581_i282_0_reg_230_fifo.DATA_WIDTH = 1;
defparam rnode_229to230_bb4_or581_i282_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_or581_i282_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_or581_i282_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or581_i282_stall_in = 1'b0;
assign rnode_229to230_bb4_or581_i282_0_stall_in_0_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_or581_i282_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_229to230_bb4_or581_i282_0_NO_SHIFT_REG = rnode_229to230_bb4_or581_i282_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_or581_i282_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_229to230_bb4_or581_i282_1_NO_SHIFT_REG = rnode_229to230_bb4_or581_i282_0_reg_230_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u61_stall_local;
wire [31:0] local_bb4_var__u61;

assign local_bb4_var__u61[31:1] = 31'h0;
assign local_bb4_var__u61[0] = rnode_229to230_bb4_cmp68_i285_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i289_stall_local;
wire [31:0] local_bb4_shl_i289;

assign local_bb4_shl_i289 = ((local_bb4_and74_i288 & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4__40_i295_valid_out;
wire local_bb4__40_i295_stall_in;
wire local_bb4__40_i295_inputs_ready;
wire local_bb4__40_i295_stall_local;
wire local_bb4__40_i295;

assign local_bb4__40_i295_inputs_ready = (rnode_228to229_bb4__33_i276_0_valid_out_0_NO_SHIFT_REG & rnode_228to229_bb4__33_i276_0_valid_out_1_NO_SHIFT_REG & rnode_228to229_bb4_and83_i292_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40_i295 = (local_bb4_cmp77_i291 | local_bb4__39_i294);
assign local_bb4__40_i295_valid_out = 1'b1;
assign rnode_228to229_bb4__33_i276_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4__33_i276_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4_and83_i292_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i284_stall_local;
wire local_bb4_reduction_2_i284;

assign local_bb4_reduction_2_i284 = (rnode_229to230_bb4_reduction_0_i283_0_NO_SHIFT_REG | rnode_229to230_bb4_or581_i282_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cond111_i310_stall_local;
wire [31:0] local_bb4_cond111_i310;

assign local_bb4_cond111_i310 = (rnode_229to230_bb4_or581_i282_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or76_i290_valid_out;
wire local_bb4_or76_i290_stall_in;
wire local_bb4_or76_i290_inputs_ready;
wire local_bb4_or76_i290_stall_local;
wire [31:0] local_bb4_or76_i290;

assign local_bb4_or76_i290_inputs_ready = (rnode_228to229_bb4__37_i280_0_valid_out_2_NO_SHIFT_REG & rnode_228to229_bb4_and75_i286_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or76_i290 = ((local_bb4_shl_i289 & 32'h7F800000) | (rnode_228to229_bb4_and75_i286_0_NO_SHIFT_REG & 32'h7FFFFF));
assign local_bb4_or76_i290_valid_out = 1'b1;
assign rnode_228to229_bb4__37_i280_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_228to229_bb4_and75_i286_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4__40_i295_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4__40_i295_0_stall_in_NO_SHIFT_REG;
 logic rnode_229to230_bb4__40_i295_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4__40_i295_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic rnode_229to230_bb4__40_i295_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4__40_i295_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4__40_i295_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4__40_i295_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4__40_i295_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4__40_i295_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4__40_i295_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4__40_i295_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4__40_i295_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in(local_bb4__40_i295),
	.data_out(rnode_229to230_bb4__40_i295_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4__40_i295_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4__40_i295_0_reg_230_fifo.DATA_WIDTH = 1;
defparam rnode_229to230_bb4__40_i295_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4__40_i295_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4__40_i295_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_i295_stall_in = 1'b0;
assign rnode_229to230_bb4__40_i295_0_NO_SHIFT_REG = rnode_229to230_bb4__40_i295_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4__40_i295_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4__40_i295_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_conv101_i305_stall_local;
wire [31:0] local_bb4_conv101_i305;

assign local_bb4_conv101_i305[31:1] = 31'h0;
assign local_bb4_conv101_i305[0] = local_bb4_reduction_2_i284;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_229to230_bb4_or76_i290_0_valid_out_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or76_i290_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_or76_i290_0_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or76_i290_0_reg_230_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_229to230_bb4_or76_i290_0_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or76_i290_0_valid_out_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or76_i290_0_stall_in_reg_230_NO_SHIFT_REG;
 logic rnode_229to230_bb4_or76_i290_0_stall_out_reg_230_NO_SHIFT_REG;

acl_data_fifo rnode_229to230_bb4_or76_i290_0_reg_230_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_229to230_bb4_or76_i290_0_reg_230_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_229to230_bb4_or76_i290_0_stall_in_reg_230_NO_SHIFT_REG),
	.valid_out(rnode_229to230_bb4_or76_i290_0_valid_out_reg_230_NO_SHIFT_REG),
	.stall_out(rnode_229to230_bb4_or76_i290_0_stall_out_reg_230_NO_SHIFT_REG),
	.data_in((local_bb4_or76_i290 & 32'h7FFFFFFF)),
	.data_out(rnode_229to230_bb4_or76_i290_0_reg_230_NO_SHIFT_REG)
);

defparam rnode_229to230_bb4_or76_i290_0_reg_230_fifo.DEPTH = 1;
defparam rnode_229to230_bb4_or76_i290_0_reg_230_fifo.DATA_WIDTH = 32;
defparam rnode_229to230_bb4_or76_i290_0_reg_230_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_229to230_bb4_or76_i290_0_reg_230_fifo.IMPL = "shift_reg";

assign rnode_229to230_bb4_or76_i290_0_reg_230_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or76_i290_stall_in = 1'b0;
assign rnode_229to230_bb4_or76_i290_0_NO_SHIFT_REG = rnode_229to230_bb4_or76_i290_0_reg_230_NO_SHIFT_REG;
assign rnode_229to230_bb4_or76_i290_0_stall_in_reg_230_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_or76_i290_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cond_i296_stall_local;
wire [31:0] local_bb4_cond_i296;

assign local_bb4_cond_i296[31:1] = 31'h0;
assign local_bb4_cond_i296[0] = rnode_229to230_bb4__40_i295_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add87_i297_stall_local;
wire [31:0] local_bb4_add87_i297;

assign local_bb4_add87_i297 = ((local_bb4_cond_i296 & 32'h1) + (rnode_229to230_bb4_or76_i290_0_NO_SHIFT_REG & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i298_stall_local;
wire [31:0] local_bb4_and88_i298;

assign local_bb4_and88_i298 = (local_bb4_add87_i297 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i300_stall_local;
wire [31:0] local_bb4_and90_i300;

assign local_bb4_and90_i300 = (local_bb4_add87_i297 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_or89_i299_stall_local;
wire [31:0] local_bb4_or89_i299;

assign local_bb4_or89_i299 = ((local_bb4_and88_i298 & 32'h7FFFFFFF) | (local_bb4_and4_i225 & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i301_stall_local;
wire local_bb4_cmp91_i301;

assign local_bb4_cmp91_i301 = ((local_bb4_and90_i300 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge14_i303_stall_local;
wire local_bb4_brmerge14_i303;

assign local_bb4_brmerge14_i303 = (local_bb4_cmp91_i301 | rnode_229to230_bb4_cmp71_not_i302_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_conv99_i304_stall_local;
wire [31:0] local_bb4_conv99_i304;

assign local_bb4_conv99_i304 = (local_bb4_brmerge14_i303 ? (local_bb4_var__u61 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or102_i306_stall_local;
wire [31:0] local_bb4_or102_i306;

assign local_bb4_or102_i306 = ((local_bb4_conv99_i304 & 32'h1) | (local_bb4_conv101_i305 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool103_i307_stall_local;
wire local_bb4_tobool103_i307;

assign local_bb4_tobool103_i307 = ((local_bb4_or102_i306 & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cond107_i308_stall_local;
wire [31:0] local_bb4_cond107_i308;

assign local_bb4_cond107_i308 = (local_bb4_tobool103_i307 ? (local_bb4_and4_i225 & 32'h80000000) : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and108_i309_stall_local;
wire [31:0] local_bb4_and108_i309;

assign local_bb4_and108_i309 = (local_bb4_cond107_i308 & local_bb4_or89_i299);

// This section implements an unregistered operation.
// 
wire local_bb4_or112_i311_stall_local;
wire [31:0] local_bb4_or112_i311;

assign local_bb4_or112_i311 = (local_bb4_and108_i309 | (local_bb4_cond111_i310 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u62_stall_local;
wire [31:0] local_bb4_var__u62;

assign local_bb4_var__u62 = local_bb4_or112_i311;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u63_stall_local;
wire [31:0] local_bb4_var__u63;

assign local_bb4_var__u63 = (rnode_229to230_bb4__29_i253_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb4_var__u62);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u64_stall_local;
wire [31:0] local_bb4_var__u64;

assign local_bb4_var__u64 = local_bb4_var__u63;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u65_stall_local;
wire [31:0] local_bb4_var__u65;

assign local_bb4_var__u65 = local_bb4_var__u63;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i193_stall_local;
wire [31:0] local_bb4_shr_i193;

assign local_bb4_shr_i193 = (local_bb4_var__u64 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i195_stall_local;
wire [31:0] local_bb4_xor_i195;

assign local_bb4_xor_i195 = (local_bb4_var__u37 ^ local_bb4_var__u64);

// This section implements an unregistered operation.
// 
wire local_bb4_and5_i_stall_local;
wire [31:0] local_bb4_and5_i;

assign local_bb4_and5_i = (local_bb4_var__u64 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i205_stall_local;
wire [31:0] local_bb4_or_i205;

assign local_bb4_or_i205 = ((local_bb4_and5_i & 32'h7FFFFF) | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_shr2_i_valid_out;
wire local_bb4_shr2_i_stall_in;
wire local_bb4_xor_i195_valid_out;
wire local_bb4_xor_i195_stall_in;
wire local_bb4_and6_i_valid_out_1;
wire local_bb4_and6_i_stall_in_1;
wire local_bb4_conv1_i_i_valid_out;
wire local_bb4_conv1_i_i_stall_in;
wire local_bb4_var__u65_valid_out;
wire local_bb4_var__u65_stall_in;
wire local_bb4_shr_i193_valid_out;
wire local_bb4_shr_i193_stall_in;
wire local_bb4_and5_i_valid_out_1;
wire local_bb4_and5_i_stall_in_1;
wire local_bb4_conv_i_i_valid_out;
wire local_bb4_conv_i_i_stall_in;
wire local_bb4_conv_i_i_inputs_ready;
wire local_bb4_conv_i_i_stall_local;
wire [63:0] local_bb4_conv_i_i;

assign local_bb4_conv_i_i_inputs_ready = (rnode_229to230_bb4_c1_ene1_0_valid_out_1_NO_SHIFT_REG & rnode_229to230_bb4_xor_i224_0_valid_out_NO_SHIFT_REG & rnode_229to230_bb4__29_i253_0_valid_out_NO_SHIFT_REG & rnode_229to230_bb4_or581_i282_0_valid_out_1_NO_SHIFT_REG & rnode_229to230_bb4_or581_i282_0_valid_out_0_NO_SHIFT_REG & rnode_229to230_bb4_reduction_0_i283_0_valid_out_NO_SHIFT_REG & rnode_229to230_bb4_cmp68_i285_0_valid_out_NO_SHIFT_REG & rnode_229to230_bb4_cmp71_not_i302_0_valid_out_NO_SHIFT_REG & rnode_229to230_bb4__40_i295_0_valid_out_NO_SHIFT_REG & rnode_229to230_bb4_or76_i290_0_valid_out_NO_SHIFT_REG);
assign local_bb4_conv_i_i[63:32] = 32'h0;
assign local_bb4_conv_i_i[31:0] = ((local_bb4_or_i205 & 32'hFFFFFF) | 32'h800000);
assign local_bb4_shr2_i_valid_out = 1'b1;
assign local_bb4_xor_i195_valid_out = 1'b1;
assign local_bb4_and6_i_valid_out_1 = 1'b1;
assign local_bb4_conv1_i_i_valid_out = 1'b1;
assign local_bb4_var__u65_valid_out = 1'b1;
assign local_bb4_shr_i193_valid_out = 1'b1;
assign local_bb4_and5_i_valid_out_1 = 1'b1;
assign local_bb4_conv_i_i_valid_out = 1'b1;
assign rnode_229to230_bb4_c1_ene1_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_xor_i224_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4__29_i253_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_or581_i282_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_or581_i282_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_reduction_0_i283_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_cmp68_i285_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_cmp71_not_i302_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4__40_i295_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_229to230_bb4_or76_i290_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_shr2_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr2_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_shr2_i_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr2_i_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_shr2_i_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr2_i_0_valid_out_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr2_i_0_stall_in_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr2_i_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_shr2_i_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_shr2_i_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_shr2_i_0_stall_in_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_shr2_i_0_valid_out_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_shr2_i_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in((local_bb4_shr2_i & 32'h1FF)),
	.data_out(rnode_230to231_bb4_shr2_i_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_shr2_i_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_shr2_i_0_reg_231_fifo.DATA_WIDTH = 32;
defparam rnode_230to231_bb4_shr2_i_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_shr2_i_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_shr2_i_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr2_i_stall_in = 1'b0;
assign rnode_230to231_bb4_shr2_i_0_NO_SHIFT_REG = rnode_230to231_bb4_shr2_i_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_shr2_i_0_stall_in_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_shr2_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_230to231_bb4_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_xor_i195_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_xor_i195_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_xor_i195_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_xor_i195_0_valid_out_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_xor_i195_0_stall_in_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_xor_i195_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_xor_i195_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_xor_i195_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_xor_i195_0_stall_in_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_xor_i195_0_valid_out_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_xor_i195_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in(local_bb4_xor_i195),
	.data_out(rnode_230to231_bb4_xor_i195_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_xor_i195_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_xor_i195_0_reg_231_fifo.DATA_WIDTH = 32;
defparam rnode_230to231_bb4_xor_i195_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_xor_i195_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_xor_i195_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor_i195_stall_in = 1'b0;
assign rnode_230to231_bb4_xor_i195_0_NO_SHIFT_REG = rnode_230to231_bb4_xor_i195_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_xor_i195_0_stall_in_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_and6_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_and6_i_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_and6_i_1_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_and6_i_2_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_and6_i_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_valid_out_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_stall_in_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and6_i_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_and6_i_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_and6_i_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_and6_i_0_stall_in_0_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_and6_i_0_valid_out_0_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_and6_i_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in((local_bb4_and6_i & 32'h7FFFFF)),
	.data_out(rnode_230to231_bb4_and6_i_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_and6_i_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_and6_i_0_reg_231_fifo.DATA_WIDTH = 32;
defparam rnode_230to231_bb4_and6_i_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_and6_i_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_and6_i_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and6_i_stall_in_1 = 1'b0;
assign rnode_230to231_bb4_and6_i_0_stall_in_0_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_and6_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_and6_i_0_NO_SHIFT_REG = rnode_230to231_bb4_and6_i_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_and6_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_and6_i_1_NO_SHIFT_REG = rnode_230to231_bb4_and6_i_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_and6_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_and6_i_2_NO_SHIFT_REG = rnode_230to231_bb4_and6_i_0_reg_231_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_var__u65_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_var__u65_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_var__u65_1_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_var__u65_2_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_var__u65_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_valid_out_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_stall_in_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_var__u65_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_var__u65_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_var__u65_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_var__u65_0_stall_in_0_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_var__u65_0_valid_out_0_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_var__u65_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in(local_bb4_var__u65),
	.data_out(rnode_230to231_bb4_var__u65_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_var__u65_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_var__u65_0_reg_231_fifo.DATA_WIDTH = 32;
defparam rnode_230to231_bb4_var__u65_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_var__u65_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_var__u65_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u65_stall_in = 1'b0;
assign rnode_230to231_bb4_var__u65_0_stall_in_0_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_var__u65_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_var__u65_0_NO_SHIFT_REG = rnode_230to231_bb4_var__u65_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_var__u65_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_var__u65_1_NO_SHIFT_REG = rnode_230to231_bb4_var__u65_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_var__u65_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_var__u65_2_NO_SHIFT_REG = rnode_230to231_bb4_var__u65_0_reg_231_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_shr_i193_0_valid_out_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr_i193_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_shr_i193_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr_i193_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_shr_i193_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr_i193_0_valid_out_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr_i193_0_stall_in_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_shr_i193_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_shr_i193_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_shr_i193_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_shr_i193_0_stall_in_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_shr_i193_0_valid_out_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_shr_i193_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in((local_bb4_shr_i193 & 32'h1FF)),
	.data_out(rnode_230to231_bb4_shr_i193_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_shr_i193_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_shr_i193_0_reg_231_fifo.DATA_WIDTH = 32;
defparam rnode_230to231_bb4_shr_i193_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_shr_i193_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_shr_i193_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr_i193_stall_in = 1'b0;
assign rnode_230to231_bb4_shr_i193_0_NO_SHIFT_REG = rnode_230to231_bb4_shr_i193_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_shr_i193_0_stall_in_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_shr_i193_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_230to231_bb4_and5_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and5_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_and5_i_0_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and5_i_0_reg_231_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_230to231_bb4_and5_i_0_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and5_i_0_valid_out_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and5_i_0_stall_in_reg_231_NO_SHIFT_REG;
 logic rnode_230to231_bb4_and5_i_0_stall_out_reg_231_NO_SHIFT_REG;

acl_data_fifo rnode_230to231_bb4_and5_i_0_reg_231_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_230to231_bb4_and5_i_0_reg_231_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_230to231_bb4_and5_i_0_stall_in_reg_231_NO_SHIFT_REG),
	.valid_out(rnode_230to231_bb4_and5_i_0_valid_out_reg_231_NO_SHIFT_REG),
	.stall_out(rnode_230to231_bb4_and5_i_0_stall_out_reg_231_NO_SHIFT_REG),
	.data_in((local_bb4_and5_i & 32'h7FFFFF)),
	.data_out(rnode_230to231_bb4_and5_i_0_reg_231_NO_SHIFT_REG)
);

defparam rnode_230to231_bb4_and5_i_0_reg_231_fifo.DEPTH = 1;
defparam rnode_230to231_bb4_and5_i_0_reg_231_fifo.DATA_WIDTH = 32;
defparam rnode_230to231_bb4_and5_i_0_reg_231_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_230to231_bb4_and5_i_0_reg_231_fifo.IMPL = "shift_reg";

assign rnode_230to231_bb4_and5_i_0_reg_231_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and5_i_stall_in_1 = 1'b0;
assign rnode_230to231_bb4_and5_i_0_NO_SHIFT_REG = rnode_230to231_bb4_and5_i_0_reg_231_NO_SHIFT_REG;
assign rnode_230to231_bb4_and5_i_0_stall_in_reg_231_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_and5_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb4_mul_i_i_inputs_ready;
 reg local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG;
wire local_bb4_mul_i_i_stall_in_0;
 reg local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i_stall_in_1;
wire local_bb4_mul_i_i_output_regs_ready;
wire [63:0] local_bb4_mul_i_i;
 reg local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb4_mul_i_i_valid_pipe_1_NO_SHIFT_REG;
wire local_bb4_mul_i_i_causedstall;

acl_int_mult int_module_local_bb4_mul_i_i (
	.clock(clock),
	.dataa(((local_bb4_conv1_i_i & 64'hFFFFFF) | 64'h800000)),
	.datab(((local_bb4_conv_i_i & 64'hFFFFFF) | 64'h800000)),
	.enable(local_bb4_mul_i_i_output_regs_ready),
	.result(local_bb4_mul_i_i)
);

defparam int_module_local_bb4_mul_i_i.INPUT1_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i.INPUT2_WIDTH = 24;
defparam int_module_local_bb4_mul_i_i.OUTPUT_WIDTH = 64;
defparam int_module_local_bb4_mul_i_i.LATENCY = 3;
defparam int_module_local_bb4_mul_i_i.SIGNED = 0;

assign local_bb4_mul_i_i_inputs_ready = 1'b1;
assign local_bb4_mul_i_i_output_regs_ready = 1'b1;
assign local_bb4_conv1_i_i_stall_in = 1'b0;
assign local_bb4_conv_i_i_stall_in = 1'b0;
assign local_bb4_mul_i_i_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i_output_regs_ready)
		begin
			local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= local_bb4_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_mul_i_i_output_regs_ready)
		begin
			local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_mul_i_i_stall_in_0))
			begin
				local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb4_mul_i_i_stall_in_1))
			begin
				local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_and3_i_stall_local;
wire [31:0] local_bb4_and3_i;

assign local_bb4_and3_i = ((rnode_230to231_bb4_shr2_i_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_231to234_bb4_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_231to234_bb4_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_231to234_bb4_xor_i195_0_NO_SHIFT_REG;
 logic rnode_231to234_bb4_xor_i195_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_231to234_bb4_xor_i195_0_reg_234_NO_SHIFT_REG;
 logic rnode_231to234_bb4_xor_i195_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_231to234_bb4_xor_i195_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_231to234_bb4_xor_i195_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_231to234_bb4_xor_i195_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to234_bb4_xor_i195_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to234_bb4_xor_i195_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_231to234_bb4_xor_i195_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_231to234_bb4_xor_i195_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(rnode_230to231_bb4_xor_i195_0_NO_SHIFT_REG),
	.data_out(rnode_231to234_bb4_xor_i195_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_231to234_bb4_xor_i195_0_reg_234_fifo.DEPTH = 3;
defparam rnode_231to234_bb4_xor_i195_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_231to234_bb4_xor_i195_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to234_bb4_xor_i195_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_231to234_bb4_xor_i195_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_231to234_bb4_xor_i195_0_NO_SHIFT_REG = rnode_231to234_bb4_xor_i195_0_reg_234_NO_SHIFT_REG;
assign rnode_231to234_bb4_xor_i195_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_231to234_bb4_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_i_stall_local;
wire local_bb4_lnot17_i;

assign local_bb4_lnot17_i = ((rnode_230to231_bb4_and6_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_stall_local;
wire [31:0] local_bb4_and_i;

assign local_bb4_and_i = (rnode_230to231_bb4_var__u65_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i_stall_local;
wire [31:0] local_bb4_and10_i;

assign local_bb4_and10_i = (rnode_230to231_bb4_var__u65_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_231to232_bb4_var__u65_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u65_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_var__u65_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u65_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u65_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_var__u65_1_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u65_0_reg_232_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_var__u65_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u65_0_valid_out_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u65_0_stall_in_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u65_0_stall_out_reg_232_NO_SHIFT_REG;

acl_data_fifo rnode_231to232_bb4_var__u65_0_reg_232_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to232_bb4_var__u65_0_reg_232_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to232_bb4_var__u65_0_stall_in_0_reg_232_NO_SHIFT_REG),
	.valid_out(rnode_231to232_bb4_var__u65_0_valid_out_0_reg_232_NO_SHIFT_REG),
	.stall_out(rnode_231to232_bb4_var__u65_0_stall_out_reg_232_NO_SHIFT_REG),
	.data_in(rnode_230to231_bb4_var__u65_2_NO_SHIFT_REG),
	.data_out(rnode_231to232_bb4_var__u65_0_reg_232_NO_SHIFT_REG)
);

defparam rnode_231to232_bb4_var__u65_0_reg_232_fifo.DEPTH = 1;
defparam rnode_231to232_bb4_var__u65_0_reg_232_fifo.DATA_WIDTH = 32;
defparam rnode_231to232_bb4_var__u65_0_reg_232_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to232_bb4_var__u65_0_reg_232_fifo.IMPL = "shift_reg";

assign rnode_231to232_bb4_var__u65_0_reg_232_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_230to231_bb4_var__u65_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u65_0_stall_in_0_reg_232_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u65_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4_var__u65_0_NO_SHIFT_REG = rnode_231to232_bb4_var__u65_0_reg_232_NO_SHIFT_REG;
assign rnode_231to232_bb4_var__u65_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4_var__u65_1_NO_SHIFT_REG = rnode_231to232_bb4_var__u65_0_reg_232_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i194_stall_local;
wire [31:0] local_bb4_and_i194;

assign local_bb4_and_i194 = ((rnode_230to231_bb4_shr_i193_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_i_stall_local;
wire local_bb4_lnot14_i;

assign local_bb4_lnot14_i = ((rnode_230to231_bb4_and5_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_conv3_i_i_stall_local;
wire [31:0] local_bb4_conv3_i_i;
wire [63:0] local_bb4_conv3_i_i$ps;

assign local_bb4_conv3_i_i$ps = (local_bb4_mul_i_i & 64'hFFFFFFFFFFFF);
assign local_bb4_conv3_i_i = local_bb4_conv3_i_i$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_var__u66_stall_local;
wire [63:0] local_bb4_var__u66;

assign local_bb4_var__u66 = ((local_bb4_mul_i_i & 64'hFFFFFFFFFFFF) >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot8_i_stall_local;
wire local_bb4_lnot8_i;

assign local_bb4_lnot8_i = ((local_bb4_and3_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_i_stall_local;
wire local_bb4_cmp11_i;

assign local_bb4_cmp11_i = ((local_bb4_and3_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u67_stall_local;
wire [31:0] local_bb4_var__u67;

assign local_bb4_var__u67 = ((local_bb4_and3_i & 32'hFF) | (rnode_230to231_bb4_and6_i_1_NO_SHIFT_REG & 32'h7FFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_xor_i195_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_xor_i195_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_xor_i195_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_xor_i195_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_xor_i195_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_xor_i195_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_xor_i195_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_xor_i195_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_xor_i195_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_xor_i195_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_xor_i195_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_xor_i195_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_xor_i195_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(rnode_231to234_bb4_xor_i195_0_NO_SHIFT_REG),
	.data_out(rnode_234to235_bb4_xor_i195_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_xor_i195_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_xor_i195_0_reg_235_fifo.DATA_WIDTH = 32;
defparam rnode_234to235_bb4_xor_i195_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_xor_i195_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_xor_i195_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_231to234_bb4_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_xor_i195_0_NO_SHIFT_REG = rnode_234to235_bb4_xor_i195_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_xor_i195_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_xor_i195_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot17_not_i_stall_local;
wire local_bb4_lnot17_not_i;

assign local_bb4_lnot17_not_i = (local_bb4_lnot17_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i1_stall_local;
wire [31:0] local_bb4_shr_i1;

assign local_bb4_shr_i1 = ((local_bb4_and_i & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i_stall_local;
wire local_bb4_cmp13_i;

assign local_bb4_cmp13_i = ((local_bb4_and10_i & 32'hFFFF) > (local_bb4_and12_i & 32'hFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i196_stall_local;
wire local_bb4_lnot_i196;

assign local_bb4_lnot_i196 = ((local_bb4_and_i194 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i197_stall_local;
wire local_bb4_cmp_i197;

assign local_bb4_cmp_i197 = ((local_bb4_and_i194 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u68_stall_local;
wire [31:0] local_bb4_var__u68;

assign local_bb4_var__u68 = ((rnode_230to231_bb4_and6_i_2_NO_SHIFT_REG & 32'h7FFFFF) | (local_bb4_and_i194 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_add_i206_stall_local;
wire [31:0] local_bb4_add_i206;

assign local_bb4_add_i206 = ((local_bb4_and3_i & 32'hFF) + (local_bb4_and_i194 & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot14_not_i_stall_local;
wire local_bb4_lnot14_not_i;

assign local_bb4_lnot14_not_i = (local_bb4_lnot14_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i16_i_stall_local;
wire [31:0] local_bb4_shr_i16_i;

assign local_bb4_shr_i16_i = (local_bb4_conv3_i_i >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i18_i_stall_local;
wire [31:0] local_bb4_shl1_i18_i;

assign local_bb4_shl1_i18_i = (local_bb4_conv3_i_i << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u69_stall_local;
wire [31:0] local_bb4_var__u69;

assign local_bb4_var__u69 = (local_bb4_conv3_i_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shl1_i_i_stall_local;
wire [31:0] local_bb4_shl1_i_i;

assign local_bb4_shl1_i_i = (local_bb4_conv3_i_i << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb4__tr_i_stall_local;
wire [31:0] local_bb4__tr_i;
wire [63:0] local_bb4__tr_i$ps;

assign local_bb4__tr_i$ps = (local_bb4_var__u66 & 64'hFFFFFF);
assign local_bb4__tr_i = local_bb4__tr_i$ps[31:0];

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge8_demorgan_i_stall_local;
wire local_bb4_brmerge8_demorgan_i;

assign local_bb4_brmerge8_demorgan_i = (local_bb4_cmp11_i & local_bb4_lnot17_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp11_not_i_stall_local;
wire local_bb4_cmp11_not_i;

assign local_bb4_cmp11_not_i = (local_bb4_cmp11_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u70_stall_local;
wire local_bb4_var__u70;

assign local_bb4_var__u70 = ((local_bb4_var__u67 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and4_i_stall_local;
wire [31:0] local_bb4_and4_i;

assign local_bb4_and4_i = (rnode_234to235_bb4_xor_i195_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i3_stall_local;
wire local_bb4_cmp_i3;

assign local_bb4_cmp_i3 = ((local_bb4_shr_i1 & 32'h7FFF) > (local_bb4_shr3_i & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i_stall_local;
wire local_bb4_cmp8_i;

assign local_bb4_cmp8_i = ((local_bb4_shr_i1 & 32'h7FFF) == (local_bb4_shr3_i & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i212_stall_local;
wire local_bb4_reduction_0_i212;

assign local_bb4_reduction_0_i212 = (local_bb4_lnot_i196 | local_bb4_lnot8_i);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u71_stall_local;
wire local_bb4_var__u71;

assign local_bb4_var__u71 = (local_bb4_cmp_i197 | local_bb4_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u72_stall_local;
wire local_bb4_var__u72;

assign local_bb4_var__u72 = ((local_bb4_var__u68 & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__28_i203_stall_local;
wire local_bb4__28_i203;

assign local_bb4__28_i203 = (local_bb4_cmp_i197 & local_bb4_lnot14_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i207_stall_local;
wire [31:0] local_bb4_shr_i_i207;

assign local_bb4_shr_i_i207 = ((local_bb4_var__u69 & 32'h1FF) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i15_i_stall_local;
wire [31:0] local_bb4_shl_i15_i;

assign local_bb4_shl_i15_i = ((local_bb4__tr_i & 32'hFFFFFF) & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb4_and48_i_stall_local;
wire [31:0] local_bb4_and48_i;

assign local_bb4_and48_i = ((local_bb4__tr_i & 32'hFFFFFF) & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge10_demorgan_i_stall_local;
wire local_bb4_brmerge10_demorgan_i;

assign local_bb4_brmerge10_demorgan_i = (local_bb4_brmerge8_demorgan_i & local_bb4_lnot_i196);

// This section implements an unregistered operation.
// 
wire local_bb4__mux9_mux_i_stall_local;
wire local_bb4__mux9_mux_i;

assign local_bb4__mux9_mux_i = (local_bb4_brmerge8_demorgan_i ^ local_bb4_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge3_i_stall_local;
wire local_bb4_brmerge3_i;

assign local_bb4_brmerge3_i = (local_bb4_var__u70 | local_bb4_cmp11_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_i_stall_local;
wire local_bb4__mux_mux_i;

assign local_bb4__mux_mux_i = (local_bb4_var__u70 | local_bb4_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb4__not_i_stall_local;
wire local_bb4__not_i;

assign local_bb4__not_i = (local_bb4_var__u70 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4___i4_stall_local;
wire local_bb4___i4;

assign local_bb4___i4 = (local_bb4_cmp8_i & local_bb4_cmp13_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i17_i_stall_local;
wire [31:0] local_bb4_or_i17_i;

assign local_bb4_or_i17_i = ((local_bb4_shl_i15_i & 32'hFFFF00) | (local_bb4_shr_i16_i & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool49_i_stall_local;
wire local_bb4_tobool49_i;

assign local_bb4_tobool49_i = ((local_bb4_and48_i & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4__26_demorgan_i_stall_local;
wire local_bb4__26_demorgan_i;

assign local_bb4__26_demorgan_i = (local_bb4_cmp_i197 | local_bb4_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge5_i_stall_local;
wire local_bb4_brmerge5_i;

assign local_bb4_brmerge5_i = (local_bb4_brmerge3_i | local_bb4_lnot17_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i198_stall_local;
wire local_bb4_reduction_3_i198;

assign local_bb4_reduction_3_i198 = (local_bb4_cmp11_i & local_bb4__not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u45_valid_out_2;
wire local_bb4_var__u45_stall_in_2;
wire local_bb4__21_i_valid_out;
wire local_bb4__21_i_stall_in;
wire local_bb4__21_i_inputs_ready;
wire local_bb4__21_i_stall_local;
wire local_bb4__21_i;

assign local_bb4__21_i_inputs_ready = (rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_valid_out_0_NO_SHIFT_REG & rnode_230to231_bb4_var__u65_0_valid_out_1_NO_SHIFT_REG & rnode_230to231_bb4_var__u65_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__21_i = (local_bb4_cmp_i3 | local_bb4___i4);
assign local_bb4_var__u45_valid_out_2 = 1'b1;
assign local_bb4__21_i_valid_out = 1'b1;
assign rnode_230to231_bb4_sum_321_pop9_c1_ene5_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_var__u65_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_var__u65_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i_i_stall_local;
wire [31:0] local_bb4_shl_i_i;

assign local_bb4_shl_i_i = ((local_bb4_or_i17_i & 32'hFFFFFF) << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__mux_mux_mux_i_stall_local;
wire local_bb4__mux_mux_mux_i;

assign local_bb4__mux_mux_mux_i = (local_bb4_brmerge5_i & local_bb4__mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i199_stall_local;
wire local_bb4_reduction_5_i199;

assign local_bb4_reduction_5_i199 = (local_bb4_lnot14_i & local_bb4_reduction_3_i198);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_231to232_bb4_var__u45_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u45_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_var__u45_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u45_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u45_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_var__u45_1_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u45_0_reg_232_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_231to232_bb4_var__u45_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u45_0_valid_out_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u45_0_stall_in_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u45_0_stall_out_reg_232_NO_SHIFT_REG;

acl_data_fifo rnode_231to232_bb4_var__u45_0_reg_232_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to232_bb4_var__u45_0_reg_232_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to232_bb4_var__u45_0_stall_in_0_reg_232_NO_SHIFT_REG),
	.valid_out(rnode_231to232_bb4_var__u45_0_valid_out_0_reg_232_NO_SHIFT_REG),
	.stall_out(rnode_231to232_bb4_var__u45_0_stall_out_reg_232_NO_SHIFT_REG),
	.data_in(local_bb4_var__u45),
	.data_out(rnode_231to232_bb4_var__u45_0_reg_232_NO_SHIFT_REG)
);

defparam rnode_231to232_bb4_var__u45_0_reg_232_fifo.DEPTH = 1;
defparam rnode_231to232_bb4_var__u45_0_reg_232_fifo.DATA_WIDTH = 32;
defparam rnode_231to232_bb4_var__u45_0_reg_232_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to232_bb4_var__u45_0_reg_232_fifo.IMPL = "shift_reg";

assign rnode_231to232_bb4_var__u45_0_reg_232_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u45_stall_in_2 = 1'b0;
assign rnode_231to232_bb4_var__u45_0_stall_in_0_reg_232_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u45_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4_var__u45_0_NO_SHIFT_REG = rnode_231to232_bb4_var__u45_0_reg_232_NO_SHIFT_REG;
assign rnode_231to232_bb4_var__u45_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4_var__u45_1_NO_SHIFT_REG = rnode_231to232_bb4_var__u45_0_reg_232_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_231to232_bb4__21_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_1_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_reg_232_inputs_ready_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_valid_out_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_stall_in_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4__21_i_0_stall_out_reg_232_NO_SHIFT_REG;

acl_data_fifo rnode_231to232_bb4__21_i_0_reg_232_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to232_bb4__21_i_0_reg_232_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to232_bb4__21_i_0_stall_in_0_reg_232_NO_SHIFT_REG),
	.valid_out(rnode_231to232_bb4__21_i_0_valid_out_0_reg_232_NO_SHIFT_REG),
	.stall_out(rnode_231to232_bb4__21_i_0_stall_out_reg_232_NO_SHIFT_REG),
	.data_in(local_bb4__21_i),
	.data_out(rnode_231to232_bb4__21_i_0_reg_232_NO_SHIFT_REG)
);

defparam rnode_231to232_bb4__21_i_0_reg_232_fifo.DEPTH = 1;
defparam rnode_231to232_bb4__21_i_0_reg_232_fifo.DATA_WIDTH = 1;
defparam rnode_231to232_bb4__21_i_0_reg_232_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to232_bb4__21_i_0_reg_232_fifo.IMPL = "shift_reg";

assign rnode_231to232_bb4__21_i_0_reg_232_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i_stall_in = 1'b0;
assign rnode_231to232_bb4__21_i_0_stall_in_0_reg_232_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4__21_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4__21_i_0_NO_SHIFT_REG = rnode_231to232_bb4__21_i_0_reg_232_NO_SHIFT_REG;
assign rnode_231to232_bb4__21_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4__21_i_1_NO_SHIFT_REG = rnode_231to232_bb4__21_i_0_reg_232_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i208_stall_local;
wire [31:0] local_bb4_or_i_i208;

assign local_bb4_or_i_i208 = ((local_bb4_shl_i_i & 32'h1FFFFFE) | (local_bb4_shr_i_i207 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i200_stall_local;
wire local_bb4_reduction_6_i200;

assign local_bb4_reduction_6_i200 = (local_bb4_var__u72 & local_bb4_reduction_5_i199);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i_stall_local;
wire [31:0] local_bb4__22_i;

assign local_bb4__22_i = (rnode_231to232_bb4__21_i_0_NO_SHIFT_REG ? rnode_231to232_bb4_var__u45_0_NO_SHIFT_REG : rnode_231to232_bb4_var__u65_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i_stall_local;
wire [31:0] local_bb4__23_i;

assign local_bb4__23_i = (rnode_231to232_bb4__21_i_1_NO_SHIFT_REG ? rnode_231to232_bb4_var__u65_1_NO_SHIFT_REG : rnode_231to232_bb4_var__u45_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i201_stall_local;
wire local_bb4__24_i201;

assign local_bb4__24_i201 = (local_bb4_cmp_i197 ? local_bb4_reduction_6_i200 : local_bb4_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i_stall_local;
wire [31:0] local_bb4_shr18_i;

assign local_bb4_shr18_i = (local_bb4__22_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i_stall_local;
wire [31:0] local_bb4_shr16_i;

assign local_bb4_shr16_i = (local_bb4__23_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4__25_i_stall_local;
wire local_bb4__25_i;

assign local_bb4__25_i = (local_bb4__24_i201 ? local_bb4_lnot14_i : local_bb4__mux_mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i_stall_local;
wire [31:0] local_bb4_and19_i;

assign local_bb4_and19_i = ((local_bb4_shr18_i & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i_stall_local;
wire [31:0] local_bb4_sub_i;

assign local_bb4_sub_i = ((local_bb4_shr16_i & 32'h1FF) - (local_bb4_shr18_i & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4__27_i202_stall_local;
wire local_bb4__27_i202;

assign local_bb4__27_i202 = (local_bb4__26_demorgan_i ? local_bb4__25_i : local_bb4__mux9_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i_stall_local;
wire local_bb4_lnot23_i;

assign local_bb4_lnot23_i = ((local_bb4_and19_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i_stall_local;
wire local_bb4_cmp27_i;

assign local_bb4_cmp27_i = ((local_bb4_and19_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and68_i_stall_local;
wire [31:0] local_bb4_and68_i;

assign local_bb4_and68_i = (local_bb4_sub_i & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_add_i206_valid_out;
wire local_bb4_add_i206_stall_in;
wire local_bb4_reduction_0_i212_valid_out;
wire local_bb4_reduction_0_i212_stall_in;
wire local_bb4_var__u71_valid_out;
wire local_bb4_var__u71_stall_in;
wire local_bb4__29_i204_valid_out;
wire local_bb4__29_i204_stall_in;
wire local_bb4__29_i204_inputs_ready;
wire local_bb4__29_i204_stall_local;
wire local_bb4__29_i204;

assign local_bb4__29_i204_inputs_ready = (rnode_230to231_bb4_shr2_i_0_valid_out_NO_SHIFT_REG & rnode_230to231_bb4_and6_i_0_valid_out_1_NO_SHIFT_REG & rnode_230to231_bb4_and6_i_0_valid_out_0_NO_SHIFT_REG & rnode_230to231_bb4_and6_i_0_valid_out_2_NO_SHIFT_REG & rnode_230to231_bb4_shr_i193_0_valid_out_NO_SHIFT_REG & rnode_230to231_bb4_and5_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4__29_i204 = (local_bb4__28_i203 | local_bb4__27_i202);
assign local_bb4_add_i206_valid_out = 1'b1;
assign local_bb4_reduction_0_i212_valid_out = 1'b1;
assign local_bb4_var__u71_valid_out = 1'b1;
assign local_bb4__29_i204_valid_out = 1'b1;
assign rnode_230to231_bb4_shr2_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_and6_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_and6_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_and6_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_shr_i193_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_230to231_bb4_and5_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp69_i_stall_local;
wire local_bb4_cmp69_i;

assign local_bb4_cmp69_i = ((local_bb4_and68_i & 32'hFF) > 32'h1F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_231to233_bb4_add_i206_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_231to233_bb4_add_i206_0_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_231to233_bb4_add_i206_1_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_231to233_bb4_add_i206_2_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_reg_233_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_231to233_bb4_add_i206_0_reg_233_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_valid_out_0_reg_233_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_stall_in_0_reg_233_NO_SHIFT_REG;
 logic rnode_231to233_bb4_add_i206_0_stall_out_reg_233_NO_SHIFT_REG;

acl_data_fifo rnode_231to233_bb4_add_i206_0_reg_233_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to233_bb4_add_i206_0_reg_233_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to233_bb4_add_i206_0_stall_in_0_reg_233_NO_SHIFT_REG),
	.valid_out(rnode_231to233_bb4_add_i206_0_valid_out_0_reg_233_NO_SHIFT_REG),
	.stall_out(rnode_231to233_bb4_add_i206_0_stall_out_reg_233_NO_SHIFT_REG),
	.data_in((local_bb4_add_i206 & 32'h1FF)),
	.data_out(rnode_231to233_bb4_add_i206_0_reg_233_NO_SHIFT_REG)
);

defparam rnode_231to233_bb4_add_i206_0_reg_233_fifo.DEPTH = 2;
defparam rnode_231to233_bb4_add_i206_0_reg_233_fifo.DATA_WIDTH = 32;
defparam rnode_231to233_bb4_add_i206_0_reg_233_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to233_bb4_add_i206_0_reg_233_fifo.IMPL = "shift_reg";

assign rnode_231to233_bb4_add_i206_0_reg_233_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add_i206_stall_in = 1'b0;
assign rnode_231to233_bb4_add_i206_0_stall_in_0_reg_233_NO_SHIFT_REG = 1'b0;
assign rnode_231to233_bb4_add_i206_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_231to233_bb4_add_i206_0_NO_SHIFT_REG = rnode_231to233_bb4_add_i206_0_reg_233_NO_SHIFT_REG;
assign rnode_231to233_bb4_add_i206_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_231to233_bb4_add_i206_1_NO_SHIFT_REG = rnode_231to233_bb4_add_i206_0_reg_233_NO_SHIFT_REG;
assign rnode_231to233_bb4_add_i206_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_231to233_bb4_add_i206_2_NO_SHIFT_REG = rnode_231to233_bb4_add_i206_0_reg_233_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_231to232_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_231to232_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_231to232_bb4_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4_reduction_0_i212_0_reg_232_inputs_ready_NO_SHIFT_REG;
 logic rnode_231to232_bb4_reduction_0_i212_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_reduction_0_i212_0_valid_out_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_reduction_0_i212_0_stall_in_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_reduction_0_i212_0_stall_out_reg_232_NO_SHIFT_REG;

acl_data_fifo rnode_231to232_bb4_reduction_0_i212_0_reg_232_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to232_bb4_reduction_0_i212_0_reg_232_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to232_bb4_reduction_0_i212_0_stall_in_reg_232_NO_SHIFT_REG),
	.valid_out(rnode_231to232_bb4_reduction_0_i212_0_valid_out_reg_232_NO_SHIFT_REG),
	.stall_out(rnode_231to232_bb4_reduction_0_i212_0_stall_out_reg_232_NO_SHIFT_REG),
	.data_in(local_bb4_reduction_0_i212),
	.data_out(rnode_231to232_bb4_reduction_0_i212_0_reg_232_NO_SHIFT_REG)
);

defparam rnode_231to232_bb4_reduction_0_i212_0_reg_232_fifo.DEPTH = 1;
defparam rnode_231to232_bb4_reduction_0_i212_0_reg_232_fifo.DATA_WIDTH = 1;
defparam rnode_231to232_bb4_reduction_0_i212_0_reg_232_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to232_bb4_reduction_0_i212_0_reg_232_fifo.IMPL = "shift_reg";

assign rnode_231to232_bb4_reduction_0_i212_0_reg_232_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_reduction_0_i212_stall_in = 1'b0;
assign rnode_231to232_bb4_reduction_0_i212_0_NO_SHIFT_REG = rnode_231to232_bb4_reduction_0_i212_0_reg_232_NO_SHIFT_REG;
assign rnode_231to232_bb4_reduction_0_i212_0_stall_in_reg_232_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_231to232_bb4_var__u71_0_valid_out_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u71_0_stall_in_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u71_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u71_0_reg_232_inputs_ready_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u71_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u71_0_valid_out_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u71_0_stall_in_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4_var__u71_0_stall_out_reg_232_NO_SHIFT_REG;

acl_data_fifo rnode_231to232_bb4_var__u71_0_reg_232_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to232_bb4_var__u71_0_reg_232_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to232_bb4_var__u71_0_stall_in_reg_232_NO_SHIFT_REG),
	.valid_out(rnode_231to232_bb4_var__u71_0_valid_out_reg_232_NO_SHIFT_REG),
	.stall_out(rnode_231to232_bb4_var__u71_0_stall_out_reg_232_NO_SHIFT_REG),
	.data_in(local_bb4_var__u71),
	.data_out(rnode_231to232_bb4_var__u71_0_reg_232_NO_SHIFT_REG)
);

defparam rnode_231to232_bb4_var__u71_0_reg_232_fifo.DEPTH = 1;
defparam rnode_231to232_bb4_var__u71_0_reg_232_fifo.DATA_WIDTH = 1;
defparam rnode_231to232_bb4_var__u71_0_reg_232_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to232_bb4_var__u71_0_reg_232_fifo.IMPL = "shift_reg";

assign rnode_231to232_bb4_var__u71_0_reg_232_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u71_stall_in = 1'b0;
assign rnode_231to232_bb4_var__u71_0_NO_SHIFT_REG = rnode_231to232_bb4_var__u71_0_reg_232_NO_SHIFT_REG;
assign rnode_231to232_bb4_var__u71_0_stall_in_reg_232_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u71_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_231to232_bb4__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_231to232_bb4__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_231to232_bb4__29_i204_0_NO_SHIFT_REG;
 logic rnode_231to232_bb4__29_i204_0_reg_232_inputs_ready_NO_SHIFT_REG;
 logic rnode_231to232_bb4__29_i204_0_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4__29_i204_0_valid_out_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4__29_i204_0_stall_in_reg_232_NO_SHIFT_REG;
 logic rnode_231to232_bb4__29_i204_0_stall_out_reg_232_NO_SHIFT_REG;

acl_data_fifo rnode_231to232_bb4__29_i204_0_reg_232_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_231to232_bb4__29_i204_0_reg_232_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_231to232_bb4__29_i204_0_stall_in_reg_232_NO_SHIFT_REG),
	.valid_out(rnode_231to232_bb4__29_i204_0_valid_out_reg_232_NO_SHIFT_REG),
	.stall_out(rnode_231to232_bb4__29_i204_0_stall_out_reg_232_NO_SHIFT_REG),
	.data_in(local_bb4__29_i204),
	.data_out(rnode_231to232_bb4__29_i204_0_reg_232_NO_SHIFT_REG)
);

defparam rnode_231to232_bb4__29_i204_0_reg_232_fifo.DEPTH = 1;
defparam rnode_231to232_bb4__29_i204_0_reg_232_fifo.DATA_WIDTH = 1;
defparam rnode_231to232_bb4__29_i204_0_reg_232_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_231to232_bb4__29_i204_0_reg_232_fifo.IMPL = "shift_reg";

assign rnode_231to232_bb4__29_i204_0_reg_232_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__29_i204_stall_in = 1'b0;
assign rnode_231to232_bb4__29_i204_0_NO_SHIFT_REG = rnode_231to232_bb4__29_i204_0_reg_232_NO_SHIFT_REG;
assign rnode_231to232_bb4__29_i204_0_stall_in_reg_232_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__22_i_valid_out_1;
wire local_bb4__22_i_stall_in_1;
wire local_bb4__23_i_valid_out_1;
wire local_bb4__23_i_stall_in_1;
wire local_bb4_shr16_i_valid_out_1;
wire local_bb4_shr16_i_stall_in_1;
wire local_bb4_lnot23_i_valid_out;
wire local_bb4_lnot23_i_stall_in;
wire local_bb4_cmp27_i_valid_out;
wire local_bb4_cmp27_i_stall_in;
wire local_bb4_align_0_i_valid_out;
wire local_bb4_align_0_i_stall_in;
wire local_bb4_align_0_i_inputs_ready;
wire local_bb4_align_0_i_stall_local;
wire [31:0] local_bb4_align_0_i;

assign local_bb4_align_0_i_inputs_ready = (rnode_231to232_bb4__21_i_0_valid_out_0_NO_SHIFT_REG & rnode_231to232_bb4_var__u45_0_valid_out_0_NO_SHIFT_REG & rnode_231to232_bb4_var__u65_0_valid_out_0_NO_SHIFT_REG & rnode_231to232_bb4__21_i_0_valid_out_1_NO_SHIFT_REG & rnode_231to232_bb4_var__u45_0_valid_out_1_NO_SHIFT_REG & rnode_231to232_bb4_var__u65_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_align_0_i = (local_bb4_cmp69_i ? 32'h1F : (local_bb4_and68_i & 32'hFF));
assign local_bb4__22_i_valid_out_1 = 1'b1;
assign local_bb4__23_i_valid_out_1 = 1'b1;
assign local_bb4_shr16_i_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i_valid_out = 1'b1;
assign local_bb4_cmp27_i_valid_out = 1'b1;
assign local_bb4_align_0_i_valid_out = 1'b1;
assign rnode_231to232_bb4__21_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u45_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u65_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4__21_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u45_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_231to232_bb4_var__u65_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_inc_i_stall_local;
wire [31:0] local_bb4_inc_i;

assign local_bb4_inc_i = ((rnode_231to233_bb4_add_i206_0_NO_SHIFT_REG & 32'h1FF) + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp50_not_i_stall_local;
wire local_bb4_cmp50_not_i;

assign local_bb4_cmp50_not_i = ((rnode_231to233_bb4_add_i206_1_NO_SHIFT_REG & 32'h1FF) != 32'h7F);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_232to234_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_232to234_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_232to234_bb4_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_232to234_bb4_reduction_0_i212_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_232to234_bb4_reduction_0_i212_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_reduction_0_i212_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_reduction_0_i212_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_reduction_0_i212_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_232to234_bb4_reduction_0_i212_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to234_bb4_reduction_0_i212_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to234_bb4_reduction_0_i212_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_232to234_bb4_reduction_0_i212_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_232to234_bb4_reduction_0_i212_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(rnode_231to232_bb4_reduction_0_i212_0_NO_SHIFT_REG),
	.data_out(rnode_232to234_bb4_reduction_0_i212_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_232to234_bb4_reduction_0_i212_0_reg_234_fifo.DEPTH = 2;
defparam rnode_232to234_bb4_reduction_0_i212_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_232to234_bb4_reduction_0_i212_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to234_bb4_reduction_0_i212_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_232to234_bb4_reduction_0_i212_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4_reduction_0_i212_0_NO_SHIFT_REG = rnode_232to234_bb4_reduction_0_i212_0_reg_234_NO_SHIFT_REG;
assign rnode_232to234_bb4_reduction_0_i212_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_232to233_bb4_var__u71_0_valid_out_NO_SHIFT_REG;
 logic rnode_232to233_bb4_var__u71_0_stall_in_NO_SHIFT_REG;
 logic rnode_232to233_bb4_var__u71_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4_var__u71_0_reg_233_inputs_ready_NO_SHIFT_REG;
 logic rnode_232to233_bb4_var__u71_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_var__u71_0_valid_out_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_var__u71_0_stall_in_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_var__u71_0_stall_out_reg_233_NO_SHIFT_REG;

acl_data_fifo rnode_232to233_bb4_var__u71_0_reg_233_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to233_bb4_var__u71_0_reg_233_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to233_bb4_var__u71_0_stall_in_reg_233_NO_SHIFT_REG),
	.valid_out(rnode_232to233_bb4_var__u71_0_valid_out_reg_233_NO_SHIFT_REG),
	.stall_out(rnode_232to233_bb4_var__u71_0_stall_out_reg_233_NO_SHIFT_REG),
	.data_in(rnode_231to232_bb4_var__u71_0_NO_SHIFT_REG),
	.data_out(rnode_232to233_bb4_var__u71_0_reg_233_NO_SHIFT_REG)
);

defparam rnode_232to233_bb4_var__u71_0_reg_233_fifo.DEPTH = 1;
defparam rnode_232to233_bb4_var__u71_0_reg_233_fifo.DATA_WIDTH = 1;
defparam rnode_232to233_bb4_var__u71_0_reg_233_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to233_bb4_var__u71_0_reg_233_fifo.IMPL = "shift_reg";

assign rnode_232to233_bb4_var__u71_0_reg_233_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4_var__u71_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_var__u71_0_NO_SHIFT_REG = rnode_232to233_bb4_var__u71_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4_var__u71_0_stall_in_reg_233_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_var__u71_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_232to234_bb4__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_232to234_bb4__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_232to234_bb4__29_i204_0_NO_SHIFT_REG;
 logic rnode_232to234_bb4__29_i204_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_232to234_bb4__29_i204_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4__29_i204_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4__29_i204_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4__29_i204_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_232to234_bb4__29_i204_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to234_bb4__29_i204_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to234_bb4__29_i204_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_232to234_bb4__29_i204_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_232to234_bb4__29_i204_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(rnode_231to232_bb4__29_i204_0_NO_SHIFT_REG),
	.data_out(rnode_232to234_bb4__29_i204_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_232to234_bb4__29_i204_0_reg_234_fifo.DEPTH = 2;
defparam rnode_232to234_bb4__29_i204_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_232to234_bb4__29_i204_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to234_bb4__29_i204_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_232to234_bb4__29_i204_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_231to232_bb4__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4__29_i204_0_NO_SHIFT_REG = rnode_232to234_bb4__29_i204_0_reg_234_NO_SHIFT_REG;
assign rnode_232to234_bb4__29_i204_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_232to233_bb4__22_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4__22_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4__22_i_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4__22_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_232to233_bb4__22_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4__22_i_1_NO_SHIFT_REG;
 logic rnode_232to233_bb4__22_i_0_reg_233_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4__22_i_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4__22_i_0_valid_out_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4__22_i_0_stall_in_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4__22_i_0_stall_out_reg_233_NO_SHIFT_REG;

acl_data_fifo rnode_232to233_bb4__22_i_0_reg_233_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to233_bb4__22_i_0_reg_233_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to233_bb4__22_i_0_stall_in_0_reg_233_NO_SHIFT_REG),
	.valid_out(rnode_232to233_bb4__22_i_0_valid_out_0_reg_233_NO_SHIFT_REG),
	.stall_out(rnode_232to233_bb4__22_i_0_stall_out_reg_233_NO_SHIFT_REG),
	.data_in(local_bb4__22_i),
	.data_out(rnode_232to233_bb4__22_i_0_reg_233_NO_SHIFT_REG)
);

defparam rnode_232to233_bb4__22_i_0_reg_233_fifo.DEPTH = 1;
defparam rnode_232to233_bb4__22_i_0_reg_233_fifo.DATA_WIDTH = 32;
defparam rnode_232to233_bb4__22_i_0_reg_233_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to233_bb4__22_i_0_reg_233_fifo.IMPL = "shift_reg";

assign rnode_232to233_bb4__22_i_0_reg_233_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i_stall_in_1 = 1'b0;
assign rnode_232to233_bb4__22_i_0_stall_in_0_reg_233_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4__22_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4__22_i_0_NO_SHIFT_REG = rnode_232to233_bb4__22_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4__22_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4__22_i_1_NO_SHIFT_REG = rnode_232to233_bb4__22_i_0_reg_233_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_232to233_bb4__23_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4__23_i_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4__23_i_1_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4__23_i_2_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_reg_233_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4__23_i_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_valid_out_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_stall_in_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4__23_i_0_stall_out_reg_233_NO_SHIFT_REG;

acl_data_fifo rnode_232to233_bb4__23_i_0_reg_233_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to233_bb4__23_i_0_reg_233_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to233_bb4__23_i_0_stall_in_0_reg_233_NO_SHIFT_REG),
	.valid_out(rnode_232to233_bb4__23_i_0_valid_out_0_reg_233_NO_SHIFT_REG),
	.stall_out(rnode_232to233_bb4__23_i_0_stall_out_reg_233_NO_SHIFT_REG),
	.data_in(local_bb4__23_i),
	.data_out(rnode_232to233_bb4__23_i_0_reg_233_NO_SHIFT_REG)
);

defparam rnode_232to233_bb4__23_i_0_reg_233_fifo.DEPTH = 1;
defparam rnode_232to233_bb4__23_i_0_reg_233_fifo.DATA_WIDTH = 32;
defparam rnode_232to233_bb4__23_i_0_reg_233_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to233_bb4__23_i_0_reg_233_fifo.IMPL = "shift_reg";

assign rnode_232to233_bb4__23_i_0_reg_233_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i_stall_in_1 = 1'b0;
assign rnode_232to233_bb4__23_i_0_stall_in_0_reg_233_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4__23_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4__23_i_0_NO_SHIFT_REG = rnode_232to233_bb4__23_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4__23_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4__23_i_1_NO_SHIFT_REG = rnode_232to233_bb4__23_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4__23_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4__23_i_2_NO_SHIFT_REG = rnode_232to233_bb4__23_i_0_reg_233_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_232to234_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_232to234_bb4_shr16_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_232to234_bb4_shr16_i_0_NO_SHIFT_REG;
 logic rnode_232to234_bb4_shr16_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_232to234_bb4_shr16_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_232to234_bb4_shr16_i_1_NO_SHIFT_REG;
 logic rnode_232to234_bb4_shr16_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_232to234_bb4_shr16_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_shr16_i_0_valid_out_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_shr16_i_0_stall_in_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_shr16_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_232to234_bb4_shr16_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to234_bb4_shr16_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to234_bb4_shr16_i_0_stall_in_0_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_232to234_bb4_shr16_i_0_valid_out_0_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_232to234_bb4_shr16_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i & 32'h1FF)),
	.data_out(rnode_232to234_bb4_shr16_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_232to234_bb4_shr16_i_0_reg_234_fifo.DEPTH = 2;
defparam rnode_232to234_bb4_shr16_i_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_232to234_bb4_shr16_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to234_bb4_shr16_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_232to234_bb4_shr16_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i_stall_in_1 = 1'b0;
assign rnode_232to234_bb4_shr16_i_0_stall_in_0_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4_shr16_i_0_NO_SHIFT_REG = rnode_232to234_bb4_shr16_i_0_reg_234_NO_SHIFT_REG;
assign rnode_232to234_bb4_shr16_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4_shr16_i_1_NO_SHIFT_REG = rnode_232to234_bb4_shr16_i_0_reg_234_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_232to233_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_232to233_bb4_lnot23_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_232to233_bb4_lnot23_i_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4_lnot23_i_0_reg_233_inputs_ready_NO_SHIFT_REG;
 logic rnode_232to233_bb4_lnot23_i_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_lnot23_i_0_valid_out_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_lnot23_i_0_stall_in_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_lnot23_i_0_stall_out_reg_233_NO_SHIFT_REG;

acl_data_fifo rnode_232to233_bb4_lnot23_i_0_reg_233_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to233_bb4_lnot23_i_0_reg_233_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to233_bb4_lnot23_i_0_stall_in_reg_233_NO_SHIFT_REG),
	.valid_out(rnode_232to233_bb4_lnot23_i_0_valid_out_reg_233_NO_SHIFT_REG),
	.stall_out(rnode_232to233_bb4_lnot23_i_0_stall_out_reg_233_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i),
	.data_out(rnode_232to233_bb4_lnot23_i_0_reg_233_NO_SHIFT_REG)
);

defparam rnode_232to233_bb4_lnot23_i_0_reg_233_fifo.DEPTH = 1;
defparam rnode_232to233_bb4_lnot23_i_0_reg_233_fifo.DATA_WIDTH = 1;
defparam rnode_232to233_bb4_lnot23_i_0_reg_233_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to233_bb4_lnot23_i_0_reg_233_fifo.IMPL = "shift_reg";

assign rnode_232to233_bb4_lnot23_i_0_reg_233_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i_stall_in = 1'b0;
assign rnode_232to233_bb4_lnot23_i_0_NO_SHIFT_REG = rnode_232to233_bb4_lnot23_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4_lnot23_i_0_stall_in_reg_233_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_232to234_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_1_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_2_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_valid_out_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_stall_in_0_reg_234_NO_SHIFT_REG;
 logic rnode_232to234_bb4_cmp27_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_232to234_bb4_cmp27_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to234_bb4_cmp27_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to234_bb4_cmp27_i_0_stall_in_0_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_232to234_bb4_cmp27_i_0_valid_out_0_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_232to234_bb4_cmp27_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i),
	.data_out(rnode_232to234_bb4_cmp27_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_232to234_bb4_cmp27_i_0_reg_234_fifo.DEPTH = 2;
defparam rnode_232to234_bb4_cmp27_i_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_232to234_bb4_cmp27_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to234_bb4_cmp27_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_232to234_bb4_cmp27_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i_stall_in = 1'b0;
assign rnode_232to234_bb4_cmp27_i_0_stall_in_0_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4_cmp27_i_0_NO_SHIFT_REG = rnode_232to234_bb4_cmp27_i_0_reg_234_NO_SHIFT_REG;
assign rnode_232to234_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4_cmp27_i_1_NO_SHIFT_REG = rnode_232to234_bb4_cmp27_i_0_reg_234_NO_SHIFT_REG;
assign rnode_232to234_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4_cmp27_i_2_NO_SHIFT_REG = rnode_232to234_bb4_cmp27_i_0_reg_234_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_232to233_bb4_align_0_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4_align_0_i_0_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4_align_0_i_1_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4_align_0_i_2_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4_align_0_i_3_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4_align_0_i_4_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_reg_233_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_232to233_bb4_align_0_i_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_valid_out_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_stall_in_0_reg_233_NO_SHIFT_REG;
 logic rnode_232to233_bb4_align_0_i_0_stall_out_reg_233_NO_SHIFT_REG;

acl_data_fifo rnode_232to233_bb4_align_0_i_0_reg_233_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_232to233_bb4_align_0_i_0_reg_233_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_232to233_bb4_align_0_i_0_stall_in_0_reg_233_NO_SHIFT_REG),
	.valid_out(rnode_232to233_bb4_align_0_i_0_valid_out_0_reg_233_NO_SHIFT_REG),
	.stall_out(rnode_232to233_bb4_align_0_i_0_stall_out_reg_233_NO_SHIFT_REG),
	.data_in((local_bb4_align_0_i & 32'hFF)),
	.data_out(rnode_232to233_bb4_align_0_i_0_reg_233_NO_SHIFT_REG)
);

defparam rnode_232to233_bb4_align_0_i_0_reg_233_fifo.DEPTH = 1;
defparam rnode_232to233_bb4_align_0_i_0_reg_233_fifo.DATA_WIDTH = 32;
defparam rnode_232to233_bb4_align_0_i_0_reg_233_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_232to233_bb4_align_0_i_0_reg_233_fifo.IMPL = "shift_reg";

assign rnode_232to233_bb4_align_0_i_0_reg_233_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_align_0_i_stall_in = 1'b0;
assign rnode_232to233_bb4_align_0_i_0_stall_in_0_reg_233_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_align_0_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4_align_0_i_0_NO_SHIFT_REG = rnode_232to233_bb4_align_0_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4_align_0_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4_align_0_i_1_NO_SHIFT_REG = rnode_232to233_bb4_align_0_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4_align_0_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4_align_0_i_2_NO_SHIFT_REG = rnode_232to233_bb4_align_0_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4_align_0_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4_align_0_i_3_NO_SHIFT_REG = rnode_232to233_bb4_align_0_i_0_reg_233_NO_SHIFT_REG;
assign rnode_232to233_bb4_align_0_i_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4_align_0_i_4_NO_SHIFT_REG = rnode_232to233_bb4_align_0_i_0_reg_233_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__31_i209_stall_local;
wire local_bb4__31_i209;

assign local_bb4__31_i209 = (local_bb4_tobool49_i & local_bb4_cmp50_not_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4_reduction_0_i212_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_reduction_0_i212_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4_reduction_0_i212_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_reduction_0_i212_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_reduction_0_i212_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_reduction_0_i212_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_reduction_0_i212_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_reduction_0_i212_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_reduction_0_i212_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_reduction_0_i212_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_reduction_0_i212_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(rnode_232to234_bb4_reduction_0_i212_0_NO_SHIFT_REG),
	.data_out(rnode_234to235_bb4_reduction_0_i212_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_reduction_0_i212_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_reduction_0_i212_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4_reduction_0_i212_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_reduction_0_i212_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_reduction_0_i212_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_reduction_0_i212_0_NO_SHIFT_REG = rnode_234to235_bb4_reduction_0_i212_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_reduction_0_i212_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_var__u71_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to234_bb4_var__u71_0_stall_in_NO_SHIFT_REG;
 logic rnode_233to234_bb4_var__u71_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_var__u71_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_233to234_bb4_var__u71_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_var__u71_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_var__u71_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_var__u71_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_var__u71_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_var__u71_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_var__u71_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_var__u71_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_var__u71_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(rnode_232to233_bb4_var__u71_0_NO_SHIFT_REG),
	.data_out(rnode_233to234_bb4_var__u71_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_var__u71_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_var__u71_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_233to234_bb4_var__u71_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_var__u71_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_var__u71_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_232to233_bb4_var__u71_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_var__u71_0_NO_SHIFT_REG = rnode_233to234_bb4_var__u71_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_var__u71_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_var__u71_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4__29_i204_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4__29_i204_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4__29_i204_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4__29_i204_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4__29_i204_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__29_i204_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__29_i204_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__29_i204_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4__29_i204_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4__29_i204_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4__29_i204_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4__29_i204_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4__29_i204_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(rnode_232to234_bb4__29_i204_0_NO_SHIFT_REG),
	.data_out(rnode_234to235_bb4__29_i204_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4__29_i204_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4__29_i204_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4__29_i204_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4__29_i204_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4__29_i204_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4__29_i204_0_NO_SHIFT_REG = rnode_234to235_bb4__29_i204_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4__29_i204_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4__29_i204_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i_stall_local;
wire [31:0] local_bb4_and21_i;

assign local_bb4_and21_i = (rnode_232to233_bb4__22_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i_valid_out;
wire local_bb4_and20_i_stall_in;
wire local_bb4_and20_i_inputs_ready;
wire local_bb4_and20_i_stall_local;
wire [31:0] local_bb4_and20_i;

assign local_bb4_and20_i_inputs_ready = rnode_232to233_bb4__23_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i = (rnode_232to233_bb4__23_i_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i_valid_out = 1'b1;
assign rnode_232to233_bb4__23_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i_valid_out;
wire local_bb4_and35_i_stall_in;
wire local_bb4_and35_i_inputs_ready;
wire local_bb4_and35_i_stall_local;
wire [31:0] local_bb4_and35_i;

assign local_bb4_and35_i_inputs_ready = rnode_232to233_bb4__23_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i = (rnode_232to233_bb4__23_i_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i_valid_out = 1'b1;
assign rnode_232to233_bb4__23_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i_stall_local;
wire [31:0] local_bb4_xor_i;

assign local_bb4_xor_i = (rnode_232to233_bb4__23_i_2_NO_SHIFT_REG ^ rnode_232to233_bb4__22_i_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i_stall_local;
wire [31:0] local_bb4_and17_i;

assign local_bb4_and17_i = ((rnode_232to234_bb4_shr16_i_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_234to236_bb4_shr16_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to236_bb4_shr16_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_234to236_bb4_shr16_i_0_NO_SHIFT_REG;
 logic rnode_234to236_bb4_shr16_i_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_234to236_bb4_shr16_i_0_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_shr16_i_0_valid_out_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_shr16_i_0_stall_in_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_shr16_i_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_234to236_bb4_shr16_i_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to236_bb4_shr16_i_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to236_bb4_shr16_i_0_stall_in_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_234to236_bb4_shr16_i_0_valid_out_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_234to236_bb4_shr16_i_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in((rnode_232to234_bb4_shr16_i_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_234to236_bb4_shr16_i_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_234to236_bb4_shr16_i_0_reg_236_fifo.DEPTH = 2;
defparam rnode_234to236_bb4_shr16_i_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_234to236_bb4_shr16_i_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to236_bb4_shr16_i_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_234to236_bb4_shr16_i_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_232to234_bb4_shr16_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_shr16_i_0_NO_SHIFT_REG = rnode_234to236_bb4_shr16_i_0_reg_236_NO_SHIFT_REG;
assign rnode_234to236_bb4_shr16_i_0_stall_in_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_shr16_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and93_i_stall_local;
wire [31:0] local_bb4_and93_i;

assign local_bb4_and93_i = ((rnode_232to233_bb4_align_0_i_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and95_i_stall_local;
wire [31:0] local_bb4_and95_i;

assign local_bb4_and95_i = ((rnode_232to233_bb4_align_0_i_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and115_i_stall_local;
wire [31:0] local_bb4_and115_i;

assign local_bb4_and115_i = ((rnode_232to233_bb4_align_0_i_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and130_i_stall_local;
wire [31:0] local_bb4_and130_i;

assign local_bb4_and130_i = ((rnode_232to233_bb4_align_0_i_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and149_i_stall_local;
wire [31:0] local_bb4_and149_i;

assign local_bb4_and149_i = ((rnode_232to233_bb4_align_0_i_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4__32_i210_stall_local;
wire [31:0] local_bb4__32_i210;

assign local_bb4__32_i210 = (local_bb4__31_i209 ? (local_bb4_shl1_i_i & 32'hFFFFFE00) : (local_bb4_shl1_i18_i & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__34_i_stall_local;
wire [31:0] local_bb4__34_i;

assign local_bb4__34_i = (local_bb4__31_i209 ? (local_bb4_or_i_i208 & 32'h1FFFFFF) : (local_bb4_or_i17_i & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__36_i_stall_local;
wire [31:0] local_bb4__36_i;

assign local_bb4__36_i = (local_bb4__31_i209 ? (rnode_231to233_bb4_add_i206_2_NO_SHIFT_REG & 32'h1FF) : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i_stall_local;
wire local_bb4_lnot33_not_i;

assign local_bb4_lnot33_not_i = ((local_bb4_and21_i & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or64_i_stall_local;
wire [31:0] local_bb4_or64_i;

assign local_bb4_or64_i = ((local_bb4_and21_i & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and20_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and20_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and20_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and20_i_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and20_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and20_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and20_i_0_valid_out_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and20_i_0_stall_in_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and20_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_and20_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_and20_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_and20_i_0_stall_in_0_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_and20_i_0_valid_out_0_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_and20_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i & 32'h7FFFFF)),
	.data_out(rnode_233to234_bb4_and20_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_and20_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_and20_i_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_233to234_bb4_and20_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_and20_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_and20_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i_stall_in = 1'b0;
assign rnode_233to234_bb4_and20_i_0_stall_in_0_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4_and20_i_0_NO_SHIFT_REG = rnode_233to234_bb4_and20_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4_and20_i_1_NO_SHIFT_REG = rnode_233to234_bb4_and20_i_0_reg_234_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and35_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and35_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and35_i_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and35_i_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and35_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_and35_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_and35_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_and35_i_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_and35_i_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_and35_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i & 32'h80000000)),
	.data_out(rnode_233to234_bb4_and35_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_and35_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_and35_i_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_233to234_bb4_and35_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_and35_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_and35_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i_stall_in = 1'b0;
assign rnode_233to234_bb4_and35_i_0_NO_SHIFT_REG = rnode_233to234_bb4_and35_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_and35_i_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp37_i_stall_local;
wire local_bb4_cmp37_i;

assign local_bb4_cmp37_i = ($signed(local_bb4_xor_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor_lobit_i_stall_local;
wire [31:0] local_bb4_xor_lobit_i;

assign local_bb4_xor_lobit_i = ($signed(local_bb4_xor_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and36_lobit_i_stall_local;
wire [31:0] local_bb4_and36_lobit_i;

assign local_bb4_and36_lobit_i = (local_bb4_xor_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i_stall_local;
wire local_bb4_lnot_i;

assign local_bb4_lnot_i = ((local_bb4_and17_i & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i5_stall_local;
wire local_bb4_cmp25_i5;

assign local_bb4_cmp25_i5 = ((local_bb4_and17_i & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp96_i_stall_local;
wire local_bb4_cmp96_i;

assign local_bb4_cmp96_i = ((local_bb4_and95_i & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp116_i_stall_local;
wire local_bb4_cmp116_i;

assign local_bb4_cmp116_i = ((local_bb4_and115_i & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp131_not_i_stall_local;
wire local_bb4_cmp131_not_i;

assign local_bb4_cmp131_not_i = ((local_bb4_and130_i & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i_stall_local;
wire local_bb4_Pivot20_i;

assign local_bb4_Pivot20_i = ((local_bb4_and149_i & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i_stall_local;
wire local_bb4_SwitchLeaf_i;

assign local_bb4_SwitchLeaf_i = ((local_bb4_and149_i & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i211_stall_local;
wire [31:0] local_bb4__33_i211;

assign local_bb4__33_i211 = (local_bb4_tobool49_i ? (local_bb4__32_i210 & 32'hFFFFFF00) : (local_bb4_shl1_i18_i & 32'hFFFFFF00));

// This section implements an unregistered operation.
// 
wire local_bb4__35_i_stall_local;
wire [31:0] local_bb4__35_i;

assign local_bb4__35_i = (local_bb4_tobool49_i ? (local_bb4__34_i & 32'h1FFFFFF) : (local_bb4_or_i17_i & 32'hFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__37_i_stall_local;
wire [31:0] local_bb4__37_i;

assign local_bb4__37_i = (local_bb4_tobool49_i ? (local_bb4__36_i & 32'h1FF) : (local_bb4_inc_i & 32'h3FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl65_i_stall_local;
wire [31:0] local_bb4_shl65_i;

assign local_bb4_shl65_i = ((local_bb4_or64_i & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i_stall_local;
wire local_bb4_lnot30_i;

assign local_bb4_lnot30_i = ((rnode_233to234_bb4_and20_i_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i6_stall_local;
wire [31:0] local_bb4_or_i6;

assign local_bb4_or_i6 = ((rnode_233to234_bb4_and20_i_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_234to236_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_234to236_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and35_i_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_234to236_bb4_and35_i_0_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and35_i_0_valid_out_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and35_i_0_stall_in_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and35_i_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_234to236_bb4_and35_i_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to236_bb4_and35_i_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to236_bb4_and35_i_0_stall_in_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_234to236_bb4_and35_i_0_valid_out_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_234to236_bb4_and35_i_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in((rnode_233to234_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_234to236_bb4_and35_i_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_234to236_bb4_and35_i_0_reg_236_fifo.DEPTH = 2;
defparam rnode_234to236_bb4_and35_i_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_234to236_bb4_and35_i_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to236_bb4_and35_i_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_234to236_bb4_and35_i_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_and35_i_0_NO_SHIFT_REG = rnode_234to236_bb4_and35_i_0_reg_236_NO_SHIFT_REG;
assign rnode_234to236_bb4_and35_i_0_stall_in_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i_stall_local;
wire local_bb4_cmp25_not_i;

assign local_bb4_cmp25_not_i = (local_bb4_cmp25_i5 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u73_stall_local;
wire local_bb4_var__u73;

assign local_bb4_var__u73 = (local_bb4_cmp25_i5 | rnode_232to234_bb4_cmp27_i_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i214_stall_local;
wire [31:0] local_bb4_and75_i214;

assign local_bb4_and75_i214 = ((local_bb4__35_i & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__33_i211_valid_out;
wire local_bb4__33_i211_stall_in;
wire local_bb4__37_i_valid_out;
wire local_bb4__37_i_stall_in;
wire local_bb4_and75_i214_valid_out;
wire local_bb4_and75_i214_stall_in;
wire local_bb4_and83_i_valid_out;
wire local_bb4_and83_i_stall_in;
wire local_bb4_and83_i_inputs_ready;
wire local_bb4_and83_i_stall_local;
wire [31:0] local_bb4_and83_i;

assign local_bb4_and83_i_inputs_ready = (local_bb4_mul_i_i_valid_out_0_NO_SHIFT_REG & rnode_231to233_bb4_add_i206_0_valid_out_1_NO_SHIFT_REG & rnode_231to233_bb4_add_i206_0_valid_out_0_NO_SHIFT_REG & rnode_231to233_bb4_add_i206_0_valid_out_2_NO_SHIFT_REG & local_bb4_mul_i_i_valid_out_1_NO_SHIFT_REG);
assign local_bb4_and83_i = ((local_bb4__35_i & 32'h1FFFFFF) & 32'h1);
assign local_bb4__33_i211_valid_out = 1'b1;
assign local_bb4__37_i_valid_out = 1'b1;
assign local_bb4_and75_i214_valid_out = 1'b1;
assign local_bb4_and83_i_valid_out = 1'b1;
assign local_bb4_mul_i_i_stall_in_0 = 1'b0;
assign rnode_231to233_bb4_add_i206_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_231to233_bb4_add_i206_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_231to233_bb4_add_i206_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign local_bb4_mul_i_i_stall_in_1 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__28_i_stall_local;
wire [31:0] local_bb4__28_i;

assign local_bb4__28_i = (rnode_232to233_bb4_lnot23_i_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl65_i & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i_stall_local;
wire local_bb4_lnot30_not_i;

assign local_bb4_lnot30_not_i = (local_bb4_lnot30_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i7_stall_local;
wire [31:0] local_bb4_shl_i7;

assign local_bb4_shl_i7 = ((local_bb4_or_i6 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_and35_i_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and35_i_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_and35_i_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and35_i_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and35_i_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and35_i_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_and35_i_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_and35_i_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_and35_i_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_and35_i_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_and35_i_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in((rnode_234to236_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_236to237_bb4_and35_i_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_and35_i_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_and35_i_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_236to237_bb4_and35_i_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_and35_i_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_and35_i_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_234to236_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_and35_i_0_NO_SHIFT_REG = rnode_236to237_bb4_and35_i_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_and35_i_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i_stall_local;
wire local_bb4_or_cond_i;

assign local_bb4_or_cond_i = (local_bb4_lnot30_i | local_bb4_cmp25_not_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4__33_i211_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4__33_i211_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__33_i211_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4__33_i211_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4__33_i211_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__33_i211_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4__33_i211_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__33_i211_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4__33_i211_0_valid_out_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4__33_i211_0_stall_in_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4__33_i211_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4__33_i211_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4__33_i211_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4__33_i211_0_stall_in_0_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4__33_i211_0_valid_out_0_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4__33_i211_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in((local_bb4__33_i211 & 32'hFFFFFF00)),
	.data_out(rnode_233to234_bb4__33_i211_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4__33_i211_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4__33_i211_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_233to234_bb4__33_i211_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4__33_i211_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4__33_i211_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__33_i211_stall_in = 1'b0;
assign rnode_233to234_bb4__33_i211_0_stall_in_0_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4__33_i211_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4__33_i211_0_NO_SHIFT_REG = rnode_233to234_bb4__33_i211_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4__33_i211_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4__33_i211_1_NO_SHIFT_REG = rnode_233to234_bb4__33_i211_0_reg_234_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4__37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__37_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__37_i_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__37_i_2_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__37_i_3_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4__37_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_valid_out_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_stall_in_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4__37_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4__37_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4__37_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4__37_i_0_stall_in_0_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4__37_i_0_valid_out_0_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4__37_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in((local_bb4__37_i & 32'h3FF)),
	.data_out(rnode_233to234_bb4__37_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4__37_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4__37_i_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_233to234_bb4__37_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4__37_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4__37_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__37_i_stall_in = 1'b0;
assign rnode_233to234_bb4__37_i_0_stall_in_0_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4__37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4__37_i_0_NO_SHIFT_REG = rnode_233to234_bb4__37_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4__37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4__37_i_1_NO_SHIFT_REG = rnode_233to234_bb4__37_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4__37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4__37_i_2_NO_SHIFT_REG = rnode_233to234_bb4__37_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4__37_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4__37_i_3_NO_SHIFT_REG = rnode_233to234_bb4__37_i_0_reg_234_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_233to235_bb4_and75_i214_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to235_bb4_and75_i214_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_233to235_bb4_and75_i214_0_NO_SHIFT_REG;
 logic rnode_233to235_bb4_and75_i214_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to235_bb4_and75_i214_0_reg_235_NO_SHIFT_REG;
 logic rnode_233to235_bb4_and75_i214_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_233to235_bb4_and75_i214_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_233to235_bb4_and75_i214_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_233to235_bb4_and75_i214_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to235_bb4_and75_i214_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to235_bb4_and75_i214_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_233to235_bb4_and75_i214_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_233to235_bb4_and75_i214_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in((local_bb4_and75_i214 & 32'h7FFFFF)),
	.data_out(rnode_233to235_bb4_and75_i214_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_233to235_bb4_and75_i214_0_reg_235_fifo.DEPTH = 2;
defparam rnode_233to235_bb4_and75_i214_0_reg_235_fifo.DATA_WIDTH = 32;
defparam rnode_233to235_bb4_and75_i214_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to235_bb4_and75_i214_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_233to235_bb4_and75_i214_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and75_i214_stall_in = 1'b0;
assign rnode_233to235_bb4_and75_i214_0_NO_SHIFT_REG = rnode_233to235_bb4_and75_i214_0_reg_235_NO_SHIFT_REG;
assign rnode_233to235_bb4_and75_i214_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_233to235_bb4_and75_i214_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_and83_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and83_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and83_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and83_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and83_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and83_i_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and83_i_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and83_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_and83_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_and83_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_and83_i_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_and83_i_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_and83_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in((local_bb4_and83_i & 32'h1)),
	.data_out(rnode_233to234_bb4_and83_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_and83_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_and83_i_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_233to234_bb4_and83_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_and83_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_and83_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and83_i_stall_in = 1'b0;
assign rnode_233to234_bb4_and83_i_0_NO_SHIFT_REG = rnode_233to234_bb4_and83_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_and83_i_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and83_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and72_i_stall_local;
wire [31:0] local_bb4_and72_i;

assign local_bb4_and72_i = ((local_bb4__28_i & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i_stall_local;
wire [31:0] local_bb4_and75_i;

assign local_bb4_and75_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and78_i_stall_local;
wire [31:0] local_bb4_and78_i;

assign local_bb4_and78_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr94_i_stall_local;
wire [31:0] local_bb4_shr94_i;

assign local_bb4_shr94_i = ((local_bb4__28_i & 32'h7FFFFF8) >> (local_bb4_and93_i & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i_stall_local;
wire [31:0] local_bb4_and90_i;

assign local_bb4_and90_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and87_i_stall_local;
wire [31:0] local_bb4_and87_i;

assign local_bb4_and87_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and84_i_stall_local;
wire [31:0] local_bb4_and84_i;

assign local_bb4_and84_i = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u74_stall_local;
wire [31:0] local_bb4_var__u74;

assign local_bb4_var__u74 = ((local_bb4__28_i & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i_stall_local;
wire local_bb4_or_cond_not_i;

assign local_bb4_or_cond_not_i = (local_bb4_cmp25_i5 & local_bb4_lnot30_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i_stall_local;
wire [31:0] local_bb4__27_i;

assign local_bb4__27_i = (local_bb4_lnot_i ? 32'h0 : ((local_bb4_shl_i7 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i_stall_local;
wire local_bb4_reduction_8_i;

assign local_bb4_reduction_8_i = (rnode_232to234_bb4_cmp27_i_1_NO_SHIFT_REG & local_bb4_or_cond_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp77_i_stall_local;
wire local_bb4_cmp77_i;

assign local_bb4_cmp77_i = ((rnode_233to234_bb4__33_i211_0_NO_SHIFT_REG & 32'hFFFFFF00) > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u75_stall_local;
wire local_bb4_var__u75;

assign local_bb4_var__u75 = ($signed((rnode_233to234_bb4__33_i211_1_NO_SHIFT_REG & 32'hFFFFFF00)) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp53_i_stall_local;
wire local_bb4_cmp53_i;

assign local_bb4_cmp53_i = ((rnode_233to234_bb4__37_i_0_NO_SHIFT_REG & 32'h3FF) > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp68_i_valid_out;
wire local_bb4_cmp68_i_stall_in;
wire local_bb4_cmp68_i_inputs_ready;
wire local_bb4_cmp68_i_stall_local;
wire local_bb4_cmp68_i;

assign local_bb4_cmp68_i_inputs_ready = rnode_233to234_bb4__37_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp68_i = ((rnode_233to234_bb4__37_i_1_NO_SHIFT_REG & 32'h3FF) < 32'h80);
assign local_bb4_cmp68_i_valid_out = 1'b1;
assign rnode_233to234_bb4__37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i215_stall_local;
wire [31:0] local_bb4_sub_i215;

assign local_bb4_sub_i215 = ((rnode_233to234_bb4__37_i_2_NO_SHIFT_REG & 32'h3FF) << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp71_not_i_valid_out;
wire local_bb4_cmp71_not_i_stall_in;
wire local_bb4_cmp71_not_i_inputs_ready;
wire local_bb4_cmp71_not_i_stall_local;
wire local_bb4_cmp71_not_i;

assign local_bb4_cmp71_not_i_inputs_ready = rnode_233to234_bb4__37_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4_cmp71_not_i = ((rnode_233to234_bb4__37_i_3_NO_SHIFT_REG & 32'h3FF) != 32'h7F);
assign local_bb4_cmp71_not_i_valid_out = 1'b1;
assign rnode_233to234_bb4__37_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool84_i_stall_local;
wire local_bb4_tobool84_i;

assign local_bb4_tobool84_i = ((rnode_233to234_bb4_and83_i_0_NO_SHIFT_REG & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and72_tr_i_stall_local;
wire [7:0] local_bb4_and72_tr_i;
wire [31:0] local_bb4_and72_tr_i$ps;

assign local_bb4_and72_tr_i$ps = (local_bb4_and72_i & 32'hFFFFFF);
assign local_bb4_and72_tr_i = local_bb4_and72_tr_i$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp76_i_stall_local;
wire local_bb4_cmp76_i;

assign local_bb4_cmp76_i = ((local_bb4_and75_i & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp79_i_stall_local;
wire local_bb4_cmp79_i;

assign local_bb4_cmp79_i = ((local_bb4_and78_i & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and142_i_stall_local;
wire [31:0] local_bb4_and142_i;

assign local_bb4_and142_i = (local_bb4_shr94_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr150_i_stall_local;
wire [31:0] local_bb4_shr150_i;

assign local_bb4_shr150_i = (local_bb4_shr94_i >> (local_bb4_and149_i & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u76_stall_local;
wire [31:0] local_bb4_var__u76;

assign local_bb4_var__u76 = (local_bb4_shr94_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and146_i_stall_local;
wire [31:0] local_bb4_and146_i;

assign local_bb4_and146_i = (local_bb4_shr94_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i_stall_local;
wire local_bb4_cmp91_i;

assign local_bb4_cmp91_i = ((local_bb4_and90_i & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp88_i_stall_local;
wire local_bb4_cmp88_i;

assign local_bb4_cmp88_i = ((local_bb4_and87_i & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp85_i_stall_local;
wire local_bb4_cmp85_i;

assign local_bb4_cmp85_i = ((local_bb4_and84_i & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u77_stall_local;
wire local_bb4_var__u77;

assign local_bb4_var__u77 = ((local_bb4_var__u74 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or581_i_valid_out;
wire local_bb4_or581_i_stall_in;
wire local_bb4_or581_i_inputs_ready;
wire local_bb4_or581_i_stall_local;
wire local_bb4_or581_i;

assign local_bb4_or581_i_inputs_ready = (rnode_233to234_bb4_var__u71_0_valid_out_NO_SHIFT_REG & rnode_233to234_bb4__37_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4_or581_i = (rnode_233to234_bb4_var__u71_0_NO_SHIFT_REG | local_bb4_cmp53_i);
assign local_bb4_or581_i_valid_out = 1'b1;
assign rnode_233to234_bb4_var__u71_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4__37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_cmp68_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp68_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp68_i_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp68_i_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp68_i_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp68_i_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp68_i_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp68_i_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_cmp68_i_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_cmp68_i_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_cmp68_i_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_cmp68_i_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_cmp68_i_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(local_bb4_cmp68_i),
	.data_out(rnode_234to235_bb4_cmp68_i_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_cmp68_i_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_cmp68_i_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4_cmp68_i_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_cmp68_i_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_cmp68_i_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp68_i_stall_in = 1'b0;
assign rnode_234to235_bb4_cmp68_i_0_NO_SHIFT_REG = rnode_234to235_bb4_cmp68_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_cmp68_i_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_cmp68_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and74_i_stall_local;
wire [31:0] local_bb4_and74_i;

assign local_bb4_and74_i = ((local_bb4_sub_i215 & 32'hFF800000) + 32'h40800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_cmp71_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp71_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp71_not_i_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp71_not_i_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp71_not_i_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp71_not_i_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp71_not_i_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_cmp71_not_i_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_cmp71_not_i_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_cmp71_not_i_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_cmp71_not_i_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_cmp71_not_i_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_cmp71_not_i_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(local_bb4_cmp71_not_i),
	.data_out(rnode_234to235_bb4_cmp71_not_i_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_cmp71_not_i_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_cmp71_not_i_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4_cmp71_not_i_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_cmp71_not_i_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_cmp71_not_i_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp71_not_i_stall_in = 1'b0;
assign rnode_234to235_bb4_cmp71_not_i_0_NO_SHIFT_REG = rnode_234to235_bb4_cmp71_not_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_cmp71_not_i_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_cmp71_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__39_i_stall_local;
wire local_bb4__39_i;

assign local_bb4__39_i = (local_bb4_tobool84_i & local_bb4_var__u75);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool74_i_stall_local;
wire [7:0] local_bb4_frombool74_i;

assign local_bb4_frombool74_i = (local_bb4_and72_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u78_stall_local;
wire [31:0] local_bb4_var__u78;

assign local_bb4_var__u78 = ((local_bb4_and146_i & 32'h3FFFFFFF) | local_bb4_shr94_i);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i_stall_local;
wire local_bb4__31_v_i;

assign local_bb4__31_v_i = (local_bb4_cmp96_i ? local_bb4_cmp79_i : local_bb4_cmp91_i);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i_stall_local;
wire local_bb4__30_v_i;

assign local_bb4__30_v_i = (local_bb4_cmp96_i ? local_bb4_cmp76_i : local_bb4_cmp88_i);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool109_i_stall_local;
wire [7:0] local_bb4_frombool109_i;

assign local_bb4_frombool109_i[7:1] = 7'h0;
assign local_bb4_frombool109_i[0] = local_bb4_cmp85_i;

// This section implements an unregistered operation.
// 
wire local_bb4_or107_i_stall_local;
wire [31:0] local_bb4_or107_i;

assign local_bb4_or107_i[31:1] = 31'h0;
assign local_bb4_or107_i[0] = local_bb4_var__u77;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_or581_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_1_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_valid_out_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_stall_in_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_or581_i_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_or581_i_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_or581_i_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_or581_i_0_stall_in_0_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_or581_i_0_valid_out_0_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_or581_i_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(local_bb4_or581_i),
	.data_out(rnode_234to235_bb4_or581_i_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_or581_i_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_or581_i_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4_or581_i_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_or581_i_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_or581_i_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or581_i_stall_in = 1'b0;
assign rnode_234to235_bb4_or581_i_0_stall_in_0_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_or581_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4_or581_i_0_NO_SHIFT_REG = rnode_234to235_bb4_or581_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_or581_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4_or581_i_1_NO_SHIFT_REG = rnode_234to235_bb4_or581_i_0_reg_235_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u79_stall_local;
wire [31:0] local_bb4_var__u79;

assign local_bb4_var__u79[31:1] = 31'h0;
assign local_bb4_var__u79[0] = rnode_234to235_bb4_cmp68_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i216_valid_out;
wire local_bb4_shl_i216_stall_in;
wire local_bb4_shl_i216_inputs_ready;
wire local_bb4_shl_i216_stall_local;
wire [31:0] local_bb4_shl_i216;

assign local_bb4_shl_i216_inputs_ready = rnode_233to234_bb4__37_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shl_i216 = ((local_bb4_and74_i & 32'hFF800000) & 32'h7F800000);
assign local_bb4_shl_i216_valid_out = 1'b1;
assign rnode_233to234_bb4__37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__40_i_valid_out;
wire local_bb4__40_i_stall_in;
wire local_bb4__40_i_inputs_ready;
wire local_bb4__40_i_stall_local;
wire local_bb4__40_i;

assign local_bb4__40_i_inputs_ready = (rnode_233to234_bb4__33_i211_0_valid_out_0_NO_SHIFT_REG & rnode_233to234_bb4__33_i211_0_valid_out_1_NO_SHIFT_REG & rnode_233to234_bb4_and83_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4__40_i = (local_bb4_cmp77_i | local_bb4__39_i);
assign local_bb4__40_i_valid_out = 1'b1;
assign rnode_233to234_bb4__33_i211_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4__33_i211_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and83_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or1596_i_stall_local;
wire [31:0] local_bb4_or1596_i;

assign local_bb4_or1596_i = (local_bb4_var__u78 | (local_bb4_and142_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i_stall_local;
wire [7:0] local_bb4__31_i;

assign local_bb4__31_i[7:1] = 7'h0;
assign local_bb4__31_i[0] = local_bb4__31_v_i;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i_stall_local;
wire [7:0] local_bb4__30_i;

assign local_bb4__30_i[7:1] = 7'h0;
assign local_bb4__30_i[0] = local_bb4__30_v_i;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i_stall_local;
wire [7:0] local_bb4__29_i;

assign local_bb4__29_i = (local_bb4_cmp96_i ? (local_bb4_frombool74_i & 8'h1) : (local_bb4_frombool109_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i_stall_local;
wire [31:0] local_bb4__32_i;

assign local_bb4__32_i = (local_bb4_cmp96_i ? 32'h0 : (local_bb4_or107_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i213_stall_local;
wire local_bb4_reduction_2_i213;

assign local_bb4_reduction_2_i213 = (rnode_234to235_bb4_reduction_0_i212_0_NO_SHIFT_REG | rnode_234to235_bb4_or581_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_cond111_i_stall_local;
wire [31:0] local_bb4_cond111_i;

assign local_bb4_cond111_i = (rnode_234to235_bb4_or581_i_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_shl_i216_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_shl_i216_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_shl_i216_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_shl_i216_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_shl_i216_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_shl_i216_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_shl_i216_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_shl_i216_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_shl_i216_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_shl_i216_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_shl_i216_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_shl_i216_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_shl_i216_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in((local_bb4_shl_i216 & 32'h7F800000)),
	.data_out(rnode_234to235_bb4_shl_i216_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_shl_i216_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_shl_i216_0_reg_235_fifo.DATA_WIDTH = 32;
defparam rnode_234to235_bb4_shl_i216_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_shl_i216_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_shl_i216_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shl_i216_stall_in = 1'b0;
assign rnode_234to235_bb4_shl_i216_0_NO_SHIFT_REG = rnode_234to235_bb4_shl_i216_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_shl_i216_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_shl_i216_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4__40_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4__40_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4__40_i_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4__40_i_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4__40_i_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__40_i_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__40_i_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__40_i_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4__40_i_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4__40_i_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4__40_i_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4__40_i_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4__40_i_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(local_bb4__40_i),
	.data_out(rnode_234to235_bb4__40_i_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4__40_i_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4__40_i_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4__40_i_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4__40_i_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4__40_i_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__40_i_stall_in = 1'b0;
assign rnode_234to235_bb4__40_i_0_NO_SHIFT_REG = rnode_234to235_bb4__40_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4__40_i_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4__40_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or162_i_stall_local;
wire [31:0] local_bb4_or162_i;

assign local_bb4_or162_i = (local_bb4_or1596_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1237_i_stall_local;
wire [7:0] local_bb4_or1237_i;

assign local_bb4_or1237_i = ((local_bb4__30_i & 8'h1) | (local_bb4__29_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i_stall_local;
wire [7:0] local_bb4__33_i;

assign local_bb4__33_i = (local_bb4_cmp116_i ? (local_bb4__29_i & 8'h1) : (local_bb4__31_i & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv101_i_stall_local;
wire [31:0] local_bb4_conv101_i;

assign local_bb4_conv101_i[31:1] = 31'h0;
assign local_bb4_conv101_i[0] = local_bb4_reduction_2_i213;

// This section implements an unregistered operation.
// 
wire local_bb4_or76_i_stall_local;
wire [31:0] local_bb4_or76_i;

assign local_bb4_or76_i = ((rnode_234to235_bb4_shl_i216_0_NO_SHIFT_REG & 32'h7F800000) | (rnode_233to235_bb4_and75_i214_0_NO_SHIFT_REG & 32'h7FFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond_i217_stall_local;
wire [31:0] local_bb4_cond_i217;

assign local_bb4_cond_i217[31:1] = 31'h0;
assign local_bb4_cond_i217[0] = rnode_234to235_bb4__40_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i_stall_local;
wire [31:0] local_bb4__37_v_i;

assign local_bb4__37_v_i = (local_bb4_Pivot20_i ? 32'h0 : (local_bb4_or162_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or123_i_stall_local;
wire [31:0] local_bb4_or123_i;

assign local_bb4_or123_i[31:8] = 24'h0;
assign local_bb4_or123_i[7:0] = (local_bb4_or1237_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u80_stall_local;
wire [7:0] local_bb4_var__u80;

assign local_bb4_var__u80 = ((local_bb4__33_i & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_add87_i_stall_local;
wire [31:0] local_bb4_add87_i;

assign local_bb4_add87_i = ((local_bb4_cond_i217 & 32'h1) + (local_bb4_or76_i & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i_stall_local;
wire [31:0] local_bb4__39_v_i;

assign local_bb4__39_v_i = (local_bb4_SwitchLeaf_i ? (local_bb4_var__u76 & 32'h1) : (local_bb4__37_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i_stall_local;
wire [31:0] local_bb4_or124_i;

assign local_bb4_or124_i = (local_bb4_cmp116_i ? 32'h0 : (local_bb4_or123_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv135_i_stall_local;
wire [31:0] local_bb4_conv135_i;

assign local_bb4_conv135_i[31:8] = 24'h0;
assign local_bb4_conv135_i[7:0] = (local_bb4_var__u80 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and88_i_stall_local;
wire [31:0] local_bb4_and88_i;

assign local_bb4_and88_i = (local_bb4_add87_i & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i218_stall_local;
wire [31:0] local_bb4_and90_i218;

assign local_bb4_and90_i218 = (local_bb4_add87_i & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i_stall_local;
wire [31:0] local_bb4_reduction_3_i;

assign local_bb4_reduction_3_i = ((local_bb4__32_i & 32'h1) | (local_bb4_or124_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or136_i_stall_local;
wire [31:0] local_bb4_or136_i;

assign local_bb4_or136_i = (local_bb4_cmp131_not_i ? (local_bb4_conv135_i & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or89_i_stall_local;
wire [31:0] local_bb4_or89_i;

assign local_bb4_or89_i = ((local_bb4_and88_i & 32'h7FFFFFFF) | (local_bb4_and4_i & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i219_stall_local;
wire local_bb4_cmp91_i219;

assign local_bb4_cmp91_i219 = ((local_bb4_and90_i218 & 32'h800000) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i_stall_local;
wire [31:0] local_bb4_reduction_5_i;

assign local_bb4_reduction_5_i = (local_bb4_shr150_i | (local_bb4_reduction_3_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i_stall_local;
wire [31:0] local_bb4_reduction_4_i;

assign local_bb4_reduction_4_i = ((local_bb4_or136_i & 32'h1) | (local_bb4__39_v_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge14_i_stall_local;
wire local_bb4_brmerge14_i;

assign local_bb4_brmerge14_i = (local_bb4_cmp91_i219 | rnode_234to235_bb4_cmp71_not_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i_stall_local;
wire [31:0] local_bb4_reduction_6_i;

assign local_bb4_reduction_6_i = ((local_bb4_reduction_4_i & 32'h1) | local_bb4_reduction_5_i);

// This section implements an unregistered operation.
// 
wire local_bb4_conv99_i_stall_local;
wire [31:0] local_bb4_conv99_i;

assign local_bb4_conv99_i = (local_bb4_brmerge14_i ? (local_bb4_var__u79 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i_valid_out;
wire local_bb4_lnot33_not_i_stall_in;
wire local_bb4_cmp37_i_valid_out;
wire local_bb4_cmp37_i_stall_in;
wire local_bb4_and36_lobit_i_valid_out;
wire local_bb4_and36_lobit_i_stall_in;
wire local_bb4_xor188_i_valid_out;
wire local_bb4_xor188_i_stall_in;
wire local_bb4_xor188_i_inputs_ready;
wire local_bb4_xor188_i_stall_local;
wire [31:0] local_bb4_xor188_i;

assign local_bb4_xor188_i_inputs_ready = (rnode_232to233_bb4__22_i_0_valid_out_0_NO_SHIFT_REG & rnode_232to233_bb4_lnot23_i_0_valid_out_NO_SHIFT_REG & rnode_232to233_bb4_align_0_i_0_valid_out_0_NO_SHIFT_REG & rnode_232to233_bb4_align_0_i_0_valid_out_4_NO_SHIFT_REG & rnode_232to233_bb4_align_0_i_0_valid_out_1_NO_SHIFT_REG & rnode_232to233_bb4_align_0_i_0_valid_out_2_NO_SHIFT_REG & rnode_232to233_bb4_align_0_i_0_valid_out_3_NO_SHIFT_REG & rnode_232to233_bb4__23_i_0_valid_out_2_NO_SHIFT_REG & rnode_232to233_bb4__22_i_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor188_i = (local_bb4_reduction_6_i ^ local_bb4_xor_lobit_i);
assign local_bb4_lnot33_not_i_valid_out = 1'b1;
assign local_bb4_cmp37_i_valid_out = 1'b1;
assign local_bb4_and36_lobit_i_valid_out = 1'b1;
assign local_bb4_xor188_i_valid_out = 1'b1;
assign rnode_232to233_bb4__22_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_lnot23_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_align_0_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_align_0_i_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_align_0_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_align_0_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4_align_0_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4__23_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_232to233_bb4__22_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or102_i_stall_local;
wire [31:0] local_bb4_or102_i;

assign local_bb4_or102_i = ((local_bb4_conv99_i & 32'h1) | (local_bb4_conv101_i & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to234_bb4_lnot33_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_233to234_bb4_lnot33_not_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_lnot33_not_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_233to234_bb4_lnot33_not_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_lnot33_not_i_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_lnot33_not_i_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_lnot33_not_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_lnot33_not_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_lnot33_not_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_lnot33_not_i_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_lnot33_not_i_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_lnot33_not_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i),
	.data_out(rnode_233to234_bb4_lnot33_not_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_lnot33_not_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_lnot33_not_i_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_233to234_bb4_lnot33_not_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_lnot33_not_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_lnot33_not_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i_stall_in = 1'b0;
assign rnode_233to234_bb4_lnot33_not_i_0_NO_SHIFT_REG = rnode_233to234_bb4_lnot33_not_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_lnot33_not_i_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_valid_out_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_stall_in_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_cmp37_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_cmp37_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_cmp37_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_cmp37_i_0_stall_in_0_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_cmp37_i_0_valid_out_0_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_cmp37_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(local_bb4_cmp37_i),
	.data_out(rnode_233to234_bb4_cmp37_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_cmp37_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_cmp37_i_0_reg_234_fifo.DATA_WIDTH = 1;
defparam rnode_233to234_bb4_cmp37_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_cmp37_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_cmp37_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp37_i_stall_in = 1'b0;
assign rnode_233to234_bb4_cmp37_i_0_stall_in_0_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4_cmp37_i_0_NO_SHIFT_REG = rnode_233to234_bb4_cmp37_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4_cmp37_i_1_NO_SHIFT_REG = rnode_233to234_bb4_cmp37_i_0_reg_234_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and36_lobit_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and36_lobit_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and36_lobit_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_and36_lobit_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and36_lobit_i_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and36_lobit_i_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_and36_lobit_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_and36_lobit_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_and36_lobit_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_and36_lobit_i_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_and36_lobit_i_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_and36_lobit_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in((local_bb4_and36_lobit_i & 32'h1)),
	.data_out(rnode_233to234_bb4_and36_lobit_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_and36_lobit_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_and36_lobit_i_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_233to234_bb4_and36_lobit_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_and36_lobit_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_and36_lobit_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and36_lobit_i_stall_in = 1'b0;
assign rnode_233to234_bb4_and36_lobit_i_0_NO_SHIFT_REG = rnode_233to234_bb4_and36_lobit_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_and36_lobit_i_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_233to234_bb4_xor188_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_233to234_bb4_xor188_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_xor188_i_0_NO_SHIFT_REG;
 logic rnode_233to234_bb4_xor188_i_0_reg_234_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_233to234_bb4_xor188_i_0_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_xor188_i_0_valid_out_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_xor188_i_0_stall_in_reg_234_NO_SHIFT_REG;
 logic rnode_233to234_bb4_xor188_i_0_stall_out_reg_234_NO_SHIFT_REG;

acl_data_fifo rnode_233to234_bb4_xor188_i_0_reg_234_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_233to234_bb4_xor188_i_0_reg_234_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_233to234_bb4_xor188_i_0_stall_in_reg_234_NO_SHIFT_REG),
	.valid_out(rnode_233to234_bb4_xor188_i_0_valid_out_reg_234_NO_SHIFT_REG),
	.stall_out(rnode_233to234_bb4_xor188_i_0_stall_out_reg_234_NO_SHIFT_REG),
	.data_in(local_bb4_xor188_i),
	.data_out(rnode_233to234_bb4_xor188_i_0_reg_234_NO_SHIFT_REG)
);

defparam rnode_233to234_bb4_xor188_i_0_reg_234_fifo.DEPTH = 1;
defparam rnode_233to234_bb4_xor188_i_0_reg_234_fifo.DATA_WIDTH = 32;
defparam rnode_233to234_bb4_xor188_i_0_reg_234_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_233to234_bb4_xor188_i_0_reg_234_fifo.IMPL = "shift_reg";

assign rnode_233to234_bb4_xor188_i_0_reg_234_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor188_i_stall_in = 1'b0;
assign rnode_233to234_bb4_xor188_i_0_NO_SHIFT_REG = rnode_233to234_bb4_xor188_i_0_reg_234_NO_SHIFT_REG;
assign rnode_233to234_bb4_xor188_i_0_stall_in_reg_234_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_xor188_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_tobool103_i_stall_local;
wire local_bb4_tobool103_i;

assign local_bb4_tobool103_i = ((local_bb4_or102_i & 32'h1) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i_stall_local;
wire local_bb4_brmerge_not_i;

assign local_bb4_brmerge_not_i = (rnode_232to234_bb4_cmp27_i_0_NO_SHIFT_REG & rnode_233to234_bb4_lnot33_not_i_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_234to236_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_2_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_valid_out_0_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_stall_in_0_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_cmp37_i_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_234to236_bb4_cmp37_i_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to236_bb4_cmp37_i_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to236_bb4_cmp37_i_0_stall_in_0_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_234to236_bb4_cmp37_i_0_valid_out_0_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_234to236_bb4_cmp37_i_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in(rnode_233to234_bb4_cmp37_i_1_NO_SHIFT_REG),
	.data_out(rnode_234to236_bb4_cmp37_i_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_234to236_bb4_cmp37_i_0_reg_236_fifo.DEPTH = 2;
defparam rnode_234to236_bb4_cmp37_i_0_reg_236_fifo.DATA_WIDTH = 1;
defparam rnode_234to236_bb4_cmp37_i_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to236_bb4_cmp37_i_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_234to236_bb4_cmp37_i_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_233to234_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_cmp37_i_0_stall_in_0_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_234to236_bb4_cmp37_i_0_NO_SHIFT_REG = rnode_234to236_bb4_cmp37_i_0_reg_236_NO_SHIFT_REG;
assign rnode_234to236_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_234to236_bb4_cmp37_i_1_NO_SHIFT_REG = rnode_234to236_bb4_cmp37_i_0_reg_236_NO_SHIFT_REG;
assign rnode_234to236_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_234to236_bb4_cmp37_i_2_NO_SHIFT_REG = rnode_234to236_bb4_cmp37_i_0_reg_236_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i8_stall_local;
wire [31:0] local_bb4_add_i8;

assign local_bb4_add_i8 = ((local_bb4__27_i & 32'h7FFFFF8) | (rnode_233to234_bb4_and36_lobit_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_cond107_i_stall_local;
wire [31:0] local_bb4_cond107_i;

assign local_bb4_cond107_i = (local_bb4_tobool103_i ? (local_bb4_and4_i & 32'h80000000) : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i_stall_local;
wire local_bb4__24_i;

assign local_bb4__24_i = (local_bb4_or_cond_not_i | local_bb4_brmerge_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i_stall_local;
wire local_bb4_brmerge_not_not_i;

assign local_bb4_brmerge_not_not_i = (local_bb4_brmerge_not_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp37_i_stall_local;
wire local_bb4_not_cmp37_i;

assign local_bb4_not_cmp37_i = (rnode_234to236_bb4_cmp37_i_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add192_i_stall_local;
wire [31:0] local_bb4_add192_i;

assign local_bb4_add192_i = ((local_bb4_add_i8 & 32'h7FFFFF9) + rnode_233to234_bb4_xor188_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and108_i_stall_local;
wire [31:0] local_bb4_and108_i;

assign local_bb4_and108_i = (local_bb4_cond107_i & local_bb4_or89_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i_stall_local;
wire local_bb4_reduction_7_i;

assign local_bb4_reduction_7_i = (local_bb4_cmp25_i5 & local_bb4_brmerge_not_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or112_i_stall_local;
wire [31:0] local_bb4_or112_i;

assign local_bb4_or112_i = (local_bb4_and108_i | (local_bb4_cond111_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i_stall_local;
wire local_bb4_reduction_9_i;

assign local_bb4_reduction_9_i = (local_bb4_reduction_7_i & local_bb4_reduction_8_i);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u81_valid_out;
wire local_bb4_var__u81_stall_in;
wire local_bb4_var__u81_inputs_ready;
wire local_bb4_var__u81_stall_local;
wire [31:0] local_bb4_var__u81;

assign local_bb4_var__u81_inputs_ready = (rnode_234to235_bb4_xor_i195_0_valid_out_NO_SHIFT_REG & rnode_234to235_bb4__29_i204_0_valid_out_NO_SHIFT_REG & rnode_234to235_bb4_or581_i_0_valid_out_1_NO_SHIFT_REG & rnode_234to235_bb4_or581_i_0_valid_out_0_NO_SHIFT_REG & rnode_234to235_bb4_reduction_0_i212_0_valid_out_NO_SHIFT_REG & rnode_234to235_bb4_cmp68_i_0_valid_out_NO_SHIFT_REG & rnode_234to235_bb4_cmp71_not_i_0_valid_out_NO_SHIFT_REG & rnode_234to235_bb4_shl_i216_0_valid_out_NO_SHIFT_REG & rnode_233to235_bb4_and75_i214_0_valid_out_NO_SHIFT_REG & rnode_234to235_bb4__40_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4_var__u81 = (rnode_234to235_bb4__29_i204_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb4_or112_i);
assign local_bb4_var__u81_valid_out = 1'b1;
assign rnode_234to235_bb4_xor_i195_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4__29_i204_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_or581_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_or581_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_reduction_0_i212_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_cmp68_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_cmp71_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_shl_i216_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_233to235_bb4_and75_i214_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4__40_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i_valid_out_2;
wire local_bb4_and17_i_stall_in_2;
wire local_bb4_var__u73_valid_out;
wire local_bb4_var__u73_stall_in;
wire local_bb4_add192_i_valid_out;
wire local_bb4_add192_i_stall_in;
wire local_bb4__26_i_valid_out;
wire local_bb4__26_i_stall_in;
wire local_bb4__26_i_inputs_ready;
wire local_bb4__26_i_stall_local;
wire local_bb4__26_i;

assign local_bb4__26_i_inputs_ready = (rnode_232to234_bb4_shr16_i_0_valid_out_0_NO_SHIFT_REG & rnode_232to234_bb4_cmp27_i_0_valid_out_2_NO_SHIFT_REG & rnode_233to234_bb4_and36_lobit_i_0_valid_out_NO_SHIFT_REG & rnode_233to234_bb4_xor188_i_0_valid_out_NO_SHIFT_REG & rnode_233to234_bb4_and20_i_0_valid_out_0_NO_SHIFT_REG & rnode_232to234_bb4_cmp27_i_0_valid_out_0_NO_SHIFT_REG & rnode_233to234_bb4_lnot33_not_i_0_valid_out_NO_SHIFT_REG & rnode_232to234_bb4_cmp27_i_0_valid_out_1_NO_SHIFT_REG & rnode_233to234_bb4_and20_i_0_valid_out_1_NO_SHIFT_REG & rnode_233to234_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i = (local_bb4_reduction_9_i ? rnode_233to234_bb4_cmp37_i_0_NO_SHIFT_REG : local_bb4__24_i);
assign local_bb4_and17_i_valid_out_2 = 1'b1;
assign local_bb4_var__u73_valid_out = 1'b1;
assign local_bb4_add192_i_valid_out = 1'b1;
assign local_bb4__26_i_valid_out = 1'b1;
assign rnode_232to234_bb4_shr16_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4_cmp27_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and36_lobit_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_xor188_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and20_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4_cmp27_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_lnot33_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_232to234_bb4_cmp27_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_and20_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_233to234_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_235to236_bb4_var__u81_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_var__u81_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_var__u81_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_var__u81_2_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_var__u81_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_valid_out_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_stall_in_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u81_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_235to236_bb4_var__u81_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to236_bb4_var__u81_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to236_bb4_var__u81_0_stall_in_0_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_235to236_bb4_var__u81_0_valid_out_0_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_235to236_bb4_var__u81_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in(local_bb4_var__u81),
	.data_out(rnode_235to236_bb4_var__u81_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_235to236_bb4_var__u81_0_reg_236_fifo.DEPTH = 1;
defparam rnode_235to236_bb4_var__u81_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_235to236_bb4_var__u81_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to236_bb4_var__u81_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_235to236_bb4_var__u81_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u81_stall_in = 1'b0;
assign rnode_235to236_bb4_var__u81_0_stall_in_0_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_var__u81_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_var__u81_0_NO_SHIFT_REG = rnode_235to236_bb4_var__u81_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_var__u81_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_var__u81_1_NO_SHIFT_REG = rnode_235to236_bb4_var__u81_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_var__u81_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_var__u81_2_NO_SHIFT_REG = rnode_235to236_bb4_var__u81_0_reg_236_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_234to236_bb4_and17_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and17_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_234to236_bb4_and17_i_0_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and17_i_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_234to236_bb4_and17_i_0_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and17_i_0_valid_out_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and17_i_0_stall_in_reg_236_NO_SHIFT_REG;
 logic rnode_234to236_bb4_and17_i_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_234to236_bb4_and17_i_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to236_bb4_and17_i_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to236_bb4_and17_i_0_stall_in_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_234to236_bb4_and17_i_0_valid_out_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_234to236_bb4_and17_i_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i & 32'hFF)),
	.data_out(rnode_234to236_bb4_and17_i_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_234to236_bb4_and17_i_0_reg_236_fifo.DEPTH = 2;
defparam rnode_234to236_bb4_and17_i_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_234to236_bb4_and17_i_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to236_bb4_and17_i_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_234to236_bb4_and17_i_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i_stall_in_2 = 1'b0;
assign rnode_234to236_bb4_and17_i_0_NO_SHIFT_REG = rnode_234to236_bb4_and17_i_0_reg_236_NO_SHIFT_REG;
assign rnode_234to236_bb4_and17_i_0_stall_in_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_and17_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_var__u73_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4_var__u73_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4_var__u73_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_var__u73_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4_var__u73_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_var__u73_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_var__u73_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_var__u73_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_var__u73_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_var__u73_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_var__u73_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_var__u73_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_var__u73_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(local_bb4_var__u73),
	.data_out(rnode_234to235_bb4_var__u73_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_var__u73_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_var__u73_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4_var__u73_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_var__u73_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_var__u73_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u73_stall_in = 1'b0;
assign rnode_234to235_bb4_var__u73_0_NO_SHIFT_REG = rnode_234to235_bb4_var__u73_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_var__u73_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_var__u73_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_add192_i_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_add192_i_1_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_add192_i_2_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_add192_i_3_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_234to235_bb4_add192_i_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_valid_out_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_stall_in_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4_add192_i_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4_add192_i_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4_add192_i_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4_add192_i_0_stall_in_0_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4_add192_i_0_valid_out_0_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4_add192_i_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(local_bb4_add192_i),
	.data_out(rnode_234to235_bb4_add192_i_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4_add192_i_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4_add192_i_0_reg_235_fifo.DATA_WIDTH = 32;
defparam rnode_234to235_bb4_add192_i_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4_add192_i_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4_add192_i_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add192_i_stall_in = 1'b0;
assign rnode_234to235_bb4_add192_i_0_stall_in_0_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4_add192_i_0_NO_SHIFT_REG = rnode_234to235_bb4_add192_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4_add192_i_1_NO_SHIFT_REG = rnode_234to235_bb4_add192_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4_add192_i_2_NO_SHIFT_REG = rnode_234to235_bb4_add192_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4_add192_i_3_NO_SHIFT_REG = rnode_234to235_bb4_add192_i_0_reg_235_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_234to235_bb4__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_234to235_bb4__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_234to235_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_234to235_bb4__26_i_0_reg_235_inputs_ready_NO_SHIFT_REG;
 logic rnode_234to235_bb4__26_i_0_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__26_i_0_valid_out_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__26_i_0_stall_in_reg_235_NO_SHIFT_REG;
 logic rnode_234to235_bb4__26_i_0_stall_out_reg_235_NO_SHIFT_REG;

acl_data_fifo rnode_234to235_bb4__26_i_0_reg_235_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_234to235_bb4__26_i_0_reg_235_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_234to235_bb4__26_i_0_stall_in_reg_235_NO_SHIFT_REG),
	.valid_out(rnode_234to235_bb4__26_i_0_valid_out_reg_235_NO_SHIFT_REG),
	.stall_out(rnode_234to235_bb4__26_i_0_stall_out_reg_235_NO_SHIFT_REG),
	.data_in(local_bb4__26_i),
	.data_out(rnode_234to235_bb4__26_i_0_reg_235_NO_SHIFT_REG)
);

defparam rnode_234to235_bb4__26_i_0_reg_235_fifo.DEPTH = 1;
defparam rnode_234to235_bb4__26_i_0_reg_235_fifo.DATA_WIDTH = 1;
defparam rnode_234to235_bb4__26_i_0_reg_235_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_234to235_bb4__26_i_0_reg_235_fifo.IMPL = "shift_reg";

assign rnode_234to235_bb4__26_i_0_reg_235_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i_stall_in = 1'b0;
assign rnode_234to235_bb4__26_i_0_NO_SHIFT_REG = rnode_234to235_bb4__26_i_0_reg_235_NO_SHIFT_REG;
assign rnode_234to235_bb4__26_i_0_stall_in_reg_235_NO_SHIFT_REG = 1'b0;
assign rnode_234to235_bb4__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i11_stall_local;
wire [31:0] local_bb4_and_i11;

assign local_bb4_and_i11 = (rnode_235to236_bb4_var__u81_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and10_i17_stall_local;
wire [31:0] local_bb4_and10_i17;

assign local_bb4_and10_i17 = (rnode_235to236_bb4_var__u81_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_var__u81_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u81_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_var__u81_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u81_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u81_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_var__u81_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u81_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_var__u81_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u81_0_valid_out_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u81_0_stall_in_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u81_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_var__u81_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_var__u81_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_var__u81_0_stall_in_0_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_var__u81_0_valid_out_0_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_var__u81_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(rnode_235to236_bb4_var__u81_2_NO_SHIFT_REG),
	.data_out(rnode_236to237_bb4_var__u81_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_var__u81_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_var__u81_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_236to237_bb4_var__u81_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_var__u81_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_var__u81_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_var__u81_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u81_0_stall_in_0_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u81_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4_var__u81_0_NO_SHIFT_REG = rnode_236to237_bb4_var__u81_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_var__u81_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4_var__u81_1_NO_SHIFT_REG = rnode_236to237_bb4_var__u81_0_reg_237_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_235to236_bb4_var__u73_0_valid_out_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u73_0_stall_in_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u73_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u73_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u73_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u73_0_valid_out_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u73_0_stall_in_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_var__u73_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_235to236_bb4_var__u73_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to236_bb4_var__u73_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to236_bb4_var__u73_0_stall_in_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_235to236_bb4_var__u73_0_valid_out_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_235to236_bb4_var__u73_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in(rnode_234to235_bb4_var__u73_0_NO_SHIFT_REG),
	.data_out(rnode_235to236_bb4_var__u73_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_235to236_bb4_var__u73_0_reg_236_fifo.DEPTH = 1;
defparam rnode_235to236_bb4_var__u73_0_reg_236_fifo.DATA_WIDTH = 1;
defparam rnode_235to236_bb4_var__u73_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to236_bb4_var__u73_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_235to236_bb4_var__u73_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4_var__u73_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_var__u73_0_NO_SHIFT_REG = rnode_235to236_bb4_var__u73_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_var__u73_0_stall_in_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_var__u73_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and193_i_valid_out;
wire local_bb4_and193_i_stall_in;
wire local_bb4_and193_i_inputs_ready;
wire local_bb4_and193_i_stall_local;
wire [31:0] local_bb4_and193_i;

assign local_bb4_and193_i_inputs_ready = rnode_234to235_bb4_add192_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and193_i = (rnode_234to235_bb4_add192_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and193_i_valid_out = 1'b1;
assign rnode_234to235_bb4_add192_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and195_i_valid_out;
wire local_bb4_and195_i_stall_in;
wire local_bb4_and195_i_inputs_ready;
wire local_bb4_and195_i_stall_local;
wire [31:0] local_bb4_and195_i;

assign local_bb4_and195_i_inputs_ready = rnode_234to235_bb4_add192_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and195_i = (rnode_234to235_bb4_add192_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and195_i_valid_out = 1'b1;
assign rnode_234to235_bb4_add192_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and198_i_valid_out;
wire local_bb4_and198_i_stall_in;
wire local_bb4_and198_i_inputs_ready;
wire local_bb4_and198_i_stall_local;
wire [31:0] local_bb4_and198_i;

assign local_bb4_and198_i_inputs_ready = rnode_234to235_bb4_add192_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and198_i = (rnode_234to235_bb4_add192_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and198_i_valid_out = 1'b1;
assign rnode_234to235_bb4_add192_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and201_i_stall_local;
wire [31:0] local_bb4_and201_i;

assign local_bb4_and201_i = (rnode_234to235_bb4_add192_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_235to237_bb4__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_235to237_bb4__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_235to237_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_235to237_bb4__26_i_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic rnode_235to237_bb4__26_i_0_reg_237_NO_SHIFT_REG;
 logic rnode_235to237_bb4__26_i_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_235to237_bb4__26_i_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_235to237_bb4__26_i_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_235to237_bb4__26_i_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to237_bb4__26_i_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to237_bb4__26_i_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_235to237_bb4__26_i_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_235to237_bb4__26_i_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(rnode_234to235_bb4__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_235to237_bb4__26_i_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_235to237_bb4__26_i_0_reg_237_fifo.DEPTH = 2;
defparam rnode_235to237_bb4__26_i_0_reg_237_fifo.DATA_WIDTH = 1;
defparam rnode_235to237_bb4__26_i_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to237_bb4__26_i_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_235to237_bb4__26_i_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_234to235_bb4__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_235to237_bb4__26_i_0_NO_SHIFT_REG = rnode_235to237_bb4__26_i_0_reg_237_NO_SHIFT_REG;
assign rnode_235to237_bb4__26_i_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_235to237_bb4__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i12_stall_local;
wire [31:0] local_bb4_shr_i12;

assign local_bb4_shr_i12 = ((local_bb4_and_i11 & 32'hFFFF) & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp13_i19_stall_local;
wire local_bb4_cmp13_i19;

assign local_bb4_cmp13_i19 = ((local_bb4_and10_i17 & 32'hFFFF) > (local_bb4_and12_i18 & 32'hFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_var__u73_0_valid_out_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u73_0_stall_in_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u73_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u73_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u73_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u73_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u73_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u73_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_var__u73_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_var__u73_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_var__u73_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_var__u73_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_var__u73_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(rnode_235to236_bb4_var__u73_0_NO_SHIFT_REG),
	.data_out(rnode_236to237_bb4_var__u73_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_var__u73_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_var__u73_0_reg_237_fifo.DATA_WIDTH = 1;
defparam rnode_236to237_bb4_var__u73_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_var__u73_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_var__u73_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_var__u73_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u73_0_NO_SHIFT_REG = rnode_236to237_bb4_var__u73_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_var__u73_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u73_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_235to236_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and193_i_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and193_i_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and193_i_2_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and193_i_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_valid_out_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_stall_in_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and193_i_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_235to236_bb4_and193_i_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to236_bb4_and193_i_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to236_bb4_and193_i_0_stall_in_0_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_235to236_bb4_and193_i_0_valid_out_0_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_235to236_bb4_and193_i_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in((local_bb4_and193_i & 32'hFFFFFFF)),
	.data_out(rnode_235to236_bb4_and193_i_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_235to236_bb4_and193_i_0_reg_236_fifo.DEPTH = 1;
defparam rnode_235to236_bb4_and193_i_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_235to236_bb4_and193_i_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to236_bb4_and193_i_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_235to236_bb4_and193_i_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and193_i_stall_in = 1'b0;
assign rnode_235to236_bb4_and193_i_0_stall_in_0_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_and193_i_0_NO_SHIFT_REG = rnode_235to236_bb4_and193_i_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_and193_i_1_NO_SHIFT_REG = rnode_235to236_bb4_and193_i_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4_and193_i_2_NO_SHIFT_REG = rnode_235to236_bb4_and193_i_0_reg_236_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_235to236_bb4_and195_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and195_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and195_i_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and195_i_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and195_i_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and195_i_0_valid_out_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and195_i_0_stall_in_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and195_i_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_235to236_bb4_and195_i_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to236_bb4_and195_i_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to236_bb4_and195_i_0_stall_in_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_235to236_bb4_and195_i_0_valid_out_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_235to236_bb4_and195_i_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in((local_bb4_and195_i & 32'h1F)),
	.data_out(rnode_235to236_bb4_and195_i_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_235to236_bb4_and195_i_0_reg_236_fifo.DEPTH = 1;
defparam rnode_235to236_bb4_and195_i_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_235to236_bb4_and195_i_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to236_bb4_and195_i_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_235to236_bb4_and195_i_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and195_i_stall_in = 1'b0;
assign rnode_235to236_bb4_and195_i_0_NO_SHIFT_REG = rnode_235to236_bb4_and195_i_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_and195_i_0_stall_in_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and195_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_235to236_bb4_and198_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and198_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and198_i_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and198_i_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4_and198_i_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and198_i_0_valid_out_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and198_i_0_stall_in_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4_and198_i_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_235to236_bb4_and198_i_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to236_bb4_and198_i_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to236_bb4_and198_i_0_stall_in_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_235to236_bb4_and198_i_0_valid_out_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_235to236_bb4_and198_i_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in((local_bb4_and198_i & 32'h1)),
	.data_out(rnode_235to236_bb4_and198_i_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_235to236_bb4_and198_i_0_reg_236_fifo.DEPTH = 1;
defparam rnode_235to236_bb4_and198_i_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_235to236_bb4_and198_i_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to236_bb4_and198_i_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_235to236_bb4_and198_i_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and198_i_stall_in = 1'b0;
assign rnode_235to236_bb4_and198_i_0_NO_SHIFT_REG = rnode_235to236_bb4_and198_i_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4_and198_i_0_stall_in_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and198_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i_stall_local;
wire [31:0] local_bb4_shr_i_i;

assign local_bb4_shr_i_i = ((local_bb4_and201_i & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4__26_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_valid_out_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_stall_in_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__26_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4__26_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4__26_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4__26_i_0_stall_in_0_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4__26_i_0_valid_out_0_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4__26_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(rnode_235to237_bb4__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_237to238_bb4__26_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4__26_i_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4__26_i_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_237to238_bb4__26_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4__26_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4__26_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_235to237_bb4__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__26_i_0_stall_in_0_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__26_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__26_i_0_NO_SHIFT_REG = rnode_237to238_bb4__26_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4__26_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__26_i_1_NO_SHIFT_REG = rnode_237to238_bb4__26_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4__26_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__26_i_2_NO_SHIFT_REG = rnode_237to238_bb4__26_i_0_reg_238_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp_i15_stall_local;
wire local_bb4_cmp_i15;

assign local_bb4_cmp_i15 = ((local_bb4_shr_i12 & 32'h7FFF) > (local_bb4_shr3_i14 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cmp8_i16_stall_local;
wire local_bb4_cmp8_i16;

assign local_bb4_cmp8_i16 = ((local_bb4_shr_i12 & 32'h7FFF) == (local_bb4_shr3_i14 & 32'h7FFF));

// This section implements an unregistered operation.
// 
wire local_bb4_shr216_i_stall_local;
wire [31:0] local_bb4_shr216_i;

assign local_bb4_shr216_i = ((rnode_235to236_bb4_and193_i_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i_stall_local;
wire [31:0] local_bb4__pre_i;

assign local_bb4__pre_i = ((rnode_235to236_bb4_and195_i_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i_stall_local;
wire [31:0] local_bb4_or_i_i;

assign local_bb4_or_i_i = ((local_bb4_shr_i_i & 32'h3FFFFFF) | (local_bb4_and201_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond292_i_stall_local;
wire [31:0] local_bb4_cond292_i;

assign local_bb4_cond292_i = (rnode_237to238_bb4__26_i_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u82_stall_local;
wire [31:0] local_bb4_var__u82;

assign local_bb4_var__u82[31:1] = 31'h0;
assign local_bb4_var__u82[0] = rnode_237to238_bb4__26_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4___i20_stall_local;
wire local_bb4___i20;

assign local_bb4___i20 = (local_bb4_cmp8_i16 & local_bb4_cmp13_i19);

// This section implements an unregistered operation.
// 
wire local_bb4_or219_i_stall_local;
wire [31:0] local_bb4_or219_i;

assign local_bb4_or219_i = ((local_bb4_shr216_i & 32'h7FFFFFF) | (rnode_235to236_bb4_and198_i_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool213_i_stall_local;
wire local_bb4_tobool213_i;

assign local_bb4_tobool213_i = ((local_bb4__pre_i & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i_stall_local;
wire [31:0] local_bb4_shr1_i_i;

assign local_bb4_shr1_i_i = ((local_bb4_or_i_i & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i_stall_local;
wire [31:0] local_bb4_lnot_ext_i;

assign local_bb4_lnot_ext_i = ((local_bb4_var__u82 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u46_valid_out_2;
wire local_bb4_var__u46_stall_in_2;
wire local_bb4__21_i21_valid_out;
wire local_bb4__21_i21_stall_in;
wire local_bb4__21_i21_inputs_ready;
wire local_bb4__21_i21_stall_local;
wire local_bb4__21_i21;

assign local_bb4__21_i21_inputs_ready = (rnode_235to236_bb4_t_322_pop8_c1_ene3_0_valid_out_0_NO_SHIFT_REG & rnode_235to236_bb4_var__u81_0_valid_out_1_NO_SHIFT_REG & rnode_235to236_bb4_var__u81_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__21_i21 = (local_bb4_cmp_i15 | local_bb4___i20);
assign local_bb4_var__u46_valid_out_2 = 1'b1;
assign local_bb4__21_i21_valid_out = 1'b1;
assign rnode_235to236_bb4_t_322_pop8_c1_ene3_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_var__u81_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_var__u81_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i_stall_local;
wire local_bb4__40_demorgan_i;

assign local_bb4__40_demorgan_i = (rnode_234to236_bb4_cmp37_i_0_NO_SHIFT_REG | local_bb4_tobool213_i);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i_stall_local;
wire local_bb4__42_i;

assign local_bb4__42_i = (local_bb4_tobool213_i & local_bb4_not_cmp37_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i_stall_local;
wire [31:0] local_bb4_or2_i_i;

assign local_bb4_or2_i_i = ((local_bb4_shr1_i_i & 32'h1FFFFFF) | (local_bb4_or_i_i & 32'h7FFFFFF));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_var__u46_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u46_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_var__u46_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u46_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u46_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_var__u46_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u46_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_var__u46_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u46_0_valid_out_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u46_0_stall_in_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_var__u46_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_var__u46_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_var__u46_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_var__u46_0_stall_in_0_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_var__u46_0_valid_out_0_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_var__u46_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(local_bb4_var__u46),
	.data_out(rnode_236to237_bb4_var__u46_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_var__u46_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_var__u46_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_236to237_bb4_var__u46_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_var__u46_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_var__u46_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u46_stall_in_2 = 1'b0;
assign rnode_236to237_bb4_var__u46_0_stall_in_0_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u46_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4_var__u46_0_NO_SHIFT_REG = rnode_236to237_bb4_var__u46_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_var__u46_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4_var__u46_1_NO_SHIFT_REG = rnode_236to237_bb4_var__u46_0_reg_237_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4__21_i21_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_valid_out_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_stall_in_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4__21_i21_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4__21_i21_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4__21_i21_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4__21_i21_0_stall_in_0_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4__21_i21_0_valid_out_0_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4__21_i21_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(local_bb4__21_i21),
	.data_out(rnode_236to237_bb4__21_i21_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4__21_i21_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4__21_i21_0_reg_237_fifo.DATA_WIDTH = 1;
defparam rnode_236to237_bb4__21_i21_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4__21_i21_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4__21_i21_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__21_i21_stall_in = 1'b0;
assign rnode_236to237_bb4__21_i21_0_stall_in_0_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4__21_i21_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4__21_i21_0_NO_SHIFT_REG = rnode_236to237_bb4__21_i21_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4__21_i21_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4__21_i21_1_NO_SHIFT_REG = rnode_236to237_bb4__21_i21_0_reg_237_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__43_i_stall_local;
wire [31:0] local_bb4__43_i;

assign local_bb4__43_i = (local_bb4__42_i ? 32'h0 : (local_bb4__pre_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i_stall_local;
wire [31:0] local_bb4_shr3_i_i;

assign local_bb4_shr3_i_i = ((local_bb4_or2_i_i & 32'h7FFFFFF) >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4__22_i22_stall_local;
wire [31:0] local_bb4__22_i22;

assign local_bb4__22_i22 = (rnode_236to237_bb4__21_i21_0_NO_SHIFT_REG ? rnode_236to237_bb4_var__u46_0_NO_SHIFT_REG : rnode_236to237_bb4_var__u81_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4__23_i23_stall_local;
wire [31:0] local_bb4__23_i23;

assign local_bb4__23_i23 = (rnode_236to237_bb4__21_i21_1_NO_SHIFT_REG ? rnode_236to237_bb4_var__u81_1_NO_SHIFT_REG : rnode_236to237_bb4_var__u46_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i_stall_local;
wire [31:0] local_bb4_or4_i_i;

assign local_bb4_or4_i_i = ((local_bb4_shr3_i_i & 32'h7FFFFF) | (local_bb4_or2_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_shr18_i26_stall_local;
wire [31:0] local_bb4_shr18_i26;

assign local_bb4_shr18_i26 = (local_bb4__22_i22 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr16_i24_stall_local;
wire [31:0] local_bb4_shr16_i24;

assign local_bb4_shr16_i24 = (local_bb4__23_i23 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i_stall_local;
wire [31:0] local_bb4_shr5_i_i;

assign local_bb4_shr5_i_i = ((local_bb4_or4_i_i & 32'h7FFFFFF) >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and19_i27_stall_local;
wire [31:0] local_bb4_and19_i27;

assign local_bb4_and19_i27 = ((local_bb4_shr18_i26 & 32'h1FF) & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_sub_i56_stall_local;
wire [31:0] local_bb4_sub_i56;

assign local_bb4_sub_i56 = ((local_bb4_shr16_i24 & 32'h1FF) - (local_bb4_shr18_i26 & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i_stall_local;
wire [31:0] local_bb4_or6_i_i;

assign local_bb4_or6_i_i = ((local_bb4_shr5_i_i & 32'h7FFFF) | (local_bb4_or4_i_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot23_i31_stall_local;
wire local_bb4_lnot23_i31;

assign local_bb4_lnot23_i31 = ((local_bb4_and19_i27 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp27_i33_stall_local;
wire local_bb4_cmp27_i33;

assign local_bb4_cmp27_i33 = ((local_bb4_and19_i27 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and68_i57_stall_local;
wire [31:0] local_bb4_and68_i57;

assign local_bb4_and68_i57 = (local_bb4_sub_i56 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i_stall_local;
wire [31:0] local_bb4_shr7_i_i;

assign local_bb4_shr7_i_i = ((local_bb4_or6_i_i & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i_stall_local;
wire [31:0] local_bb4_or6_masked_i_i;

assign local_bb4_or6_masked_i_i = ((local_bb4_or6_i_i & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp69_i58_stall_local;
wire local_bb4_cmp69_i58;

assign local_bb4_cmp69_i58 = ((local_bb4_and68_i57 & 32'hFF) > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i_stall_local;
wire [31:0] local_bb4_neg_i_i;

assign local_bb4_neg_i_i = ((local_bb4_or6_masked_i_i & 32'h7FFFFFF) | (local_bb4_shr7_i_i & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb4__22_i22_valid_out_1;
wire local_bb4__22_i22_stall_in_1;
wire local_bb4__23_i23_valid_out_1;
wire local_bb4__23_i23_stall_in_1;
wire local_bb4_shr16_i24_valid_out_1;
wire local_bb4_shr16_i24_stall_in_1;
wire local_bb4_lnot23_i31_valid_out;
wire local_bb4_lnot23_i31_stall_in;
wire local_bb4_cmp27_i33_valid_out;
wire local_bb4_cmp27_i33_stall_in;
wire local_bb4_align_0_i59_valid_out;
wire local_bb4_align_0_i59_stall_in;
wire local_bb4_align_0_i59_inputs_ready;
wire local_bb4_align_0_i59_stall_local;
wire [31:0] local_bb4_align_0_i59;

assign local_bb4_align_0_i59_inputs_ready = (rnode_236to237_bb4__21_i21_0_valid_out_0_NO_SHIFT_REG & rnode_236to237_bb4_var__u46_0_valid_out_0_NO_SHIFT_REG & rnode_236to237_bb4_var__u81_0_valid_out_0_NO_SHIFT_REG & rnode_236to237_bb4__21_i21_0_valid_out_1_NO_SHIFT_REG & rnode_236to237_bb4_var__u46_0_valid_out_1_NO_SHIFT_REG & rnode_236to237_bb4_var__u81_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_align_0_i59 = (local_bb4_cmp69_i58 ? 32'h1F : (local_bb4_and68_i57 & 32'hFF));
assign local_bb4__22_i22_valid_out_1 = 1'b1;
assign local_bb4__23_i23_valid_out_1 = 1'b1;
assign local_bb4_shr16_i24_valid_out_1 = 1'b1;
assign local_bb4_lnot23_i31_valid_out = 1'b1;
assign local_bb4_cmp27_i33_valid_out = 1'b1;
assign local_bb4_align_0_i59_valid_out = 1'b1;
assign rnode_236to237_bb4__21_i21_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u46_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u81_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4__21_i21_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u46_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u81_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i9_stall_local;
wire [31:0] local_bb4_and_i_i9;

assign local_bb4_and_i_i9 = ((local_bb4_neg_i_i & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4__22_i22_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__22_i22_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4__22_i22_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__22_i22_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__22_i22_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4__22_i22_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__22_i22_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4__22_i22_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__22_i22_0_valid_out_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__22_i22_0_stall_in_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__22_i22_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4__22_i22_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4__22_i22_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4__22_i22_0_stall_in_0_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4__22_i22_0_valid_out_0_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4__22_i22_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(local_bb4__22_i22),
	.data_out(rnode_237to238_bb4__22_i22_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4__22_i22_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4__22_i22_0_reg_238_fifo.DATA_WIDTH = 32;
defparam rnode_237to238_bb4__22_i22_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4__22_i22_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4__22_i22_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__22_i22_stall_in_1 = 1'b0;
assign rnode_237to238_bb4__22_i22_0_stall_in_0_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__22_i22_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__22_i22_0_NO_SHIFT_REG = rnode_237to238_bb4__22_i22_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4__22_i22_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__22_i22_1_NO_SHIFT_REG = rnode_237to238_bb4__22_i22_0_reg_238_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4__23_i23_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4__23_i23_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4__23_i23_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4__23_i23_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4__23_i23_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_valid_out_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_stall_in_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__23_i23_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4__23_i23_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4__23_i23_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4__23_i23_0_stall_in_0_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4__23_i23_0_valid_out_0_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4__23_i23_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(local_bb4__23_i23),
	.data_out(rnode_237to238_bb4__23_i23_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4__23_i23_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4__23_i23_0_reg_238_fifo.DATA_WIDTH = 32;
defparam rnode_237to238_bb4__23_i23_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4__23_i23_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4__23_i23_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__23_i23_stall_in_1 = 1'b0;
assign rnode_237to238_bb4__23_i23_0_stall_in_0_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__23_i23_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__23_i23_0_NO_SHIFT_REG = rnode_237to238_bb4__23_i23_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4__23_i23_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__23_i23_1_NO_SHIFT_REG = rnode_237to238_bb4__23_i23_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4__23_i23_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__23_i23_2_NO_SHIFT_REG = rnode_237to238_bb4__23_i23_0_reg_238_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_237to239_bb4_shr16_i24_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to239_bb4_shr16_i24_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_237to239_bb4_shr16_i24_0_NO_SHIFT_REG;
 logic rnode_237to239_bb4_shr16_i24_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to239_bb4_shr16_i24_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_237to239_bb4_shr16_i24_1_NO_SHIFT_REG;
 logic rnode_237to239_bb4_shr16_i24_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to239_bb4_shr16_i24_0_reg_239_NO_SHIFT_REG;
 logic rnode_237to239_bb4_shr16_i24_0_valid_out_0_reg_239_NO_SHIFT_REG;
 logic rnode_237to239_bb4_shr16_i24_0_stall_in_0_reg_239_NO_SHIFT_REG;
 logic rnode_237to239_bb4_shr16_i24_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_237to239_bb4_shr16_i24_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to239_bb4_shr16_i24_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to239_bb4_shr16_i24_0_stall_in_0_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_237to239_bb4_shr16_i24_0_valid_out_0_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_237to239_bb4_shr16_i24_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in((local_bb4_shr16_i24 & 32'h1FF)),
	.data_out(rnode_237to239_bb4_shr16_i24_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_237to239_bb4_shr16_i24_0_reg_239_fifo.DEPTH = 2;
defparam rnode_237to239_bb4_shr16_i24_0_reg_239_fifo.DATA_WIDTH = 32;
defparam rnode_237to239_bb4_shr16_i24_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to239_bb4_shr16_i24_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_237to239_bb4_shr16_i24_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr16_i24_stall_in_1 = 1'b0;
assign rnode_237to239_bb4_shr16_i24_0_stall_in_0_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_237to239_bb4_shr16_i24_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to239_bb4_shr16_i24_0_NO_SHIFT_REG = rnode_237to239_bb4_shr16_i24_0_reg_239_NO_SHIFT_REG;
assign rnode_237to239_bb4_shr16_i24_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to239_bb4_shr16_i24_1_NO_SHIFT_REG = rnode_237to239_bb4_shr16_i24_0_reg_239_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_lnot23_i31_0_valid_out_NO_SHIFT_REG;
 logic rnode_237to238_bb4_lnot23_i31_0_stall_in_NO_SHIFT_REG;
 logic rnode_237to238_bb4_lnot23_i31_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_lnot23_i31_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to238_bb4_lnot23_i31_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_lnot23_i31_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_lnot23_i31_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_lnot23_i31_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_lnot23_i31_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_lnot23_i31_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_lnot23_i31_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_lnot23_i31_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_lnot23_i31_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(local_bb4_lnot23_i31),
	.data_out(rnode_237to238_bb4_lnot23_i31_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_lnot23_i31_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_lnot23_i31_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_237to238_bb4_lnot23_i31_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_lnot23_i31_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_lnot23_i31_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot23_i31_stall_in = 1'b0;
assign rnode_237to238_bb4_lnot23_i31_0_NO_SHIFT_REG = rnode_237to238_bb4_lnot23_i31_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_lnot23_i31_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_lnot23_i31_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_237to239_bb4_cmp27_i33_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_1_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_2_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_reg_239_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_valid_out_0_reg_239_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_stall_in_0_reg_239_NO_SHIFT_REG;
 logic rnode_237to239_bb4_cmp27_i33_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_237to239_bb4_cmp27_i33_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to239_bb4_cmp27_i33_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to239_bb4_cmp27_i33_0_stall_in_0_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_237to239_bb4_cmp27_i33_0_valid_out_0_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_237to239_bb4_cmp27_i33_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in(local_bb4_cmp27_i33),
	.data_out(rnode_237to239_bb4_cmp27_i33_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_237to239_bb4_cmp27_i33_0_reg_239_fifo.DEPTH = 2;
defparam rnode_237to239_bb4_cmp27_i33_0_reg_239_fifo.DATA_WIDTH = 1;
defparam rnode_237to239_bb4_cmp27_i33_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to239_bb4_cmp27_i33_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_237to239_bb4_cmp27_i33_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp27_i33_stall_in = 1'b0;
assign rnode_237to239_bb4_cmp27_i33_0_stall_in_0_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_237to239_bb4_cmp27_i33_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to239_bb4_cmp27_i33_0_NO_SHIFT_REG = rnode_237to239_bb4_cmp27_i33_0_reg_239_NO_SHIFT_REG;
assign rnode_237to239_bb4_cmp27_i33_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to239_bb4_cmp27_i33_1_NO_SHIFT_REG = rnode_237to239_bb4_cmp27_i33_0_reg_239_NO_SHIFT_REG;
assign rnode_237to239_bb4_cmp27_i33_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_237to239_bb4_cmp27_i33_2_NO_SHIFT_REG = rnode_237to239_bb4_cmp27_i33_0_reg_239_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_align_0_i59_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_align_0_i59_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_align_0_i59_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_align_0_i59_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_align_0_i59_3_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_align_0_i59_4_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_align_0_i59_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_valid_out_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_stall_in_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_align_0_i59_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_align_0_i59_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_align_0_i59_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_align_0_i59_0_stall_in_0_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_align_0_i59_0_valid_out_0_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_align_0_i59_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in((local_bb4_align_0_i59 & 32'hFF)),
	.data_out(rnode_237to238_bb4_align_0_i59_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_align_0_i59_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_align_0_i59_0_reg_238_fifo.DATA_WIDTH = 32;
defparam rnode_237to238_bb4_align_0_i59_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_align_0_i59_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_align_0_i59_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_align_0_i59_stall_in = 1'b0;
assign rnode_237to238_bb4_align_0_i59_0_stall_in_0_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_align_0_i59_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_align_0_i59_0_NO_SHIFT_REG = rnode_237to238_bb4_align_0_i59_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_align_0_i59_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_align_0_i59_1_NO_SHIFT_REG = rnode_237to238_bb4_align_0_i59_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_align_0_i59_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_align_0_i59_2_NO_SHIFT_REG = rnode_237to238_bb4_align_0_i59_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_align_0_i59_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_align_0_i59_3_NO_SHIFT_REG = rnode_237to238_bb4_align_0_i59_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_align_0_i59_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_align_0_i59_4_NO_SHIFT_REG = rnode_237to238_bb4_align_0_i59_0_reg_238_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i9_valid_out;
wire local_bb4__and_i_i9_stall_in;
wire local_bb4__and_i_i9_inputs_ready;
wire local_bb4__and_i_i9_stall_local;
wire [31:0] local_bb4__and_i_i9;

thirtysix_six_comp local_bb4__and_i_i9_popcnt_instance (
	.data((local_bb4_and_i_i9 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i9)
);


assign local_bb4__and_i_i9_inputs_ready = rnode_234to235_bb4_add192_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i9_valid_out = 1'b1;
assign rnode_234to235_bb4_add192_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and21_i29_stall_local;
wire [31:0] local_bb4_and21_i29;

assign local_bb4_and21_i29 = (rnode_237to238_bb4__22_i22_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and20_i28_valid_out;
wire local_bb4_and20_i28_stall_in;
wire local_bb4_and20_i28_inputs_ready;
wire local_bb4_and20_i28_stall_local;
wire [31:0] local_bb4_and20_i28;

assign local_bb4_and20_i28_inputs_ready = rnode_237to238_bb4__23_i23_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and20_i28 = (rnode_237to238_bb4__23_i23_0_NO_SHIFT_REG & 32'h7FFFFF);
assign local_bb4_and20_i28_valid_out = 1'b1;
assign rnode_237to238_bb4__23_i23_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and35_i34_valid_out;
wire local_bb4_and35_i34_stall_in;
wire local_bb4_and35_i34_inputs_ready;
wire local_bb4_and35_i34_stall_local;
wire [31:0] local_bb4_and35_i34;

assign local_bb4_and35_i34_inputs_ready = rnode_237to238_bb4__23_i23_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and35_i34 = (rnode_237to238_bb4__23_i23_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb4_and35_i34_valid_out = 1'b1;
assign rnode_237to238_bb4__23_i23_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_xor_i35_stall_local;
wire [31:0] local_bb4_xor_i35;

assign local_bb4_xor_i35 = (rnode_237to238_bb4__23_i23_2_NO_SHIFT_REG ^ rnode_237to238_bb4__22_i22_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i25_stall_local;
wire [31:0] local_bb4_and17_i25;

assign local_bb4_and17_i25 = ((rnode_237to239_bb4_shr16_i24_0_NO_SHIFT_REG & 32'h1FF) & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_239to241_bb4_shr16_i24_0_valid_out_NO_SHIFT_REG;
 logic rnode_239to241_bb4_shr16_i24_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_239to241_bb4_shr16_i24_0_NO_SHIFT_REG;
 logic rnode_239to241_bb4_shr16_i24_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_239to241_bb4_shr16_i24_0_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_shr16_i24_0_valid_out_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_shr16_i24_0_stall_in_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_shr16_i24_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_239to241_bb4_shr16_i24_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to241_bb4_shr16_i24_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to241_bb4_shr16_i24_0_stall_in_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_239to241_bb4_shr16_i24_0_valid_out_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_239to241_bb4_shr16_i24_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in((rnode_237to239_bb4_shr16_i24_1_NO_SHIFT_REG & 32'h1FF)),
	.data_out(rnode_239to241_bb4_shr16_i24_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_239to241_bb4_shr16_i24_0_reg_241_fifo.DEPTH = 2;
defparam rnode_239to241_bb4_shr16_i24_0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_239to241_bb4_shr16_i24_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to241_bb4_shr16_i24_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_239to241_bb4_shr16_i24_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_237to239_bb4_shr16_i24_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_shr16_i24_0_NO_SHIFT_REG = rnode_239to241_bb4_shr16_i24_0_reg_241_NO_SHIFT_REG;
assign rnode_239to241_bb4_shr16_i24_0_stall_in_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_shr16_i24_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and93_i67_stall_local;
wire [31:0] local_bb4_and93_i67;

assign local_bb4_and93_i67 = ((rnode_237to238_bb4_align_0_i59_0_NO_SHIFT_REG & 32'hFF) & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb4_and95_i69_stall_local;
wire [31:0] local_bb4_and95_i69;

assign local_bb4_and95_i69 = ((rnode_237to238_bb4_align_0_i59_1_NO_SHIFT_REG & 32'hFF) & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_and115_i85_stall_local;
wire [31:0] local_bb4_and115_i85;

assign local_bb4_and115_i85 = ((rnode_237to238_bb4_align_0_i59_2_NO_SHIFT_REG & 32'hFF) & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb4_and130_i91_stall_local;
wire [31:0] local_bb4_and130_i91;

assign local_bb4_and130_i91 = ((rnode_237to238_bb4_align_0_i59_3_NO_SHIFT_REG & 32'hFF) & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_and149_i96_stall_local;
wire [31:0] local_bb4_and149_i96;

assign local_bb4_and149_i96 = ((rnode_237to238_bb4_align_0_i59_4_NO_SHIFT_REG & 32'hFF) & 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_235to236_bb4__and_i_i9_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4__and_i_i9_0_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4__and_i_i9_1_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4__and_i_i9_2_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_reg_236_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_235to236_bb4__and_i_i9_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_valid_out_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_stall_in_0_reg_236_NO_SHIFT_REG;
 logic rnode_235to236_bb4__and_i_i9_0_stall_out_reg_236_NO_SHIFT_REG;

acl_data_fifo rnode_235to236_bb4__and_i_i9_0_reg_236_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_235to236_bb4__and_i_i9_0_reg_236_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_235to236_bb4__and_i_i9_0_stall_in_0_reg_236_NO_SHIFT_REG),
	.valid_out(rnode_235to236_bb4__and_i_i9_0_valid_out_0_reg_236_NO_SHIFT_REG),
	.stall_out(rnode_235to236_bb4__and_i_i9_0_stall_out_reg_236_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i9 & 32'h3F)),
	.data_out(rnode_235to236_bb4__and_i_i9_0_reg_236_NO_SHIFT_REG)
);

defparam rnode_235to236_bb4__and_i_i9_0_reg_236_fifo.DEPTH = 1;
defparam rnode_235to236_bb4__and_i_i9_0_reg_236_fifo.DATA_WIDTH = 32;
defparam rnode_235to236_bb4__and_i_i9_0_reg_236_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_235to236_bb4__and_i_i9_0_reg_236_fifo.IMPL = "shift_reg";

assign rnode_235to236_bb4__and_i_i9_0_reg_236_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i9_stall_in = 1'b0;
assign rnode_235to236_bb4__and_i_i9_0_stall_in_0_reg_236_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4__and_i_i9_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4__and_i_i9_0_NO_SHIFT_REG = rnode_235to236_bb4__and_i_i9_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4__and_i_i9_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4__and_i_i9_1_NO_SHIFT_REG = rnode_235to236_bb4__and_i_i9_0_reg_236_NO_SHIFT_REG;
assign rnode_235to236_bb4__and_i_i9_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_235to236_bb4__and_i_i9_2_NO_SHIFT_REG = rnode_235to236_bb4__and_i_i9_0_reg_236_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i40_stall_local;
wire local_bb4_lnot33_not_i40;

assign local_bb4_lnot33_not_i40 = ((local_bb4_and21_i29 & 32'h7FFFFF) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or64_i53_stall_local;
wire [31:0] local_bb4_or64_i53;

assign local_bb4_or64_i53 = ((local_bb4_and21_i29 & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_and20_i28_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and20_i28_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_and20_i28_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and20_i28_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and20_i28_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_and20_i28_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and20_i28_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_and20_i28_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and20_i28_0_valid_out_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and20_i28_0_stall_in_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and20_i28_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_and20_i28_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_and20_i28_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_and20_i28_0_stall_in_0_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_and20_i28_0_valid_out_0_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_and20_i28_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in((local_bb4_and20_i28 & 32'h7FFFFF)),
	.data_out(rnode_238to239_bb4_and20_i28_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_and20_i28_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_and20_i28_0_reg_239_fifo.DATA_WIDTH = 32;
defparam rnode_238to239_bb4_and20_i28_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_and20_i28_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_and20_i28_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and20_i28_stall_in = 1'b0;
assign rnode_238to239_bb4_and20_i28_0_stall_in_0_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_and20_i28_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_and20_i28_0_NO_SHIFT_REG = rnode_238to239_bb4_and20_i28_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_and20_i28_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_and20_i28_1_NO_SHIFT_REG = rnode_238to239_bb4_and20_i28_0_reg_239_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_and35_i34_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and35_i34_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_and35_i34_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and35_i34_0_valid_out_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and35_i34_0_stall_in_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and35_i34_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_and35_i34_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_and35_i34_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_and35_i34_0_stall_in_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_and35_i34_0_valid_out_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_and35_i34_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in((local_bb4_and35_i34 & 32'h80000000)),
	.data_out(rnode_238to239_bb4_and35_i34_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_and35_i34_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_and35_i34_0_reg_239_fifo.DATA_WIDTH = 32;
defparam rnode_238to239_bb4_and35_i34_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_and35_i34_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_and35_i34_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and35_i34_stall_in = 1'b0;
assign rnode_238to239_bb4_and35_i34_0_NO_SHIFT_REG = rnode_238to239_bb4_and35_i34_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_and35_i34_0_stall_in_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp37_i36_stall_local;
wire local_bb4_cmp37_i36;

assign local_bb4_cmp37_i36 = ($signed(local_bb4_xor_i35) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb4_xor_lobit_i109_stall_local;
wire [31:0] local_bb4_xor_lobit_i109;

assign local_bb4_xor_lobit_i109 = ($signed(local_bb4_xor_i35) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and36_lobit_i111_stall_local;
wire [31:0] local_bb4_and36_lobit_i111;

assign local_bb4_and36_lobit_i111 = (local_bb4_xor_i35 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_i30_stall_local;
wire local_bb4_lnot_i30;

assign local_bb4_lnot_i30 = ((local_bb4_and17_i25 & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_i32_stall_local;
wire local_bb4_cmp25_i32;

assign local_bb4_cmp25_i32 = ((local_bb4_and17_i25 & 32'hFF) == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp96_i70_stall_local;
wire local_bb4_cmp96_i70;

assign local_bb4_cmp96_i70 = ((local_bb4_and95_i69 & 32'h10) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp116_i86_stall_local;
wire local_bb4_cmp116_i86;

assign local_bb4_cmp116_i86 = ((local_bb4_and115_i85 & 32'h8) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp131_not_i93_stall_local;
wire local_bb4_cmp131_not_i93;

assign local_bb4_cmp131_not_i93 = ((local_bb4_and130_i91 & 32'h4) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_Pivot20_i98_stall_local;
wire local_bb4_Pivot20_i98;

assign local_bb4_Pivot20_i98 = ((local_bb4_and149_i96 & 32'h3) < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_SwitchLeaf_i99_stall_local;
wire local_bb4_SwitchLeaf_i99;

assign local_bb4_SwitchLeaf_i99 = ((local_bb4_and149_i96 & 32'h3) == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i_stall_local;
wire [31:0] local_bb4_and9_i_i;

assign local_bb4_and9_i_i = ((rnode_235to236_bb4__and_i_i9_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and203_i_stall_local;
wire [31:0] local_bb4_and203_i;

assign local_bb4_and203_i = ((rnode_235to236_bb4__and_i_i9_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i_stall_local;
wire [31:0] local_bb4_and206_i;

assign local_bb4_and206_i = ((rnode_235to236_bb4__and_i_i9_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shl65_i54_stall_local;
wire [31:0] local_bb4_shl65_i54;

assign local_bb4_shl65_i54 = ((local_bb4_or64_i53 & 32'h3FFFFF8) | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_i38_stall_local;
wire local_bb4_lnot30_i38;

assign local_bb4_lnot30_i38 = ((rnode_238to239_bb4_and20_i28_0_NO_SHIFT_REG & 32'h7FFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i50_stall_local;
wire [31:0] local_bb4_or_i50;

assign local_bb4_or_i50 = ((rnode_238to239_bb4_and20_i28_1_NO_SHIFT_REG & 32'h7FFFFF) << 32'h3);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_239to241_bb4_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_239to241_bb4_and35_i34_0_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and35_i34_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_239to241_bb4_and35_i34_0_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and35_i34_0_valid_out_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and35_i34_0_stall_in_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and35_i34_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_239to241_bb4_and35_i34_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to241_bb4_and35_i34_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to241_bb4_and35_i34_0_stall_in_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_239to241_bb4_and35_i34_0_valid_out_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_239to241_bb4_and35_i34_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in((rnode_238to239_bb4_and35_i34_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_239to241_bb4_and35_i34_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_239to241_bb4_and35_i34_0_reg_241_fifo.DEPTH = 2;
defparam rnode_239to241_bb4_and35_i34_0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_239to241_bb4_and35_i34_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to241_bb4_and35_i34_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_239to241_bb4_and35_i34_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_and35_i34_0_NO_SHIFT_REG = rnode_239to241_bb4_and35_i34_0_reg_241_NO_SHIFT_REG;
assign rnode_239to241_bb4_and35_i34_0_stall_in_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_cmp25_not_i37_stall_local;
wire local_bb4_cmp25_not_i37;

assign local_bb4_cmp25_not_i37 = (local_bb4_cmp25_i32 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u83_stall_local;
wire local_bb4_var__u83;

assign local_bb4_var__u83 = (local_bb4_cmp25_i32 | rnode_237to239_bb4_cmp27_i33_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_sub239_i_stall_local;
wire [31:0] local_bb4_sub239_i;

assign local_bb4_sub239_i = (32'h0 - (local_bb4_and9_i_i & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl204_i_stall_local;
wire [31:0] local_bb4_shl204_i;

assign local_bb4_shl204_i = ((rnode_235to236_bb4_and193_i_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and203_i & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb4__28_i55_stall_local;
wire [31:0] local_bb4__28_i55;

assign local_bb4__28_i55 = (rnode_237to238_bb4_lnot23_i31_0_NO_SHIFT_REG ? 32'h0 : ((local_bb4_shl65_i54 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot30_not_i42_stall_local;
wire local_bb4_lnot30_not_i42;

assign local_bb4_lnot30_not_i42 = (local_bb4_lnot30_i38 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_shl_i51_stall_local;
wire [31:0] local_bb4_shl_i51;

assign local_bb4_shl_i51 = ((local_bb4_or_i50 & 32'h3FFFFF8) | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_241to242_bb4_and35_i34_0_valid_out_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and35_i34_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4_and35_i34_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and35_i34_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4_and35_i34_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and35_i34_0_valid_out_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and35_i34_0_stall_in_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and35_i34_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_241to242_bb4_and35_i34_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to242_bb4_and35_i34_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to242_bb4_and35_i34_0_stall_in_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_241to242_bb4_and35_i34_0_valid_out_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_241to242_bb4_and35_i34_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in((rnode_239to241_bb4_and35_i34_0_NO_SHIFT_REG & 32'h80000000)),
	.data_out(rnode_241to242_bb4_and35_i34_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_241to242_bb4_and35_i34_0_reg_242_fifo.DEPTH = 1;
defparam rnode_241to242_bb4_and35_i34_0_reg_242_fifo.DATA_WIDTH = 32;
defparam rnode_241to242_bb4_and35_i34_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to242_bb4_and35_i34_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_241to242_bb4_and35_i34_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_239to241_bb4_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_and35_i34_0_NO_SHIFT_REG = rnode_241to242_bb4_and35_i34_0_reg_242_NO_SHIFT_REG;
assign rnode_241to242_bb4_and35_i34_0_stall_in_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_and35_i34_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_i39_stall_local;
wire local_bb4_or_cond_i39;

assign local_bb4_or_cond_i39 = (local_bb4_lnot30_i38 | local_bb4_cmp25_not_i37);

// This section implements an unregistered operation.
// 
wire local_bb4_cond244_i_stall_local;
wire [31:0] local_bb4_cond244_i;

assign local_bb4_cond244_i = (rnode_234to236_bb4_cmp37_i_2_NO_SHIFT_REG ? local_bb4_sub239_i : (local_bb4__43_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and205_i_stall_local;
wire [31:0] local_bb4_and205_i;

assign local_bb4_and205_i = (local_bb4_shl204_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and72_i60_stall_local;
wire [31:0] local_bb4_and72_i60;

assign local_bb4_and72_i60 = ((local_bb4__28_i55 & 32'h7FFFFF8) >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb4_and75_i63_stall_local;
wire [31:0] local_bb4_and75_i63;

assign local_bb4_and75_i63 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb4_and78_i65_stall_local;
wire [31:0] local_bb4_and78_i65;

assign local_bb4_and78_i65 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb4_shr94_i68_stall_local;
wire [31:0] local_bb4_shr94_i68;

assign local_bb4_shr94_i68 = ((local_bb4__28_i55 & 32'h7FFFFF8) >> (local_bb4_and93_i67 & 32'h1C));

// This section implements an unregistered operation.
// 
wire local_bb4_and90_i71_stall_local;
wire [31:0] local_bb4_and90_i71;

assign local_bb4_and90_i71 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb4_and87_i72_stall_local;
wire [31:0] local_bb4_and87_i72;

assign local_bb4_and87_i72 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb4_and84_i73_stall_local;
wire [31:0] local_bb4_and84_i73;

assign local_bb4_and84_i73 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u84_stall_local;
wire [31:0] local_bb4_var__u84;

assign local_bb4_var__u84 = ((local_bb4__28_i55 & 32'h7FFFFF8) & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb4_or_cond_not_i43_stall_local;
wire local_bb4_or_cond_not_i43;

assign local_bb4_or_cond_not_i43 = (local_bb4_cmp25_i32 & local_bb4_lnot30_not_i42);

// This section implements an unregistered operation.
// 
wire local_bb4__27_i52_stall_local;
wire [31:0] local_bb4__27_i52;

assign local_bb4__27_i52 = (local_bb4_lnot_i30 ? 32'h0 : ((local_bb4_shl_i51 & 32'h7FFFFF8) | 32'h4000000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_8_i47_stall_local;
wire local_bb4_reduction_8_i47;

assign local_bb4_reduction_8_i47 = (rnode_237to239_bb4_cmp27_i33_1_NO_SHIFT_REG & local_bb4_or_cond_i39);

// This section implements an unregistered operation.
// 
wire local_bb4_add245_i_stall_local;
wire [31:0] local_bb4_add245_i;

assign local_bb4_add245_i = (local_bb4_cond244_i + (rnode_234to236_bb4_and17_i_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i10_stall_local;
wire [31:0] local_bb4_fold_i10;

assign local_bb4_fold_i10 = (local_bb4_cond244_i + (rnode_234to236_bb4_shr16_i_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl207_i_stall_local;
wire [31:0] local_bb4_shl207_i;

assign local_bb4_shl207_i = ((local_bb4_and205_i & 32'h7FFFFFF) << (local_bb4_and206_i & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb4_and72_tr_i61_stall_local;
wire [7:0] local_bb4_and72_tr_i61;
wire [31:0] local_bb4_and72_tr_i61$ps;

assign local_bb4_and72_tr_i61$ps = (local_bb4_and72_i60 & 32'hFFFFFF);
assign local_bb4_and72_tr_i61 = local_bb4_and72_tr_i61$ps[7:0];

// This section implements an unregistered operation.
// 
wire local_bb4_cmp76_i64_stall_local;
wire local_bb4_cmp76_i64;

assign local_bb4_cmp76_i64 = ((local_bb4_and75_i63 & 32'hF0) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp79_i66_stall_local;
wire local_bb4_cmp79_i66;

assign local_bb4_cmp79_i66 = ((local_bb4_and78_i65 & 32'hF00) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and142_i95_stall_local;
wire [31:0] local_bb4_and142_i95;

assign local_bb4_and142_i95 = (local_bb4_shr94_i68 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_shr150_i97_stall_local;
wire [31:0] local_bb4_shr150_i97;

assign local_bb4_shr150_i97 = (local_bb4_shr94_i68 >> (local_bb4_and149_i96 & 32'h3));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u85_stall_local;
wire [31:0] local_bb4_var__u85;

assign local_bb4_var__u85 = (local_bb4_shr94_i68 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and146_i100_stall_local;
wire [31:0] local_bb4_and146_i100;

assign local_bb4_and146_i100 = (local_bb4_shr94_i68 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp91_i74_stall_local;
wire local_bb4_cmp91_i74;

assign local_bb4_cmp91_i74 = ((local_bb4_and90_i71 & 32'h7000000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp88_i75_stall_local;
wire local_bb4_cmp88_i75;

assign local_bb4_cmp88_i75 = ((local_bb4_and87_i72 & 32'hF00000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp85_i76_stall_local;
wire local_bb4_cmp85_i76;

assign local_bb4_cmp85_i76 = ((local_bb4_and84_i73 & 32'hF0000) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u86_stall_local;
wire local_bb4_var__u86;

assign local_bb4_var__u86 = ((local_bb4_var__u84 & 32'hFFF8) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i_stall_local;
wire [31:0] local_bb4_and250_i;

assign local_bb4_and250_i = (local_bb4_fold_i10 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and269_i_stall_local;
wire [31:0] local_bb4_and269_i;

assign local_bb4_and269_i = (local_bb4_fold_i10 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and208_i_stall_local;
wire [31:0] local_bb4_and208_i;

assign local_bb4_and208_i = (local_bb4_shl207_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool74_i62_stall_local;
wire [7:0] local_bb4_frombool74_i62;

assign local_bb4_frombool74_i62 = (local_bb4_and72_tr_i61 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u87_stall_local;
wire [31:0] local_bb4_var__u87;

assign local_bb4_var__u87 = ((local_bb4_and146_i100 & 32'h3FFFFFFF) | local_bb4_shr94_i68);

// This section implements an unregistered operation.
// 
wire local_bb4__31_v_i82_stall_local;
wire local_bb4__31_v_i82;

assign local_bb4__31_v_i82 = (local_bb4_cmp96_i70 ? local_bb4_cmp79_i66 : local_bb4_cmp91_i74);

// This section implements an unregistered operation.
// 
wire local_bb4__30_v_i80_stall_local;
wire local_bb4__30_v_i80;

assign local_bb4__30_v_i80 = (local_bb4_cmp96_i70 ? local_bb4_cmp76_i64 : local_bb4_cmp88_i75);

// This section implements an unregistered operation.
// 
wire local_bb4_frombool109_i78_stall_local;
wire [7:0] local_bb4_frombool109_i78;

assign local_bb4_frombool109_i78[7:1] = 7'h0;
assign local_bb4_frombool109_i78[0] = local_bb4_cmp85_i76;

// This section implements an unregistered operation.
// 
wire local_bb4_or107_i77_stall_local;
wire [31:0] local_bb4_or107_i77;

assign local_bb4_or107_i77[31:1] = 31'h0;
assign local_bb4_or107_i77[0] = local_bb4_var__u86;

// This section implements an unregistered operation.
// 
wire local_bb4__44_i_stall_local;
wire [31:0] local_bb4__44_i;

assign local_bb4__44_i = (local_bb4__40_demorgan_i ? (local_bb4_and208_i & 32'h7FFFFFF) : (local_bb4_or219_i & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_or1596_i101_stall_local;
wire [31:0] local_bb4_or1596_i101;

assign local_bb4_or1596_i101 = (local_bb4_var__u87 | (local_bb4_and142_i95 & 32'h7FFFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4__31_i83_stall_local;
wire [7:0] local_bb4__31_i83;

assign local_bb4__31_i83[7:1] = 7'h0;
assign local_bb4__31_i83[0] = local_bb4__31_v_i82;

// This section implements an unregistered operation.
// 
wire local_bb4__30_i81_stall_local;
wire [7:0] local_bb4__30_i81;

assign local_bb4__30_i81[7:1] = 7'h0;
assign local_bb4__30_i81[0] = local_bb4__30_v_i80;

// This section implements an unregistered operation.
// 
wire local_bb4__29_i79_stall_local;
wire [7:0] local_bb4__29_i79;

assign local_bb4__29_i79 = (local_bb4_cmp96_i70 ? (local_bb4_frombool74_i62 & 8'h1) : (local_bb4_frombool109_i78 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__32_i84_stall_local;
wire [31:0] local_bb4__32_i84;

assign local_bb4__32_i84 = (local_bb4_cmp96_i70 ? 32'h0 : (local_bb4_or107_i77 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i_valid_out;
wire local_bb4_and250_i_stall_in;
wire local_bb4_and269_i_valid_out;
wire local_bb4_and269_i_stall_in;
wire local_bb4_add245_i_valid_out;
wire local_bb4_add245_i_stall_in;
wire local_bb4__45_i_valid_out;
wire local_bb4__45_i_stall_in;
wire local_bb4_not_cmp37_i_valid_out_1;
wire local_bb4_not_cmp37_i_stall_in_1;
wire local_bb4__45_i_inputs_ready;
wire local_bb4__45_i_stall_local;
wire [31:0] local_bb4__45_i;

assign local_bb4__45_i_inputs_ready = (rnode_234to236_bb4_shr16_i_0_valid_out_NO_SHIFT_REG & rnode_234to236_bb4_and17_i_0_valid_out_NO_SHIFT_REG & rnode_234to236_bb4_cmp37_i_0_valid_out_2_NO_SHIFT_REG & rnode_234to236_bb4_cmp37_i_0_valid_out_0_NO_SHIFT_REG & rnode_235to236_bb4_and193_i_0_valid_out_2_NO_SHIFT_REG & rnode_234to236_bb4_cmp37_i_0_valid_out_1_NO_SHIFT_REG & rnode_235to236_bb4_and195_i_0_valid_out_NO_SHIFT_REG & rnode_235to236_bb4_and193_i_0_valid_out_1_NO_SHIFT_REG & rnode_235to236_bb4_and198_i_0_valid_out_NO_SHIFT_REG & rnode_235to236_bb4_and193_i_0_valid_out_0_NO_SHIFT_REG & rnode_235to236_bb4__and_i_i9_0_valid_out_1_NO_SHIFT_REG & rnode_235to236_bb4__and_i_i9_0_valid_out_2_NO_SHIFT_REG & rnode_235to236_bb4__and_i_i9_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i = (local_bb4__42_i ? (rnode_235to236_bb4_and193_i_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i & 32'h7FFFFFF));
assign local_bb4_and250_i_valid_out = 1'b1;
assign local_bb4_and269_i_valid_out = 1'b1;
assign local_bb4_add245_i_valid_out = 1'b1;
assign local_bb4__45_i_valid_out = 1'b1;
assign local_bb4_not_cmp37_i_valid_out_1 = 1'b1;
assign rnode_234to236_bb4_shr16_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_and17_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_cmp37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_234to236_bb4_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and195_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and198_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4_and193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4__and_i_i9_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4__and_i_i9_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_235to236_bb4__and_i_i9_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or162_i102_stall_local;
wire [31:0] local_bb4_or162_i102;

assign local_bb4_or162_i102 = (local_bb4_or1596_i101 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or1237_i87_stall_local;
wire [7:0] local_bb4_or1237_i87;

assign local_bb4_or1237_i87 = ((local_bb4__30_i81 & 8'h1) | (local_bb4__29_i79 & 8'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__33_i89_stall_local;
wire [7:0] local_bb4__33_i89;

assign local_bb4__33_i89 = (local_bb4_cmp116_i86 ? (local_bb4__29_i79 & 8'h1) : (local_bb4__31_i83 & 8'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_and250_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and250_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_and250_i_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and250_i_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_and250_i_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and250_i_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and250_i_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_and250_i_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_and250_i_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_and250_i_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_and250_i_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_and250_i_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_and250_i_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in((local_bb4_and250_i & 32'hFF)),
	.data_out(rnode_236to237_bb4_and250_i_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_and250_i_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_and250_i_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_236to237_bb4_and250_i_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_and250_i_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_and250_i_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and250_i_stall_in = 1'b0;
assign rnode_236to237_bb4_and250_i_0_NO_SHIFT_REG = rnode_236to237_bb4_and250_i_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_and250_i_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_and250_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_236to238_bb4_and269_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_236to238_bb4_and269_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_236to238_bb4_and269_i_0_NO_SHIFT_REG;
 logic rnode_236to238_bb4_and269_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to238_bb4_and269_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_236to238_bb4_and269_i_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_236to238_bb4_and269_i_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_236to238_bb4_and269_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_236to238_bb4_and269_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to238_bb4_and269_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to238_bb4_and269_i_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_236to238_bb4_and269_i_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_236to238_bb4_and269_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in((local_bb4_and269_i & 32'hFF800000)),
	.data_out(rnode_236to238_bb4_and269_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_236to238_bb4_and269_i_0_reg_238_fifo.DEPTH = 2;
defparam rnode_236to238_bb4_and269_i_0_reg_238_fifo.DATA_WIDTH = 32;
defparam rnode_236to238_bb4_and269_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to238_bb4_and269_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_236to238_bb4_and269_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and269_i_stall_in = 1'b0;
assign rnode_236to238_bb4_and269_i_0_NO_SHIFT_REG = rnode_236to238_bb4_and269_i_0_reg_238_NO_SHIFT_REG;
assign rnode_236to238_bb4_and269_i_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_236to238_bb4_and269_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_add245_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_add245_i_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4_add245_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_add245_i_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4_add245_i_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4_add245_i_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_add245_i_0_valid_out_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_add245_i_0_stall_in_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_add245_i_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_add245_i_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_add245_i_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_add245_i_0_stall_in_0_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_add245_i_0_valid_out_0_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_add245_i_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(local_bb4_add245_i),
	.data_out(rnode_236to237_bb4_add245_i_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_add245_i_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_add245_i_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_236to237_bb4_add245_i_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_add245_i_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_add245_i_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add245_i_stall_in = 1'b0;
assign rnode_236to237_bb4_add245_i_0_stall_in_0_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4_add245_i_0_NO_SHIFT_REG = rnode_236to237_bb4_add245_i_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4_add245_i_1_NO_SHIFT_REG = rnode_236to237_bb4_add245_i_0_reg_237_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4__45_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4__45_i_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4__45_i_1_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4__45_i_2_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_236to237_bb4__45_i_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_valid_out_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_stall_in_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4__45_i_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4__45_i_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4__45_i_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4__45_i_0_stall_in_0_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4__45_i_0_valid_out_0_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4__45_i_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in((local_bb4__45_i & 32'hFFFFFFF)),
	.data_out(rnode_236to237_bb4__45_i_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4__45_i_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4__45_i_0_reg_237_fifo.DATA_WIDTH = 32;
defparam rnode_236to237_bb4__45_i_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4__45_i_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4__45_i_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i_stall_in = 1'b0;
assign rnode_236to237_bb4__45_i_0_stall_in_0_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4__45_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4__45_i_0_NO_SHIFT_REG = rnode_236to237_bb4__45_i_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4__45_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4__45_i_1_NO_SHIFT_REG = rnode_236to237_bb4__45_i_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4__45_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_236to237_bb4__45_i_2_NO_SHIFT_REG = rnode_236to237_bb4__45_i_0_reg_237_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_236to237_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_236to237_bb4_not_cmp37_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_236to237_bb4_not_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_236to237_bb4_not_cmp37_i_0_reg_237_inputs_ready_NO_SHIFT_REG;
 logic rnode_236to237_bb4_not_cmp37_i_0_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_not_cmp37_i_0_valid_out_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_not_cmp37_i_0_stall_in_reg_237_NO_SHIFT_REG;
 logic rnode_236to237_bb4_not_cmp37_i_0_stall_out_reg_237_NO_SHIFT_REG;

acl_data_fifo rnode_236to237_bb4_not_cmp37_i_0_reg_237_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_236to237_bb4_not_cmp37_i_0_reg_237_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_236to237_bb4_not_cmp37_i_0_stall_in_reg_237_NO_SHIFT_REG),
	.valid_out(rnode_236to237_bb4_not_cmp37_i_0_valid_out_reg_237_NO_SHIFT_REG),
	.stall_out(rnode_236to237_bb4_not_cmp37_i_0_stall_out_reg_237_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp37_i),
	.data_out(rnode_236to237_bb4_not_cmp37_i_0_reg_237_NO_SHIFT_REG)
);

defparam rnode_236to237_bb4_not_cmp37_i_0_reg_237_fifo.DEPTH = 1;
defparam rnode_236to237_bb4_not_cmp37_i_0_reg_237_fifo.DATA_WIDTH = 1;
defparam rnode_236to237_bb4_not_cmp37_i_0_reg_237_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_236to237_bb4_not_cmp37_i_0_reg_237_fifo.IMPL = "shift_reg";

assign rnode_236to237_bb4_not_cmp37_i_0_reg_237_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp37_i_stall_in_1 = 1'b0;
assign rnode_236to237_bb4_not_cmp37_i_0_NO_SHIFT_REG = rnode_236to237_bb4_not_cmp37_i_0_reg_237_NO_SHIFT_REG;
assign rnode_236to237_bb4_not_cmp37_i_0_stall_in_reg_237_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__37_v_i103_stall_local;
wire [31:0] local_bb4__37_v_i103;

assign local_bb4__37_v_i103 = (local_bb4_Pivot20_i98 ? 32'h0 : (local_bb4_or162_i102 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or123_i88_stall_local;
wire [31:0] local_bb4_or123_i88;

assign local_bb4_or123_i88[31:8] = 24'h0;
assign local_bb4_or123_i88[7:0] = (local_bb4_or1237_i87 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u88_stall_local;
wire [7:0] local_bb4_var__u88;

assign local_bb4_var__u88 = ((local_bb4__33_i89 & 8'h1) & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i_stall_local;
wire local_bb4_notrhs_i;

assign local_bb4_notrhs_i = ((rnode_236to237_bb4_and250_i_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl273_i_stall_local;
wire [31:0] local_bb4_shl273_i;

assign local_bb4_shl273_i = ((rnode_236to238_bb4_and269_i_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and247_i_stall_local;
wire [31:0] local_bb4_and247_i;

assign local_bb4_and247_i = (rnode_236to237_bb4_add245_i_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp258_i_stall_local;
wire local_bb4_cmp258_i;

assign local_bb4_cmp258_i = ($signed(rnode_236to237_bb4_add245_i_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and225_i_stall_local;
wire [31:0] local_bb4_and225_i;

assign local_bb4_and225_i = ((rnode_236to237_bb4__45_i_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i_stall_local;
wire [31:0] local_bb4_and270_i;

assign local_bb4_and270_i = ((rnode_236to237_bb4__45_i_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr271_i_valid_out;
wire local_bb4_shr271_i_stall_in;
wire local_bb4_shr271_i_inputs_ready;
wire local_bb4_shr271_i_stall_local;
wire [31:0] local_bb4_shr271_i;

assign local_bb4_shr271_i_inputs_ready = rnode_236to237_bb4__45_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr271_i = ((rnode_236to237_bb4__45_i_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr271_i_valid_out = 1'b1;
assign rnode_236to237_bb4__45_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4__39_v_i104_stall_local;
wire [31:0] local_bb4__39_v_i104;

assign local_bb4__39_v_i104 = (local_bb4_SwitchLeaf_i99 ? (local_bb4_var__u85 & 32'h1) : (local_bb4__37_v_i103 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or124_i90_stall_local;
wire [31:0] local_bb4_or124_i90;

assign local_bb4_or124_i90 = (local_bb4_cmp116_i86 ? 32'h0 : (local_bb4_or123_i88 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_conv135_i92_stall_local;
wire [31:0] local_bb4_conv135_i92;

assign local_bb4_conv135_i92[31:8] = 24'h0;
assign local_bb4_conv135_i92[7:0] = (local_bb4_var__u88 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i_stall_local;
wire local_bb4_notlhs_i;

assign local_bb4_notlhs_i = ((local_bb4_and247_i & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_i_stall_local;
wire local_bb4_cmp226_i;

assign local_bb4_cmp226_i = ((local_bb4_and225_i & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i_stall_local;
wire local_bb4_cmp296_i;

assign local_bb4_cmp296_i = ((local_bb4_and270_i & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i_valid_out;
wire local_bb4_cmp296_i_stall_in;
wire local_bb4_cmp299_i_valid_out;
wire local_bb4_cmp299_i_stall_in;
wire local_bb4_cmp299_i_inputs_ready;
wire local_bb4_cmp299_i_stall_local;
wire local_bb4_cmp299_i;

assign local_bb4_cmp299_i_inputs_ready = rnode_236to237_bb4__45_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp299_i = ((local_bb4_and270_i & 32'h7) == 32'h4);
assign local_bb4_cmp296_i_valid_out = 1'b1;
assign local_bb4_cmp299_i_valid_out = 1'b1;
assign rnode_236to237_bb4__45_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_shr271_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_237to238_bb4_shr271_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_shr271_i_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_shr271_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_shr271_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_shr271_i_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_shr271_i_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_shr271_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_shr271_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_shr271_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_shr271_i_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_shr271_i_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_shr271_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in((local_bb4_shr271_i & 32'h1FFFFFF)),
	.data_out(rnode_237to238_bb4_shr271_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_shr271_i_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_shr271_i_0_reg_238_fifo.DATA_WIDTH = 32;
defparam rnode_237to238_bb4_shr271_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_shr271_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_shr271_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr271_i_stall_in = 1'b0;
assign rnode_237to238_bb4_shr271_i_0_NO_SHIFT_REG = rnode_237to238_bb4_shr271_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_shr271_i_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_shr271_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_3_i105_stall_local;
wire [31:0] local_bb4_reduction_3_i105;

assign local_bb4_reduction_3_i105 = ((local_bb4__32_i84 & 32'h1) | (local_bb4_or124_i90 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_or136_i94_stall_local;
wire [31:0] local_bb4_or136_i94;

assign local_bb4_or136_i94 = (local_bb4_cmp131_not_i93 ? (local_bb4_conv135_i92 & 32'h1) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i_stall_local;
wire local_bb4_not__46_i;

assign local_bb4_not__46_i = (local_bb4_notrhs_i | local_bb4_notlhs_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_not_i_stall_local;
wire local_bb4_cmp226_not_i;

assign local_bb4_cmp226_not_i = (local_bb4_cmp226_i ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp296_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp296_i_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp296_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp296_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp296_i_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp296_i_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp296_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_cmp296_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_cmp296_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_cmp296_i_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_cmp296_i_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_cmp296_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(local_bb4_cmp296_i),
	.data_out(rnode_237to238_bb4_cmp296_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_cmp296_i_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_cmp296_i_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_237to238_bb4_cmp296_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_cmp296_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_cmp296_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp296_i_stall_in = 1'b0;
assign rnode_237to238_bb4_cmp296_i_0_NO_SHIFT_REG = rnode_237to238_bb4_cmp296_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_cmp296_i_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp299_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp299_i_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp299_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp299_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp299_i_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp299_i_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_cmp299_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_cmp299_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_cmp299_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_cmp299_i_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_cmp299_i_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_cmp299_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(local_bb4_cmp299_i),
	.data_out(rnode_237to238_bb4_cmp299_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_cmp299_i_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_cmp299_i_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_237to238_bb4_cmp299_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_cmp299_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_cmp299_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp299_i_stall_in = 1'b0;
assign rnode_237to238_bb4_cmp299_i_0_NO_SHIFT_REG = rnode_237to238_bb4_cmp299_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_cmp299_i_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and272_i_stall_local;
wire [31:0] local_bb4_and272_i;

assign local_bb4_and272_i = ((rnode_237to238_bb4_shr271_i_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_5_i107_stall_local;
wire [31:0] local_bb4_reduction_5_i107;

assign local_bb4_reduction_5_i107 = (local_bb4_shr150_i97 | (local_bb4_reduction_3_i105 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_4_i106_stall_local;
wire [31:0] local_bb4_reduction_4_i106;

assign local_bb4_reduction_4_i106 = ((local_bb4_or136_i94 & 32'h1) | (local_bb4__39_v_i104 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4__47_i_stall_local;
wire local_bb4__47_i;

assign local_bb4__47_i = (local_bb4_cmp226_i | local_bb4_not__46_i);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i_stall_local;
wire local_bb4_brmerge12_i;

assign local_bb4_brmerge12_i = (local_bb4_cmp226_not_i | rnode_236to237_bb4_not_cmp37_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot262__i_stall_local;
wire local_bb4_lnot262__i;

assign local_bb4_lnot262__i = (local_bb4_cmp258_i & local_bb4_cmp226_not_i);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29649_i_stall_local;
wire [31:0] local_bb4_cmp29649_i;

assign local_bb4_cmp29649_i[31:1] = 31'h0;
assign local_bb4_cmp29649_i[0] = rnode_237to238_bb4_cmp296_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv300_i_stall_local;
wire [31:0] local_bb4_conv300_i;

assign local_bb4_conv300_i[31:1] = 31'h0;
assign local_bb4_conv300_i[0] = rnode_237to238_bb4_cmp299_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or274_i_stall_local;
wire [31:0] local_bb4_or274_i;

assign local_bb4_or274_i = ((local_bb4_and272_i & 32'h7FFFFF) | (local_bb4_shl273_i & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_6_i108_stall_local;
wire [31:0] local_bb4_reduction_6_i108;

assign local_bb4_reduction_6_i108 = ((local_bb4_reduction_4_i106 & 32'h1) | local_bb4_reduction_5_i107);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i_stall_local;
wire [31:0] local_bb4_resultSign_0_i;

assign local_bb4_resultSign_0_i = (local_bb4_brmerge12_i ? (rnode_236to237_bb4_and35_i_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i_valid_out;
wire local_bb4_resultSign_0_i_stall_in;
wire local_bb4__47_i_valid_out;
wire local_bb4__47_i_stall_in;
wire local_bb4_or2662_i_valid_out;
wire local_bb4_or2662_i_stall_in;
wire local_bb4_or2662_i_inputs_ready;
wire local_bb4_or2662_i_stall_local;
wire local_bb4_or2662_i;

assign local_bb4_or2662_i_inputs_ready = (rnode_236to237_bb4_and35_i_0_valid_out_NO_SHIFT_REG & rnode_236to237_bb4_not_cmp37_i_0_valid_out_NO_SHIFT_REG & rnode_236to237_bb4_add245_i_0_valid_out_0_NO_SHIFT_REG & rnode_236to237_bb4_and250_i_0_valid_out_NO_SHIFT_REG & rnode_236to237_bb4__45_i_0_valid_out_0_NO_SHIFT_REG & rnode_236to237_bb4_add245_i_0_valid_out_1_NO_SHIFT_REG & rnode_236to237_bb4_var__u73_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2662_i = (rnode_236to237_bb4_var__u73_0_NO_SHIFT_REG | local_bb4_lnot262__i);
assign local_bb4_resultSign_0_i_valid_out = 1'b1;
assign local_bb4__47_i_valid_out = 1'b1;
assign local_bb4_or2662_i_valid_out = 1'b1;
assign rnode_236to237_bb4_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_not_cmp37_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_add245_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_and250_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4__45_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_add245_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_236to237_bb4_var__u73_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot33_not_i40_valid_out;
wire local_bb4_lnot33_not_i40_stall_in;
wire local_bb4_cmp37_i36_valid_out;
wire local_bb4_cmp37_i36_stall_in;
wire local_bb4_and36_lobit_i111_valid_out;
wire local_bb4_and36_lobit_i111_stall_in;
wire local_bb4_xor188_i110_valid_out;
wire local_bb4_xor188_i110_stall_in;
wire local_bb4_xor188_i110_inputs_ready;
wire local_bb4_xor188_i110_stall_local;
wire [31:0] local_bb4_xor188_i110;

assign local_bb4_xor188_i110_inputs_ready = (rnode_237to238_bb4__22_i22_0_valid_out_0_NO_SHIFT_REG & rnode_237to238_bb4_lnot23_i31_0_valid_out_NO_SHIFT_REG & rnode_237to238_bb4_align_0_i59_0_valid_out_0_NO_SHIFT_REG & rnode_237to238_bb4_align_0_i59_0_valid_out_4_NO_SHIFT_REG & rnode_237to238_bb4_align_0_i59_0_valid_out_1_NO_SHIFT_REG & rnode_237to238_bb4_align_0_i59_0_valid_out_2_NO_SHIFT_REG & rnode_237to238_bb4_align_0_i59_0_valid_out_3_NO_SHIFT_REG & rnode_237to238_bb4__23_i23_0_valid_out_2_NO_SHIFT_REG & rnode_237to238_bb4__22_i22_0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_xor188_i110 = (local_bb4_reduction_6_i108 ^ local_bb4_xor_lobit_i109);
assign local_bb4_lnot33_not_i40_valid_out = 1'b1;
assign local_bb4_cmp37_i36_valid_out = 1'b1;
assign local_bb4_and36_lobit_i111_valid_out = 1'b1;
assign local_bb4_xor188_i110_valid_out = 1'b1;
assign rnode_237to238_bb4__22_i22_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_lnot23_i31_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_align_0_i59_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_align_0_i59_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_align_0_i59_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_align_0_i59_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_align_0_i59_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__23_i23_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__22_i22_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_237to238_bb4_resultSign_0_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_resultSign_0_i_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_resultSign_0_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_237to238_bb4_resultSign_0_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_resultSign_0_i_0_valid_out_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_resultSign_0_i_0_stall_in_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_resultSign_0_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_resultSign_0_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_resultSign_0_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_resultSign_0_i_0_stall_in_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_resultSign_0_i_0_valid_out_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_resultSign_0_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i & 32'h80000000)),
	.data_out(rnode_237to238_bb4_resultSign_0_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_resultSign_0_i_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_resultSign_0_i_0_reg_238_fifo.DATA_WIDTH = 32;
defparam rnode_237to238_bb4_resultSign_0_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_resultSign_0_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_resultSign_0_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i_stall_in = 1'b0;
assign rnode_237to238_bb4_resultSign_0_i_0_NO_SHIFT_REG = rnode_237to238_bb4_resultSign_0_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_resultSign_0_i_0_stall_in_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4__47_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_valid_out_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_stall_in_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4__47_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4__47_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4__47_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4__47_i_0_stall_in_0_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4__47_i_0_valid_out_0_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4__47_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(local_bb4__47_i),
	.data_out(rnode_237to238_bb4__47_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4__47_i_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4__47_i_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_237to238_bb4__47_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4__47_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4__47_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i_stall_in = 1'b0;
assign rnode_237to238_bb4__47_i_0_stall_in_0_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__47_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__47_i_0_NO_SHIFT_REG = rnode_237to238_bb4__47_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4__47_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4__47_i_1_NO_SHIFT_REG = rnode_237to238_bb4__47_i_0_reg_238_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_237to238_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_1_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_2_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_reg_238_inputs_ready_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_valid_out_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_stall_in_0_reg_238_NO_SHIFT_REG;
 logic rnode_237to238_bb4_or2662_i_0_stall_out_reg_238_NO_SHIFT_REG;

acl_data_fifo rnode_237to238_bb4_or2662_i_0_reg_238_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_237to238_bb4_or2662_i_0_reg_238_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_237to238_bb4_or2662_i_0_stall_in_0_reg_238_NO_SHIFT_REG),
	.valid_out(rnode_237to238_bb4_or2662_i_0_valid_out_0_reg_238_NO_SHIFT_REG),
	.stall_out(rnode_237to238_bb4_or2662_i_0_stall_out_reg_238_NO_SHIFT_REG),
	.data_in(local_bb4_or2662_i),
	.data_out(rnode_237to238_bb4_or2662_i_0_reg_238_NO_SHIFT_REG)
);

defparam rnode_237to238_bb4_or2662_i_0_reg_238_fifo.DEPTH = 1;
defparam rnode_237to238_bb4_or2662_i_0_reg_238_fifo.DATA_WIDTH = 1;
defparam rnode_237to238_bb4_or2662_i_0_reg_238_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_237to238_bb4_or2662_i_0_reg_238_fifo.IMPL = "shift_reg";

assign rnode_237to238_bb4_or2662_i_0_reg_238_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2662_i_stall_in = 1'b0;
assign rnode_237to238_bb4_or2662_i_0_stall_in_0_reg_238_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_or2662_i_0_NO_SHIFT_REG = rnode_237to238_bb4_or2662_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_or2662_i_1_NO_SHIFT_REG = rnode_237to238_bb4_or2662_i_0_reg_238_NO_SHIFT_REG;
assign rnode_237to238_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_237to238_bb4_or2662_i_2_NO_SHIFT_REG = rnode_237to238_bb4_or2662_i_0_reg_238_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_lnot33_not_i40_0_valid_out_NO_SHIFT_REG;
 logic rnode_238to239_bb4_lnot33_not_i40_0_stall_in_NO_SHIFT_REG;
 logic rnode_238to239_bb4_lnot33_not_i40_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_lnot33_not_i40_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic rnode_238to239_bb4_lnot33_not_i40_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_lnot33_not_i40_0_valid_out_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_lnot33_not_i40_0_stall_in_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_lnot33_not_i40_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_lnot33_not_i40_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_lnot33_not_i40_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_lnot33_not_i40_0_stall_in_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_lnot33_not_i40_0_valid_out_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_lnot33_not_i40_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in(local_bb4_lnot33_not_i40),
	.data_out(rnode_238to239_bb4_lnot33_not_i40_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_lnot33_not_i40_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_lnot33_not_i40_0_reg_239_fifo.DATA_WIDTH = 1;
defparam rnode_238to239_bb4_lnot33_not_i40_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_lnot33_not_i40_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_lnot33_not_i40_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_lnot33_not_i40_stall_in = 1'b0;
assign rnode_238to239_bb4_lnot33_not_i40_0_NO_SHIFT_REG = rnode_238to239_bb4_lnot33_not_i40_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_lnot33_not_i40_0_stall_in_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_lnot33_not_i40_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_valid_out_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_stall_in_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_cmp37_i36_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_cmp37_i36_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_cmp37_i36_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_cmp37_i36_0_stall_in_0_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_cmp37_i36_0_valid_out_0_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_cmp37_i36_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in(local_bb4_cmp37_i36),
	.data_out(rnode_238to239_bb4_cmp37_i36_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_cmp37_i36_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_cmp37_i36_0_reg_239_fifo.DATA_WIDTH = 1;
defparam rnode_238to239_bb4_cmp37_i36_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_cmp37_i36_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_cmp37_i36_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp37_i36_stall_in = 1'b0;
assign rnode_238to239_bb4_cmp37_i36_0_stall_in_0_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_cmp37_i36_0_NO_SHIFT_REG = rnode_238to239_bb4_cmp37_i36_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_cmp37_i36_1_NO_SHIFT_REG = rnode_238to239_bb4_cmp37_i36_0_reg_239_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_and36_lobit_i111_0_valid_out_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and36_lobit_i111_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_and36_lobit_i111_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and36_lobit_i111_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_and36_lobit_i111_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and36_lobit_i111_0_valid_out_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and36_lobit_i111_0_stall_in_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_and36_lobit_i111_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_and36_lobit_i111_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_and36_lobit_i111_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_and36_lobit_i111_0_stall_in_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_and36_lobit_i111_0_valid_out_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_and36_lobit_i111_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in((local_bb4_and36_lobit_i111 & 32'h1)),
	.data_out(rnode_238to239_bb4_and36_lobit_i111_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_and36_lobit_i111_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_and36_lobit_i111_0_reg_239_fifo.DATA_WIDTH = 32;
defparam rnode_238to239_bb4_and36_lobit_i111_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_and36_lobit_i111_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_and36_lobit_i111_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and36_lobit_i111_stall_in = 1'b0;
assign rnode_238to239_bb4_and36_lobit_i111_0_NO_SHIFT_REG = rnode_238to239_bb4_and36_lobit_i111_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_and36_lobit_i111_0_stall_in_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_and36_lobit_i111_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4_xor188_i110_0_valid_out_NO_SHIFT_REG;
 logic rnode_238to239_bb4_xor188_i110_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_xor188_i110_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4_xor188_i110_0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4_xor188_i110_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_xor188_i110_0_valid_out_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_xor188_i110_0_stall_in_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4_xor188_i110_0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4_xor188_i110_0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4_xor188_i110_0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4_xor188_i110_0_stall_in_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4_xor188_i110_0_valid_out_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4_xor188_i110_0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in(local_bb4_xor188_i110),
	.data_out(rnode_238to239_bb4_xor188_i110_0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4_xor188_i110_0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4_xor188_i110_0_reg_239_fifo.DATA_WIDTH = 32;
defparam rnode_238to239_bb4_xor188_i110_0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4_xor188_i110_0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4_xor188_i110_0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_xor188_i110_stall_in = 1'b0;
assign rnode_238to239_bb4_xor188_i110_0_NO_SHIFT_REG = rnode_238to239_bb4_xor188_i110_0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4_xor188_i110_0_stall_in_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_xor188_i110_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i_stall_local;
wire [31:0] local_bb4_or275_i;

assign local_bb4_or275_i = ((local_bb4_or274_i & 32'h7FFFFFFF) | (rnode_237to238_bb4_resultSign_0_i_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u89_stall_local;
wire [31:0] local_bb4_var__u89;

assign local_bb4_var__u89[31:1] = 31'h0;
assign local_bb4_var__u89[0] = rnode_237to238_bb4__47_i_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2804_i_stall_local;
wire local_bb4_or2804_i;

assign local_bb4_or2804_i = (rnode_237to238_bb4__47_i_0_NO_SHIFT_REG | rnode_237to238_bb4_or2662_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2875_i_stall_local;
wire local_bb4_or2875_i;

assign local_bb4_or2875_i = (rnode_237to238_bb4_or2662_i_1_NO_SHIFT_REG | rnode_237to238_bb4__26_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u90_stall_local;
wire [31:0] local_bb4_var__u90;

assign local_bb4_var__u90[31:1] = 31'h0;
assign local_bb4_var__u90[0] = rnode_237to238_bb4_or2662_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_i41_stall_local;
wire local_bb4_brmerge_not_i41;

assign local_bb4_brmerge_not_i41 = (rnode_237to239_bb4_cmp27_i33_0_NO_SHIFT_REG & rnode_238to239_bb4_lnot33_not_i40_0_NO_SHIFT_REG);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_239to241_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_1_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_2_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_valid_out_0_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_stall_in_0_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_cmp37_i36_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_239to241_bb4_cmp37_i36_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to241_bb4_cmp37_i36_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to241_bb4_cmp37_i36_0_stall_in_0_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_239to241_bb4_cmp37_i36_0_valid_out_0_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_239to241_bb4_cmp37_i36_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in(rnode_238to239_bb4_cmp37_i36_1_NO_SHIFT_REG),
	.data_out(rnode_239to241_bb4_cmp37_i36_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_239to241_bb4_cmp37_i36_0_reg_241_fifo.DEPTH = 2;
defparam rnode_239to241_bb4_cmp37_i36_0_reg_241_fifo.DATA_WIDTH = 1;
defparam rnode_239to241_bb4_cmp37_i36_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to241_bb4_cmp37_i36_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_239to241_bb4_cmp37_i36_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_cmp37_i36_0_stall_in_0_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_239to241_bb4_cmp37_i36_0_NO_SHIFT_REG = rnode_239to241_bb4_cmp37_i36_0_reg_241_NO_SHIFT_REG;
assign rnode_239to241_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_239to241_bb4_cmp37_i36_1_NO_SHIFT_REG = rnode_239to241_bb4_cmp37_i36_0_reg_241_NO_SHIFT_REG;
assign rnode_239to241_bb4_cmp37_i36_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_239to241_bb4_cmp37_i36_2_NO_SHIFT_REG = rnode_239to241_bb4_cmp37_i36_0_reg_241_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_add_i112_stall_local;
wire [31:0] local_bb4_add_i112;

assign local_bb4_add_i112 = ((local_bb4__27_i52 & 32'h7FFFFF8) | (rnode_238to239_bb4_and36_lobit_i111_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext314_i_stall_local;
wire [31:0] local_bb4_lnot_ext314_i;

assign local_bb4_lnot_ext314_i = ((local_bb4_var__u89 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond282_i_stall_local;
wire [31:0] local_bb4_cond282_i;

assign local_bb4_cond282_i = (local_bb4_or2804_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond289_i_stall_local;
wire [31:0] local_bb4_cond289_i;

assign local_bb4_cond289_i = (local_bb4_or2875_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext310_i_stall_local;
wire [31:0] local_bb4_lnot_ext310_i;

assign local_bb4_lnot_ext310_i = ((local_bb4_var__u90 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__24_i44_stall_local;
wire local_bb4__24_i44;

assign local_bb4__24_i44 = (local_bb4_or_cond_not_i43 | local_bb4_brmerge_not_i41);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge_not_not_i45_stall_local;
wire local_bb4_brmerge_not_not_i45;

assign local_bb4_brmerge_not_not_i45 = (local_bb4_brmerge_not_i41 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_not_cmp37_i142_stall_local;
wire local_bb4_not_cmp37_i142;

assign local_bb4_not_cmp37_i142 = (rnode_239to241_bb4_cmp37_i36_1_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb4_add192_i113_stall_local;
wire [31:0] local_bb4_add192_i113;

assign local_bb4_add192_i113 = ((local_bb4_add_i112 & 32'h7FFFFF9) + rnode_238to239_bb4_xor188_i110_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_and293_i_stall_local;
wire [31:0] local_bb4_and293_i;

assign local_bb4_and293_i = ((local_bb4_cond282_i | 32'h80000000) & local_bb4_or275_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or294_i_stall_local;
wire [31:0] local_bb4_or294_i;

assign local_bb4_or294_i = ((local_bb4_cond289_i & 32'h7F800000) | (local_bb4_cond292_i & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i_stall_local;
wire [31:0] local_bb4_reduction_0_i;

assign local_bb4_reduction_0_i = ((local_bb4_lnot_ext310_i & 32'h1) & (local_bb4_lnot_ext_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_7_i46_stall_local;
wire local_bb4_reduction_7_i46;

assign local_bb4_reduction_7_i46 = (local_bb4_cmp25_i32 & local_bb4_brmerge_not_not_i45);

// This section implements an unregistered operation.
// 
wire local_bb4_and302_i_stall_local;
wire [31:0] local_bb4_and302_i;

assign local_bb4_and302_i = ((local_bb4_conv300_i & 32'h1) & local_bb4_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i_stall_local;
wire [31:0] local_bb4_or295_i;

assign local_bb4_or295_i = ((local_bb4_or294_i & 32'h7FC00000) | local_bb4_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_9_i48_stall_local;
wire local_bb4_reduction_9_i48;

assign local_bb4_reduction_9_i48 = (local_bb4_reduction_7_i46 & local_bb4_reduction_8_i47);

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i_stall_local;
wire [31:0] local_bb4_lor_ext_i;

assign local_bb4_lor_ext_i = ((local_bb4_cmp29649_i & 32'h1) | (local_bb4_and302_i & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and17_i25_valid_out_2;
wire local_bb4_and17_i25_stall_in_2;
wire local_bb4_var__u83_valid_out;
wire local_bb4_var__u83_stall_in;
wire local_bb4_add192_i113_valid_out;
wire local_bb4_add192_i113_stall_in;
wire local_bb4__26_i49_valid_out;
wire local_bb4__26_i49_stall_in;
wire local_bb4__26_i49_inputs_ready;
wire local_bb4__26_i49_stall_local;
wire local_bb4__26_i49;

assign local_bb4__26_i49_inputs_ready = (rnode_237to239_bb4_shr16_i24_0_valid_out_0_NO_SHIFT_REG & rnode_237to239_bb4_cmp27_i33_0_valid_out_2_NO_SHIFT_REG & rnode_238to239_bb4_and36_lobit_i111_0_valid_out_NO_SHIFT_REG & rnode_238to239_bb4_xor188_i110_0_valid_out_NO_SHIFT_REG & rnode_238to239_bb4_and20_i28_0_valid_out_0_NO_SHIFT_REG & rnode_237to239_bb4_cmp27_i33_0_valid_out_0_NO_SHIFT_REG & rnode_238to239_bb4_lnot33_not_i40_0_valid_out_NO_SHIFT_REG & rnode_237to239_bb4_cmp27_i33_0_valid_out_1_NO_SHIFT_REG & rnode_238to239_bb4_and20_i28_0_valid_out_1_NO_SHIFT_REG & rnode_238to239_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__26_i49 = (local_bb4_reduction_9_i48 ? rnode_238to239_bb4_cmp37_i36_0_NO_SHIFT_REG : local_bb4__24_i44);
assign local_bb4_and17_i25_valid_out_2 = 1'b1;
assign local_bb4_var__u83_valid_out = 1'b1;
assign local_bb4_add192_i113_valid_out = 1'b1;
assign local_bb4__26_i49_valid_out = 1'b1;
assign rnode_237to239_bb4_shr16_i24_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to239_bb4_cmp27_i33_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_and36_lobit_i111_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_xor188_i110_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_and20_i28_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to239_bb4_cmp27_i33_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_lnot33_not_i40_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to239_bb4_cmp27_i33_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_and20_i28_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i_stall_local;
wire [31:0] local_bb4_reduction_1_i;

assign local_bb4_reduction_1_i = ((local_bb4_lnot_ext314_i & 32'h1) & (local_bb4_lor_ext_i & 32'h1));

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_239to241_bb4_and17_i25_0_valid_out_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and17_i25_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_239to241_bb4_and17_i25_0_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and17_i25_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_239to241_bb4_and17_i25_0_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and17_i25_0_valid_out_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and17_i25_0_stall_in_reg_241_NO_SHIFT_REG;
 logic rnode_239to241_bb4_and17_i25_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_239to241_bb4_and17_i25_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to241_bb4_and17_i25_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to241_bb4_and17_i25_0_stall_in_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_239to241_bb4_and17_i25_0_valid_out_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_239to241_bb4_and17_i25_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in((local_bb4_and17_i25 & 32'hFF)),
	.data_out(rnode_239to241_bb4_and17_i25_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_239to241_bb4_and17_i25_0_reg_241_fifo.DEPTH = 2;
defparam rnode_239to241_bb4_and17_i25_0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_239to241_bb4_and17_i25_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to241_bb4_and17_i25_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_239to241_bb4_and17_i25_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and17_i25_stall_in_2 = 1'b0;
assign rnode_239to241_bb4_and17_i25_0_NO_SHIFT_REG = rnode_239to241_bb4_and17_i25_0_reg_241_NO_SHIFT_REG;
assign rnode_239to241_bb4_and17_i25_0_stall_in_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_and17_i25_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_239to240_bb4_var__u83_0_valid_out_NO_SHIFT_REG;
 logic rnode_239to240_bb4_var__u83_0_stall_in_NO_SHIFT_REG;
 logic rnode_239to240_bb4_var__u83_0_NO_SHIFT_REG;
 logic rnode_239to240_bb4_var__u83_0_reg_240_inputs_ready_NO_SHIFT_REG;
 logic rnode_239to240_bb4_var__u83_0_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_var__u83_0_valid_out_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_var__u83_0_stall_in_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_var__u83_0_stall_out_reg_240_NO_SHIFT_REG;

acl_data_fifo rnode_239to240_bb4_var__u83_0_reg_240_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to240_bb4_var__u83_0_reg_240_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to240_bb4_var__u83_0_stall_in_reg_240_NO_SHIFT_REG),
	.valid_out(rnode_239to240_bb4_var__u83_0_valid_out_reg_240_NO_SHIFT_REG),
	.stall_out(rnode_239to240_bb4_var__u83_0_stall_out_reg_240_NO_SHIFT_REG),
	.data_in(local_bb4_var__u83),
	.data_out(rnode_239to240_bb4_var__u83_0_reg_240_NO_SHIFT_REG)
);

defparam rnode_239to240_bb4_var__u83_0_reg_240_fifo.DEPTH = 1;
defparam rnode_239to240_bb4_var__u83_0_reg_240_fifo.DATA_WIDTH = 1;
defparam rnode_239to240_bb4_var__u83_0_reg_240_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to240_bb4_var__u83_0_reg_240_fifo.IMPL = "shift_reg";

assign rnode_239to240_bb4_var__u83_0_reg_240_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_var__u83_stall_in = 1'b0;
assign rnode_239to240_bb4_var__u83_0_NO_SHIFT_REG = rnode_239to240_bb4_var__u83_0_reg_240_NO_SHIFT_REG;
assign rnode_239to240_bb4_var__u83_0_stall_in_reg_240_NO_SHIFT_REG = 1'b0;
assign rnode_239to240_bb4_var__u83_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_239to240_bb4_add192_i113_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_239to240_bb4_add192_i113_0_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_239to240_bb4_add192_i113_1_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_239to240_bb4_add192_i113_2_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_239to240_bb4_add192_i113_3_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_reg_240_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_239to240_bb4_add192_i113_0_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_valid_out_0_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_stall_in_0_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4_add192_i113_0_stall_out_reg_240_NO_SHIFT_REG;

acl_data_fifo rnode_239to240_bb4_add192_i113_0_reg_240_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to240_bb4_add192_i113_0_reg_240_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to240_bb4_add192_i113_0_stall_in_0_reg_240_NO_SHIFT_REG),
	.valid_out(rnode_239to240_bb4_add192_i113_0_valid_out_0_reg_240_NO_SHIFT_REG),
	.stall_out(rnode_239to240_bb4_add192_i113_0_stall_out_reg_240_NO_SHIFT_REG),
	.data_in(local_bb4_add192_i113),
	.data_out(rnode_239to240_bb4_add192_i113_0_reg_240_NO_SHIFT_REG)
);

defparam rnode_239to240_bb4_add192_i113_0_reg_240_fifo.DEPTH = 1;
defparam rnode_239to240_bb4_add192_i113_0_reg_240_fifo.DATA_WIDTH = 32;
defparam rnode_239to240_bb4_add192_i113_0_reg_240_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to240_bb4_add192_i113_0_reg_240_fifo.IMPL = "shift_reg";

assign rnode_239to240_bb4_add192_i113_0_reg_240_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add192_i113_stall_in = 1'b0;
assign rnode_239to240_bb4_add192_i113_0_stall_in_0_reg_240_NO_SHIFT_REG = 1'b0;
assign rnode_239to240_bb4_add192_i113_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4_add192_i113_0_NO_SHIFT_REG = rnode_239to240_bb4_add192_i113_0_reg_240_NO_SHIFT_REG;
assign rnode_239to240_bb4_add192_i113_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4_add192_i113_1_NO_SHIFT_REG = rnode_239to240_bb4_add192_i113_0_reg_240_NO_SHIFT_REG;
assign rnode_239to240_bb4_add192_i113_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4_add192_i113_2_NO_SHIFT_REG = rnode_239to240_bb4_add192_i113_0_reg_240_NO_SHIFT_REG;
assign rnode_239to240_bb4_add192_i113_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4_add192_i113_3_NO_SHIFT_REG = rnode_239to240_bb4_add192_i113_0_reg_240_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_239to240_bb4__26_i49_0_valid_out_NO_SHIFT_REG;
 logic rnode_239to240_bb4__26_i49_0_stall_in_NO_SHIFT_REG;
 logic rnode_239to240_bb4__26_i49_0_NO_SHIFT_REG;
 logic rnode_239to240_bb4__26_i49_0_reg_240_inputs_ready_NO_SHIFT_REG;
 logic rnode_239to240_bb4__26_i49_0_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4__26_i49_0_valid_out_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4__26_i49_0_stall_in_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4__26_i49_0_stall_out_reg_240_NO_SHIFT_REG;

acl_data_fifo rnode_239to240_bb4__26_i49_0_reg_240_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to240_bb4__26_i49_0_reg_240_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to240_bb4__26_i49_0_stall_in_reg_240_NO_SHIFT_REG),
	.valid_out(rnode_239to240_bb4__26_i49_0_valid_out_reg_240_NO_SHIFT_REG),
	.stall_out(rnode_239to240_bb4__26_i49_0_stall_out_reg_240_NO_SHIFT_REG),
	.data_in(local_bb4__26_i49),
	.data_out(rnode_239to240_bb4__26_i49_0_reg_240_NO_SHIFT_REG)
);

defparam rnode_239to240_bb4__26_i49_0_reg_240_fifo.DEPTH = 1;
defparam rnode_239to240_bb4__26_i49_0_reg_240_fifo.DATA_WIDTH = 1;
defparam rnode_239to240_bb4__26_i49_0_reg_240_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to240_bb4__26_i49_0_reg_240_fifo.IMPL = "shift_reg";

assign rnode_239to240_bb4__26_i49_0_reg_240_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__26_i49_stall_in = 1'b0;
assign rnode_239to240_bb4__26_i49_0_NO_SHIFT_REG = rnode_239to240_bb4__26_i49_0_reg_240_NO_SHIFT_REG;
assign rnode_239to240_bb4__26_i49_0_stall_in_reg_240_NO_SHIFT_REG = 1'b0;
assign rnode_239to240_bb4__26_i49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i_stall_local;
wire [31:0] local_bb4_reduction_2_i;

assign local_bb4_reduction_2_i = ((local_bb4_reduction_0_i & 32'h1) & (local_bb4_reduction_1_i & 32'h1));

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_240to241_bb4_var__u83_0_valid_out_NO_SHIFT_REG;
 logic rnode_240to241_bb4_var__u83_0_stall_in_NO_SHIFT_REG;
 logic rnode_240to241_bb4_var__u83_0_NO_SHIFT_REG;
 logic rnode_240to241_bb4_var__u83_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic rnode_240to241_bb4_var__u83_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_var__u83_0_valid_out_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_var__u83_0_stall_in_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_var__u83_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_240to241_bb4_var__u83_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to241_bb4_var__u83_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to241_bb4_var__u83_0_stall_in_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_240to241_bb4_var__u83_0_valid_out_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_240to241_bb4_var__u83_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in(rnode_239to240_bb4_var__u83_0_NO_SHIFT_REG),
	.data_out(rnode_240to241_bb4_var__u83_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_240to241_bb4_var__u83_0_reg_241_fifo.DEPTH = 1;
defparam rnode_240to241_bb4_var__u83_0_reg_241_fifo.DATA_WIDTH = 1;
defparam rnode_240to241_bb4_var__u83_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to241_bb4_var__u83_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_240to241_bb4_var__u83_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4_var__u83_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_var__u83_0_NO_SHIFT_REG = rnode_240to241_bb4_var__u83_0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4_var__u83_0_stall_in_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_var__u83_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and193_i114_valid_out;
wire local_bb4_and193_i114_stall_in;
wire local_bb4_and193_i114_inputs_ready;
wire local_bb4_and193_i114_stall_local;
wire [31:0] local_bb4_and193_i114;

assign local_bb4_and193_i114_inputs_ready = rnode_239to240_bb4_add192_i113_0_valid_out_0_NO_SHIFT_REG;
assign local_bb4_and193_i114 = (rnode_239to240_bb4_add192_i113_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb4_and193_i114_valid_out = 1'b1;
assign rnode_239to240_bb4_add192_i113_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and195_i115_valid_out;
wire local_bb4_and195_i115_stall_in;
wire local_bb4_and195_i115_inputs_ready;
wire local_bb4_and195_i115_stall_local;
wire [31:0] local_bb4_and195_i115;

assign local_bb4_and195_i115_inputs_ready = rnode_239to240_bb4_add192_i113_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_and195_i115 = (rnode_239to240_bb4_add192_i113_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb4_and195_i115_valid_out = 1'b1;
assign rnode_239to240_bb4_add192_i113_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and198_i116_valid_out;
wire local_bb4_and198_i116_stall_in;
wire local_bb4_and198_i116_inputs_ready;
wire local_bb4_and198_i116_stall_local;
wire [31:0] local_bb4_and198_i116;

assign local_bb4_and198_i116_inputs_ready = rnode_239to240_bb4_add192_i113_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_and198_i116 = (rnode_239to240_bb4_add192_i113_2_NO_SHIFT_REG & 32'h1);
assign local_bb4_and198_i116_valid_out = 1'b1;
assign rnode_239to240_bb4_add192_i113_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_and201_i117_stall_local;
wire [31:0] local_bb4_and201_i117;

assign local_bb4_and201_i117 = (rnode_239to240_bb4_add192_i113_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_240to242_bb4__26_i49_0_valid_out_NO_SHIFT_REG;
 logic rnode_240to242_bb4__26_i49_0_stall_in_NO_SHIFT_REG;
 logic rnode_240to242_bb4__26_i49_0_NO_SHIFT_REG;
 logic rnode_240to242_bb4__26_i49_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic rnode_240to242_bb4__26_i49_0_reg_242_NO_SHIFT_REG;
 logic rnode_240to242_bb4__26_i49_0_valid_out_reg_242_NO_SHIFT_REG;
 logic rnode_240to242_bb4__26_i49_0_stall_in_reg_242_NO_SHIFT_REG;
 logic rnode_240to242_bb4__26_i49_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_240to242_bb4__26_i49_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to242_bb4__26_i49_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to242_bb4__26_i49_0_stall_in_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_240to242_bb4__26_i49_0_valid_out_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_240to242_bb4__26_i49_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in(rnode_239to240_bb4__26_i49_0_NO_SHIFT_REG),
	.data_out(rnode_240to242_bb4__26_i49_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_240to242_bb4__26_i49_0_reg_242_fifo.DEPTH = 2;
defparam rnode_240to242_bb4__26_i49_0_reg_242_fifo.DATA_WIDTH = 1;
defparam rnode_240to242_bb4__26_i49_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to242_bb4__26_i49_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_240to242_bb4__26_i49_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4__26_i49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_240to242_bb4__26_i49_0_NO_SHIFT_REG = rnode_240to242_bb4__26_i49_0_reg_242_NO_SHIFT_REG;
assign rnode_240to242_bb4__26_i49_0_stall_in_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_240to242_bb4__26_i49_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_add320_i_stall_local;
wire [31:0] local_bb4_add320_i;

assign local_bb4_add320_i = ((local_bb4_reduction_2_i & 32'h1) + local_bb4_or295_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_241to242_bb4_var__u83_0_valid_out_NO_SHIFT_REG;
 logic rnode_241to242_bb4_var__u83_0_stall_in_NO_SHIFT_REG;
 logic rnode_241to242_bb4_var__u83_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4_var__u83_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic rnode_241to242_bb4_var__u83_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_var__u83_0_valid_out_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_var__u83_0_stall_in_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_var__u83_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_241to242_bb4_var__u83_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to242_bb4_var__u83_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to242_bb4_var__u83_0_stall_in_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_241to242_bb4_var__u83_0_valid_out_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_241to242_bb4_var__u83_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in(rnode_240to241_bb4_var__u83_0_NO_SHIFT_REG),
	.data_out(rnode_241to242_bb4_var__u83_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_241to242_bb4_var__u83_0_reg_242_fifo.DEPTH = 1;
defparam rnode_241to242_bb4_var__u83_0_reg_242_fifo.DATA_WIDTH = 1;
defparam rnode_241to242_bb4_var__u83_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to242_bb4_var__u83_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_241to242_bb4_var__u83_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4_var__u83_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_var__u83_0_NO_SHIFT_REG = rnode_241to242_bb4_var__u83_0_reg_242_NO_SHIFT_REG;
assign rnode_241to242_bb4_var__u83_0_stall_in_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_var__u83_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_240to241_bb4_and193_i114_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and193_i114_0_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and193_i114_1_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and193_i114_2_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and193_i114_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_valid_out_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_stall_in_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and193_i114_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_240to241_bb4_and193_i114_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to241_bb4_and193_i114_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to241_bb4_and193_i114_0_stall_in_0_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_240to241_bb4_and193_i114_0_valid_out_0_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_240to241_bb4_and193_i114_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in((local_bb4_and193_i114 & 32'hFFFFFFF)),
	.data_out(rnode_240to241_bb4_and193_i114_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_240to241_bb4_and193_i114_0_reg_241_fifo.DEPTH = 1;
defparam rnode_240to241_bb4_and193_i114_0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_240to241_bb4_and193_i114_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to241_bb4_and193_i114_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_240to241_bb4_and193_i114_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and193_i114_stall_in = 1'b0;
assign rnode_240to241_bb4_and193_i114_0_stall_in_0_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and193_i114_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4_and193_i114_0_NO_SHIFT_REG = rnode_240to241_bb4_and193_i114_0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4_and193_i114_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4_and193_i114_1_NO_SHIFT_REG = rnode_240to241_bb4_and193_i114_0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4_and193_i114_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4_and193_i114_2_NO_SHIFT_REG = rnode_240to241_bb4_and193_i114_0_reg_241_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_240to241_bb4_and195_i115_0_valid_out_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and195_i115_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and195_i115_0_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and195_i115_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and195_i115_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and195_i115_0_valid_out_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and195_i115_0_stall_in_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and195_i115_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_240to241_bb4_and195_i115_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to241_bb4_and195_i115_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to241_bb4_and195_i115_0_stall_in_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_240to241_bb4_and195_i115_0_valid_out_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_240to241_bb4_and195_i115_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in((local_bb4_and195_i115 & 32'h1F)),
	.data_out(rnode_240to241_bb4_and195_i115_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_240to241_bb4_and195_i115_0_reg_241_fifo.DEPTH = 1;
defparam rnode_240to241_bb4_and195_i115_0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_240to241_bb4_and195_i115_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to241_bb4_and195_i115_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_240to241_bb4_and195_i115_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and195_i115_stall_in = 1'b0;
assign rnode_240to241_bb4_and195_i115_0_NO_SHIFT_REG = rnode_240to241_bb4_and195_i115_0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4_and195_i115_0_stall_in_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and195_i115_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_240to241_bb4_and198_i116_0_valid_out_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and198_i116_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and198_i116_0_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and198_i116_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_and198_i116_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and198_i116_0_valid_out_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and198_i116_0_stall_in_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_and198_i116_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_240to241_bb4_and198_i116_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to241_bb4_and198_i116_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to241_bb4_and198_i116_0_stall_in_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_240to241_bb4_and198_i116_0_valid_out_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_240to241_bb4_and198_i116_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in((local_bb4_and198_i116 & 32'h1)),
	.data_out(rnode_240to241_bb4_and198_i116_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_240to241_bb4_and198_i116_0_reg_241_fifo.DEPTH = 1;
defparam rnode_240to241_bb4_and198_i116_0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_240to241_bb4_and198_i116_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to241_bb4_and198_i116_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_240to241_bb4_and198_i116_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and198_i116_stall_in = 1'b0;
assign rnode_240to241_bb4_and198_i116_0_NO_SHIFT_REG = rnode_240to241_bb4_and198_i116_0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4_and198_i116_0_stall_in_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and198_i116_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_shr_i_i118_stall_local;
wire [31:0] local_bb4_shr_i_i118;

assign local_bb4_shr_i_i118 = ((local_bb4_and201_i117 & 32'h7FFFFFF) >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4__26_i49_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_2_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_valid_out_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_stall_in_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4__26_i49_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4__26_i49_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4__26_i49_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4__26_i49_0_stall_in_0_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4__26_i49_0_valid_out_0_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4__26_i49_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(rnode_240to242_bb4__26_i49_0_NO_SHIFT_REG),
	.data_out(rnode_242to243_bb4__26_i49_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4__26_i49_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4__26_i49_0_reg_243_fifo.DATA_WIDTH = 1;
defparam rnode_242to243_bb4__26_i49_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4__26_i49_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4__26_i49_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_240to242_bb4__26_i49_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__26_i49_0_stall_in_0_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__26_i49_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4__26_i49_0_NO_SHIFT_REG = rnode_242to243_bb4__26_i49_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4__26_i49_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4__26_i49_1_NO_SHIFT_REG = rnode_242to243_bb4__26_i49_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4__26_i49_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4__26_i49_2_NO_SHIFT_REG = rnode_242to243_bb4__26_i49_0_reg_243_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_var__u91_stall_local;
wire [31:0] local_bb4_var__u91;

assign local_bb4_var__u91 = local_bb4_add320_i;

// This section implements an unregistered operation.
// 
wire local_bb4_shr216_i139_stall_local;
wire [31:0] local_bb4_shr216_i139;

assign local_bb4_shr216_i139 = ((rnode_240to241_bb4_and193_i114_1_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4__pre_i137_stall_local;
wire [31:0] local_bb4__pre_i137;

assign local_bb4__pre_i137 = ((rnode_240to241_bb4_and195_i115_0_NO_SHIFT_REG & 32'h1F) & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_or_i_i119_stall_local;
wire [31:0] local_bb4_or_i_i119;

assign local_bb4_or_i_i119 = ((local_bb4_shr_i_i118 & 32'h3FFFFFF) | (local_bb4_and201_i117 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_cond292_i176_stall_local;
wire [31:0] local_bb4_cond292_i176;

assign local_bb4_cond292_i176 = (rnode_242to243_bb4__26_i49_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u92_stall_local;
wire [31:0] local_bb4_var__u92;

assign local_bb4_var__u92[31:1] = 31'h0;
assign local_bb4_var__u92[0] = rnode_242to243_bb4__26_i49_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4___valid_out;
wire local_bb4___stall_in;
wire local_bb4___inputs_ready;
wire local_bb4___stall_local;
wire [31:0] local_bb4__;

assign local_bb4___inputs_ready = (rnode_237to238_bb4_cmp34_0_valid_out_0_NO_SHIFT_REG & rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_valid_out_NO_SHIFT_REG & rnode_236to238_bb4_and269_i_0_valid_out_NO_SHIFT_REG & rnode_237to238_bb4_resultSign_0_i_0_valid_out_NO_SHIFT_REG & rnode_237to238_bb4_or2662_i_0_valid_out_1_NO_SHIFT_REG & rnode_237to238_bb4__26_i_0_valid_out_0_NO_SHIFT_REG & rnode_237to238_bb4__26_i_0_valid_out_1_NO_SHIFT_REG & rnode_237to238_bb4__47_i_0_valid_out_0_NO_SHIFT_REG & rnode_237to238_bb4_or2662_i_0_valid_out_0_NO_SHIFT_REG & rnode_237to238_bb4__26_i_0_valid_out_2_NO_SHIFT_REG & rnode_237to238_bb4_or2662_i_0_valid_out_2_NO_SHIFT_REG & rnode_237to238_bb4_shr271_i_0_valid_out_NO_SHIFT_REG & rnode_237to238_bb4__47_i_0_valid_out_1_NO_SHIFT_REG & rnode_237to238_bb4_cmp296_i_0_valid_out_NO_SHIFT_REG & rnode_237to238_bb4_cmp299_i_0_valid_out_NO_SHIFT_REG);
assign local_bb4__ = (rnode_237to238_bb4_cmp34_0_NO_SHIFT_REG ? local_bb4_var__u91 : rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_NO_SHIFT_REG);
assign local_bb4___valid_out = 1'b1;
assign rnode_237to238_bb4_cmp34_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_sum_321_pop9_c1_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_236to238_bb4_and269_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_resultSign_0_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_or2662_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__26_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__26_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__47_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_or2662_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__26_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_or2662_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_shr271_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4__47_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_cmp296_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_237to238_bb4_cmp299_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_or219_i140_stall_local;
wire [31:0] local_bb4_or219_i140;

assign local_bb4_or219_i140 = ((local_bb4_shr216_i139 & 32'h7FFFFFF) | (rnode_240to241_bb4_and198_i116_0_NO_SHIFT_REG & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_tobool213_i138_stall_local;
wire local_bb4_tobool213_i138;

assign local_bb4_tobool213_i138 = ((local_bb4__pre_i137 & 32'h1) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shr1_i_i120_stall_local;
wire [31:0] local_bb4_shr1_i_i120;

assign local_bb4_shr1_i_i120 = ((local_bb4_or_i_i119 & 32'h7FFFFFF) >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext_i186_stall_local;
wire [31:0] local_bb4_lnot_ext_i186;

assign local_bb4_lnot_ext_i186 = ((local_bb4_var__u92 & 32'h1) ^ 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_238to239_bb4___0_valid_out_0_NO_SHIFT_REG;
 logic rnode_238to239_bb4___0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4___0_NO_SHIFT_REG;
 logic rnode_238to239_bb4___0_valid_out_1_NO_SHIFT_REG;
 logic rnode_238to239_bb4___0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4___1_NO_SHIFT_REG;
 logic rnode_238to239_bb4___0_reg_239_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_238to239_bb4___0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4___0_valid_out_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4___0_stall_in_0_reg_239_NO_SHIFT_REG;
 logic rnode_238to239_bb4___0_stall_out_reg_239_NO_SHIFT_REG;

acl_data_fifo rnode_238to239_bb4___0_reg_239_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_238to239_bb4___0_reg_239_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_238to239_bb4___0_stall_in_0_reg_239_NO_SHIFT_REG),
	.valid_out(rnode_238to239_bb4___0_valid_out_0_reg_239_NO_SHIFT_REG),
	.stall_out(rnode_238to239_bb4___0_stall_out_reg_239_NO_SHIFT_REG),
	.data_in(local_bb4__),
	.data_out(rnode_238to239_bb4___0_reg_239_NO_SHIFT_REG)
);

defparam rnode_238to239_bb4___0_reg_239_fifo.DEPTH = 1;
defparam rnode_238to239_bb4___0_reg_239_fifo.DATA_WIDTH = 32;
defparam rnode_238to239_bb4___0_reg_239_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_238to239_bb4___0_reg_239_fifo.IMPL = "shift_reg";

assign rnode_238to239_bb4___0_reg_239_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4___stall_in = 1'b0;
assign rnode_238to239_bb4___0_stall_in_0_reg_239_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4___0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4___0_NO_SHIFT_REG = rnode_238to239_bb4___0_reg_239_NO_SHIFT_REG;
assign rnode_238to239_bb4___0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4___1_NO_SHIFT_REG = rnode_238to239_bb4___0_reg_239_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4__40_demorgan_i141_stall_local;
wire local_bb4__40_demorgan_i141;

assign local_bb4__40_demorgan_i141 = (rnode_239to241_bb4_cmp37_i36_0_NO_SHIFT_REG | local_bb4_tobool213_i138);

// This section implements an unregistered operation.
// 
wire local_bb4__42_i143_stall_local;
wire local_bb4__42_i143;

assign local_bb4__42_i143 = (local_bb4_tobool213_i138 & local_bb4_not_cmp37_i142);

// This section implements an unregistered operation.
// 
wire local_bb4_or2_i_i121_stall_local;
wire [31:0] local_bb4_or2_i_i121;

assign local_bb4_or2_i_i121 = ((local_bb4_shr1_i_i120 & 32'h1FFFFFF) | (local_bb4_or_i_i119 & 32'h7FFFFFF));

// This section implements a registered operation.
// 
wire local_bb4_sum_321_push9___inputs_ready;
 reg local_bb4_sum_321_push9___valid_out_NO_SHIFT_REG;
wire local_bb4_sum_321_push9___stall_in;
wire local_bb4_sum_321_push9___output_regs_ready;
wire [31:0] local_bb4_sum_321_push9___result;
wire local_bb4_sum_321_push9___fu_valid_out;
wire local_bb4_sum_321_push9___fu_stall_out;
 reg [31:0] local_bb4_sum_321_push9___NO_SHIFT_REG;
wire local_bb4_sum_321_push9___causedstall;

acl_push local_bb4_sum_321_push9___feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_238to239_bb4_c1_ene6_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_238to239_bb4___0_NO_SHIFT_REG),
	.stall_out(local_bb4_sum_321_push9___fu_stall_out),
	.valid_in(SFC_3_VALID_238_239_0_NO_SHIFT_REG),
	.valid_out(local_bb4_sum_321_push9___fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_sum_321_push9___result),
	.feedback_out(feedback_data_out_9),
	.feedback_valid_out(feedback_valid_out_9),
	.feedback_stall_in(feedback_stall_in_9)
);

defparam local_bb4_sum_321_push9___feedback.STALLFREE = 1;
defparam local_bb4_sum_321_push9___feedback.DATA_WIDTH = 32;
defparam local_bb4_sum_321_push9___feedback.FIFO_DEPTH = 9;
defparam local_bb4_sum_321_push9___feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_sum_321_push9___feedback.STYLE = "REGULAR";

assign local_bb4_sum_321_push9___inputs_ready = 1'b1;
assign local_bb4_sum_321_push9___output_regs_ready = 1'b1;
assign SFC_3_VALID_238_239_0_stall_in_1 = 1'b0;
assign rnode_238to239_bb4___0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_238to239_bb4_c1_ene6_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign local_bb4_sum_321_push9___causedstall = (SFC_3_VALID_238_239_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_sum_321_push9___NO_SHIFT_REG <= 'x;
		local_bb4_sum_321_push9___valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_sum_321_push9___output_regs_ready)
		begin
			local_bb4_sum_321_push9___NO_SHIFT_REG <= local_bb4_sum_321_push9___result;
			local_bb4_sum_321_push9___valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_sum_321_push9___stall_in))
			begin
				local_bb4_sum_321_push9___valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_239to240_bb4___0_valid_out_NO_SHIFT_REG;
 logic rnode_239to240_bb4___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_239to240_bb4___0_NO_SHIFT_REG;
 logic rnode_239to240_bb4___0_reg_240_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_239to240_bb4___0_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4___0_valid_out_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4___0_stall_in_reg_240_NO_SHIFT_REG;
 logic rnode_239to240_bb4___0_stall_out_reg_240_NO_SHIFT_REG;

acl_data_fifo rnode_239to240_bb4___0_reg_240_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_239to240_bb4___0_reg_240_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_239to240_bb4___0_stall_in_reg_240_NO_SHIFT_REG),
	.valid_out(rnode_239to240_bb4___0_valid_out_reg_240_NO_SHIFT_REG),
	.stall_out(rnode_239to240_bb4___0_stall_out_reg_240_NO_SHIFT_REG),
	.data_in(rnode_238to239_bb4___1_NO_SHIFT_REG),
	.data_out(rnode_239to240_bb4___0_reg_240_NO_SHIFT_REG)
);

defparam rnode_239to240_bb4___0_reg_240_fifo.DEPTH = 1;
defparam rnode_239to240_bb4___0_reg_240_fifo.DATA_WIDTH = 32;
defparam rnode_239to240_bb4___0_reg_240_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_239to240_bb4___0_reg_240_fifo.IMPL = "shift_reg";

assign rnode_239to240_bb4___0_reg_240_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_238to239_bb4___0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_239to240_bb4___0_NO_SHIFT_REG = rnode_239to240_bb4___0_reg_240_NO_SHIFT_REG;
assign rnode_239to240_bb4___0_stall_in_reg_240_NO_SHIFT_REG = 1'b0;
assign rnode_239to240_bb4___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4__43_i144_stall_local;
wire [31:0] local_bb4__43_i144;

assign local_bb4__43_i144 = (local_bb4__42_i143 ? 32'h0 : (local_bb4__pre_i137 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_shr3_i_i122_stall_local;
wire [31:0] local_bb4_shr3_i_i122;

assign local_bb4_shr3_i_i122 = ((local_bb4_or2_i_i121 & 32'h7FFFFFF) >> 32'h4);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_240to241_bb4_sum_321_push9___0_valid_out_NO_SHIFT_REG;
 logic rnode_240to241_bb4_sum_321_push9___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_sum_321_push9___0_NO_SHIFT_REG;
 logic rnode_240to241_bb4_sum_321_push9___0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4_sum_321_push9___0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_sum_321_push9___0_valid_out_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_sum_321_push9___0_stall_in_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4_sum_321_push9___0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_240to241_bb4_sum_321_push9___0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to241_bb4_sum_321_push9___0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to241_bb4_sum_321_push9___0_stall_in_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_240to241_bb4_sum_321_push9___0_valid_out_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_240to241_bb4_sum_321_push9___0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in(local_bb4_sum_321_push9___NO_SHIFT_REG),
	.data_out(rnode_240to241_bb4_sum_321_push9___0_reg_241_NO_SHIFT_REG)
);

defparam rnode_240to241_bb4_sum_321_push9___0_reg_241_fifo.DEPTH = 1;
defparam rnode_240to241_bb4_sum_321_push9___0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_240to241_bb4_sum_321_push9___0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to241_bb4_sum_321_push9___0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_240to241_bb4_sum_321_push9___0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_sum_321_push9___stall_in = 1'b0;
assign rnode_240to241_bb4_sum_321_push9___0_NO_SHIFT_REG = rnode_240to241_bb4_sum_321_push9___0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4_sum_321_push9___0_stall_in_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_sum_321_push9___0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_240to244_bb4___0_valid_out_NO_SHIFT_REG;
 logic rnode_240to244_bb4___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_240to244_bb4___0_NO_SHIFT_REG;
 logic rnode_240to244_bb4___0_reg_244_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_240to244_bb4___0_reg_244_NO_SHIFT_REG;
 logic rnode_240to244_bb4___0_valid_out_reg_244_NO_SHIFT_REG;
 logic rnode_240to244_bb4___0_stall_in_reg_244_NO_SHIFT_REG;
 logic rnode_240to244_bb4___0_stall_out_reg_244_NO_SHIFT_REG;

acl_data_fifo rnode_240to244_bb4___0_reg_244_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to244_bb4___0_reg_244_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to244_bb4___0_stall_in_reg_244_NO_SHIFT_REG),
	.valid_out(rnode_240to244_bb4___0_valid_out_reg_244_NO_SHIFT_REG),
	.stall_out(rnode_240to244_bb4___0_stall_out_reg_244_NO_SHIFT_REG),
	.data_in(rnode_239to240_bb4___0_NO_SHIFT_REG),
	.data_out(rnode_240to244_bb4___0_reg_244_NO_SHIFT_REG)
);

defparam rnode_240to244_bb4___0_reg_244_fifo.DEPTH = 4;
defparam rnode_240to244_bb4___0_reg_244_fifo.DATA_WIDTH = 32;
defparam rnode_240to244_bb4___0_reg_244_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to244_bb4___0_reg_244_fifo.IMPL = "shift_reg";

assign rnode_240to244_bb4___0_reg_244_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_239to240_bb4___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_240to244_bb4___0_NO_SHIFT_REG = rnode_240to244_bb4___0_reg_244_NO_SHIFT_REG;
assign rnode_240to244_bb4___0_stall_in_reg_244_NO_SHIFT_REG = 1'b0;
assign rnode_240to244_bb4___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_or4_i_i123_stall_local;
wire [31:0] local_bb4_or4_i_i123;

assign local_bb4_or4_i_i123 = ((local_bb4_shr3_i_i122 & 32'h7FFFFF) | (local_bb4_or2_i_i121 & 32'h7FFFFFF));

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_241to244_bb4_sum_321_push9___0_valid_out_NO_SHIFT_REG;
 logic rnode_241to244_bb4_sum_321_push9___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_241to244_bb4_sum_321_push9___0_NO_SHIFT_REG;
 logic rnode_241to244_bb4_sum_321_push9___0_reg_244_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_241to244_bb4_sum_321_push9___0_reg_244_NO_SHIFT_REG;
 logic rnode_241to244_bb4_sum_321_push9___0_valid_out_reg_244_NO_SHIFT_REG;
 logic rnode_241to244_bb4_sum_321_push9___0_stall_in_reg_244_NO_SHIFT_REG;
 logic rnode_241to244_bb4_sum_321_push9___0_stall_out_reg_244_NO_SHIFT_REG;

acl_data_fifo rnode_241to244_bb4_sum_321_push9___0_reg_244_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to244_bb4_sum_321_push9___0_reg_244_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to244_bb4_sum_321_push9___0_stall_in_reg_244_NO_SHIFT_REG),
	.valid_out(rnode_241to244_bb4_sum_321_push9___0_valid_out_reg_244_NO_SHIFT_REG),
	.stall_out(rnode_241to244_bb4_sum_321_push9___0_stall_out_reg_244_NO_SHIFT_REG),
	.data_in(rnode_240to241_bb4_sum_321_push9___0_NO_SHIFT_REG),
	.data_out(rnode_241to244_bb4_sum_321_push9___0_reg_244_NO_SHIFT_REG)
);

defparam rnode_241to244_bb4_sum_321_push9___0_reg_244_fifo.DEPTH = 3;
defparam rnode_241to244_bb4_sum_321_push9___0_reg_244_fifo.DATA_WIDTH = 32;
defparam rnode_241to244_bb4_sum_321_push9___0_reg_244_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to244_bb4_sum_321_push9___0_reg_244_fifo.IMPL = "shift_reg";

assign rnode_241to244_bb4_sum_321_push9___0_reg_244_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4_sum_321_push9___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_241to244_bb4_sum_321_push9___0_NO_SHIFT_REG = rnode_241to244_bb4_sum_321_push9___0_reg_244_NO_SHIFT_REG;
assign rnode_241to244_bb4_sum_321_push9___0_stall_in_reg_244_NO_SHIFT_REG = 1'b0;
assign rnode_241to244_bb4_sum_321_push9___0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_244to245_bb4___0_valid_out_0_NO_SHIFT_REG;
 logic rnode_244to245_bb4___0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4___0_NO_SHIFT_REG;
 logic rnode_244to245_bb4___0_valid_out_1_NO_SHIFT_REG;
 logic rnode_244to245_bb4___0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4___1_NO_SHIFT_REG;
 logic rnode_244to245_bb4___0_reg_245_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4___0_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4___0_valid_out_0_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4___0_stall_in_0_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4___0_stall_out_reg_245_NO_SHIFT_REG;

acl_data_fifo rnode_244to245_bb4___0_reg_245_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_244to245_bb4___0_reg_245_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_244to245_bb4___0_stall_in_0_reg_245_NO_SHIFT_REG),
	.valid_out(rnode_244to245_bb4___0_valid_out_0_reg_245_NO_SHIFT_REG),
	.stall_out(rnode_244to245_bb4___0_stall_out_reg_245_NO_SHIFT_REG),
	.data_in(rnode_240to244_bb4___0_NO_SHIFT_REG),
	.data_out(rnode_244to245_bb4___0_reg_245_NO_SHIFT_REG)
);

defparam rnode_244to245_bb4___0_reg_245_fifo.DEPTH = 1;
defparam rnode_244to245_bb4___0_reg_245_fifo.DATA_WIDTH = 32;
defparam rnode_244to245_bb4___0_reg_245_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_244to245_bb4___0_reg_245_fifo.IMPL = "shift_reg";

assign rnode_244to245_bb4___0_reg_245_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_240to244_bb4___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_244to245_bb4___0_stall_in_0_reg_245_NO_SHIFT_REG = 1'b0;
assign rnode_244to245_bb4___0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_244to245_bb4___0_NO_SHIFT_REG = rnode_244to245_bb4___0_reg_245_NO_SHIFT_REG;
assign rnode_244to245_bb4___0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_244to245_bb4___1_NO_SHIFT_REG = rnode_244to245_bb4___0_reg_245_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_shr5_i_i124_stall_local;
wire [31:0] local_bb4_shr5_i_i124;

assign local_bb4_shr5_i_i124 = ((local_bb4_or4_i_i123 & 32'h7FFFFFF) >> 32'h8);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_244to245_bb4_sum_321_push9___0_valid_out_NO_SHIFT_REG;
 logic rnode_244to245_bb4_sum_321_push9___0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4_sum_321_push9___0_NO_SHIFT_REG;
 logic rnode_244to245_bb4_sum_321_push9___0_reg_245_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4_sum_321_push9___0_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4_sum_321_push9___0_valid_out_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4_sum_321_push9___0_stall_in_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4_sum_321_push9___0_stall_out_reg_245_NO_SHIFT_REG;

acl_data_fifo rnode_244to245_bb4_sum_321_push9___0_reg_245_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_244to245_bb4_sum_321_push9___0_reg_245_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_244to245_bb4_sum_321_push9___0_stall_in_reg_245_NO_SHIFT_REG),
	.valid_out(rnode_244to245_bb4_sum_321_push9___0_valid_out_reg_245_NO_SHIFT_REG),
	.stall_out(rnode_244to245_bb4_sum_321_push9___0_stall_out_reg_245_NO_SHIFT_REG),
	.data_in(rnode_241to244_bb4_sum_321_push9___0_NO_SHIFT_REG),
	.data_out(rnode_244to245_bb4_sum_321_push9___0_reg_245_NO_SHIFT_REG)
);

defparam rnode_244to245_bb4_sum_321_push9___0_reg_245_fifo.DEPTH = 1;
defparam rnode_244to245_bb4_sum_321_push9___0_reg_245_fifo.DATA_WIDTH = 32;
defparam rnode_244to245_bb4_sum_321_push9___0_reg_245_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_244to245_bb4_sum_321_push9___0_reg_245_fifo.IMPL = "shift_reg";

assign rnode_244to245_bb4_sum_321_push9___0_reg_245_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_241to244_bb4_sum_321_push9___0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_244to245_bb4_sum_321_push9___0_NO_SHIFT_REG = rnode_244to245_bb4_sum_321_push9___0_reg_245_NO_SHIFT_REG;
assign rnode_244to245_bb4_sum_321_push9___0_stall_in_reg_245_NO_SHIFT_REG = 1'b0;
assign rnode_244to245_bb4_sum_321_push9___0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4____valid_out;
wire local_bb4____stall_in;
wire local_bb4____inputs_ready;
wire local_bb4____stall_local;
 reg [31:0] ffwd_10_0_reg_NO_SHIFT_REG;

assign local_bb4____inputs_ready = (SFC_3_VALID_244_245_0_valid_out_1_NO_SHIFT_REG & rnode_244to245_bb4___0_valid_out_0_NO_SHIFT_REG);
assign ffwd_10_0 = ffwd_10_0_reg_NO_SHIFT_REG;
assign local_bb4____valid_out = 1'b1;
assign SFC_3_VALID_244_245_0_stall_in_1 = 1'b0;
assign rnode_244to245_bb4___0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock)
begin
	if ((1'b1 & SFC_3_VALID_244_245_0_NO_SHIFT_REG))
	begin
		ffwd_10_0_reg_NO_SHIFT_REG <= rnode_244to245_bb4___0_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_exi1_stall_local;
wire [95:0] local_bb4_c1_exi1;

assign local_bb4_c1_exi1[31:0] = 32'bx;
assign local_bb4_c1_exi1[63:32] = rnode_244to245_bb4___1_NO_SHIFT_REG;
assign local_bb4_c1_exi1[95:64] = 32'bx;

// This section implements an unregistered operation.
// 
wire local_bb4_or6_i_i125_stall_local;
wire [31:0] local_bb4_or6_i_i125;

assign local_bb4_or6_i_i125 = ((local_bb4_shr5_i_i124 & 32'h7FFFF) | (local_bb4_or4_i_i123 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_shr7_i_i126_stall_local;
wire [31:0] local_bb4_shr7_i_i126;

assign local_bb4_shr7_i_i126 = ((local_bb4_or6_i_i125 & 32'h7FFFFFF) >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb4_or6_masked_i_i127_stall_local;
wire [31:0] local_bb4_or6_masked_i_i127;

assign local_bb4_or6_masked_i_i127 = ((local_bb4_or6_i_i125 & 32'h7FFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_neg_i_i128_stall_local;
wire [31:0] local_bb4_neg_i_i128;

assign local_bb4_neg_i_i128 = ((local_bb4_or6_masked_i_i127 & 32'h7FFFFFF) | (local_bb4_shr7_i_i126 & 32'h7FF));

// This section implements an unregistered operation.
// 
wire local_bb4_and_i_i129_stall_local;
wire [31:0] local_bb4_and_i_i129;

assign local_bb4_and_i_i129 = ((local_bb4_neg_i_i128 & 32'h7FFFFFF) ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__and_i_i129_valid_out;
wire local_bb4__and_i_i129_stall_in;
wire local_bb4__and_i_i129_inputs_ready;
wire local_bb4__and_i_i129_stall_local;
wire [31:0] local_bb4__and_i_i129;

thirtysix_six_comp local_bb4__and_i_i129_popcnt_instance (
	.data((local_bb4_and_i_i129 & 32'h7FFFFFF)),
	.sum(local_bb4__and_i_i129)
);


assign local_bb4__and_i_i129_inputs_ready = rnode_239to240_bb4_add192_i113_0_valid_out_3_NO_SHIFT_REG;
assign local_bb4__and_i_i129_valid_out = 1'b1;
assign rnode_239to240_bb4_add192_i113_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_240to241_bb4__and_i_i129_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4__and_i_i129_0_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4__and_i_i129_1_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4__and_i_i129_2_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_reg_241_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_240to241_bb4__and_i_i129_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_valid_out_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_stall_in_0_reg_241_NO_SHIFT_REG;
 logic rnode_240to241_bb4__and_i_i129_0_stall_out_reg_241_NO_SHIFT_REG;

acl_data_fifo rnode_240to241_bb4__and_i_i129_0_reg_241_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_240to241_bb4__and_i_i129_0_reg_241_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_240to241_bb4__and_i_i129_0_stall_in_0_reg_241_NO_SHIFT_REG),
	.valid_out(rnode_240to241_bb4__and_i_i129_0_valid_out_0_reg_241_NO_SHIFT_REG),
	.stall_out(rnode_240to241_bb4__and_i_i129_0_stall_out_reg_241_NO_SHIFT_REG),
	.data_in((local_bb4__and_i_i129 & 32'h3F)),
	.data_out(rnode_240to241_bb4__and_i_i129_0_reg_241_NO_SHIFT_REG)
);

defparam rnode_240to241_bb4__and_i_i129_0_reg_241_fifo.DEPTH = 1;
defparam rnode_240to241_bb4__and_i_i129_0_reg_241_fifo.DATA_WIDTH = 32;
defparam rnode_240to241_bb4__and_i_i129_0_reg_241_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_240to241_bb4__and_i_i129_0_reg_241_fifo.IMPL = "shift_reg";

assign rnode_240to241_bb4__and_i_i129_0_reg_241_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__and_i_i129_stall_in = 1'b0;
assign rnode_240to241_bb4__and_i_i129_0_stall_in_0_reg_241_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4__and_i_i129_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4__and_i_i129_0_NO_SHIFT_REG = rnode_240to241_bb4__and_i_i129_0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4__and_i_i129_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4__and_i_i129_1_NO_SHIFT_REG = rnode_240to241_bb4__and_i_i129_0_reg_241_NO_SHIFT_REG;
assign rnode_240to241_bb4__and_i_i129_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_240to241_bb4__and_i_i129_2_NO_SHIFT_REG = rnode_240to241_bb4__and_i_i129_0_reg_241_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_and9_i_i130_stall_local;
wire [31:0] local_bb4_and9_i_i130;

assign local_bb4_and9_i_i130 = ((rnode_240to241_bb4__and_i_i129_0_NO_SHIFT_REG & 32'h3F) & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb4_and203_i131_stall_local;
wire [31:0] local_bb4_and203_i131;

assign local_bb4_and203_i131 = ((rnode_240to241_bb4__and_i_i129_1_NO_SHIFT_REG & 32'h3F) & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb4_and206_i133_stall_local;
wire [31:0] local_bb4_and206_i133;

assign local_bb4_and206_i133 = ((rnode_240to241_bb4__and_i_i129_2_NO_SHIFT_REG & 32'h3F) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_sub239_i152_stall_local;
wire [31:0] local_bb4_sub239_i152;

assign local_bb4_sub239_i152 = (32'h0 - (local_bb4_and9_i_i130 & 32'h1F));

// This section implements an unregistered operation.
// 
wire local_bb4_shl204_i132_stall_local;
wire [31:0] local_bb4_shl204_i132;

assign local_bb4_shl204_i132 = ((rnode_240to241_bb4_and193_i114_0_NO_SHIFT_REG & 32'hFFFFFFF) << (local_bb4_and203_i131 & 32'h18));

// This section implements an unregistered operation.
// 
wire local_bb4_cond244_i153_stall_local;
wire [31:0] local_bb4_cond244_i153;

assign local_bb4_cond244_i153 = (rnode_239to241_bb4_cmp37_i36_2_NO_SHIFT_REG ? local_bb4_sub239_i152 : (local_bb4__43_i144 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and205_i134_stall_local;
wire [31:0] local_bb4_and205_i134;

assign local_bb4_and205_i134 = (local_bb4_shl204_i132 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_add245_i154_stall_local;
wire [31:0] local_bb4_add245_i154;

assign local_bb4_add245_i154 = (local_bb4_cond244_i153 + (rnode_239to241_bb4_and17_i25_0_NO_SHIFT_REG & 32'hFF));

// This section implements an unregistered operation.
// 
wire local_bb4_fold_i156_stall_local;
wire [31:0] local_bb4_fold_i156;

assign local_bb4_fold_i156 = (local_bb4_cond244_i153 + (rnode_239to241_bb4_shr16_i24_0_NO_SHIFT_REG & 32'h1FF));

// This section implements an unregistered operation.
// 
wire local_bb4_shl207_i135_stall_local;
wire [31:0] local_bb4_shl207_i135;

assign local_bb4_shl207_i135 = ((local_bb4_and205_i134 & 32'h7FFFFFF) << (local_bb4_and206_i133 & 32'h7));

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i157_stall_local;
wire [31:0] local_bb4_and250_i157;

assign local_bb4_and250_i157 = (local_bb4_fold_i156 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and269_i168_stall_local;
wire [31:0] local_bb4_and269_i168;

assign local_bb4_and269_i168 = (local_bb4_fold_i156 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb4_and208_i136_stall_local;
wire [31:0] local_bb4_and208_i136;

assign local_bb4_and208_i136 = (local_bb4_shl207_i135 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__44_i145_stall_local;
wire [31:0] local_bb4__44_i145;

assign local_bb4__44_i145 = (local_bb4__40_demorgan_i141 ? (local_bb4_and208_i136 & 32'h7FFFFFF) : (local_bb4_or219_i140 & 32'h7FFFFFF));

// This section implements an unregistered operation.
// 
wire local_bb4_and250_i157_valid_out;
wire local_bb4_and250_i157_stall_in;
wire local_bb4_and269_i168_valid_out;
wire local_bb4_and269_i168_stall_in;
wire local_bb4_add245_i154_valid_out;
wire local_bb4_add245_i154_stall_in;
wire local_bb4__45_i146_valid_out;
wire local_bb4__45_i146_stall_in;
wire local_bb4_not_cmp37_i142_valid_out_1;
wire local_bb4_not_cmp37_i142_stall_in_1;
wire local_bb4__45_i146_inputs_ready;
wire local_bb4__45_i146_stall_local;
wire [31:0] local_bb4__45_i146;

assign local_bb4__45_i146_inputs_ready = (rnode_239to241_bb4_shr16_i24_0_valid_out_NO_SHIFT_REG & rnode_239to241_bb4_and17_i25_0_valid_out_NO_SHIFT_REG & rnode_239to241_bb4_cmp37_i36_0_valid_out_2_NO_SHIFT_REG & rnode_239to241_bb4_cmp37_i36_0_valid_out_0_NO_SHIFT_REG & rnode_240to241_bb4_and193_i114_0_valid_out_2_NO_SHIFT_REG & rnode_239to241_bb4_cmp37_i36_0_valid_out_1_NO_SHIFT_REG & rnode_240to241_bb4_and195_i115_0_valid_out_NO_SHIFT_REG & rnode_240to241_bb4_and193_i114_0_valid_out_1_NO_SHIFT_REG & rnode_240to241_bb4_and198_i116_0_valid_out_NO_SHIFT_REG & rnode_240to241_bb4_and193_i114_0_valid_out_0_NO_SHIFT_REG & rnode_240to241_bb4__and_i_i129_0_valid_out_1_NO_SHIFT_REG & rnode_240to241_bb4__and_i_i129_0_valid_out_2_NO_SHIFT_REG & rnode_240to241_bb4__and_i_i129_0_valid_out_0_NO_SHIFT_REG);
assign local_bb4__45_i146 = (local_bb4__42_i143 ? (rnode_240to241_bb4_and193_i114_2_NO_SHIFT_REG & 32'hFFFFFFF) : (local_bb4__44_i145 & 32'h7FFFFFF));
assign local_bb4_and250_i157_valid_out = 1'b1;
assign local_bb4_and269_i168_valid_out = 1'b1;
assign local_bb4_add245_i154_valid_out = 1'b1;
assign local_bb4__45_i146_valid_out = 1'b1;
assign local_bb4_not_cmp37_i142_valid_out_1 = 1'b1;
assign rnode_239to241_bb4_shr16_i24_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_and17_i25_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_cmp37_i36_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_cmp37_i36_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and193_i114_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_239to241_bb4_cmp37_i36_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and195_i115_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and193_i114_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and198_i116_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4_and193_i114_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4__and_i_i129_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4__and_i_i129_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_240to241_bb4__and_i_i129_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_241to242_bb4_and250_i157_0_valid_out_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and250_i157_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4_and250_i157_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and250_i157_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4_and250_i157_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and250_i157_0_valid_out_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and250_i157_0_stall_in_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_and250_i157_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_241to242_bb4_and250_i157_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to242_bb4_and250_i157_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to242_bb4_and250_i157_0_stall_in_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_241to242_bb4_and250_i157_0_valid_out_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_241to242_bb4_and250_i157_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in((local_bb4_and250_i157 & 32'hFF)),
	.data_out(rnode_241to242_bb4_and250_i157_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_241to242_bb4_and250_i157_0_reg_242_fifo.DEPTH = 1;
defparam rnode_241to242_bb4_and250_i157_0_reg_242_fifo.DATA_WIDTH = 32;
defparam rnode_241to242_bb4_and250_i157_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to242_bb4_and250_i157_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_241to242_bb4_and250_i157_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and250_i157_stall_in = 1'b0;
assign rnode_241to242_bb4_and250_i157_0_NO_SHIFT_REG = rnode_241to242_bb4_and250_i157_0_reg_242_NO_SHIFT_REG;
assign rnode_241to242_bb4_and250_i157_0_stall_in_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_and250_i157_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_241to243_bb4_and269_i168_0_valid_out_NO_SHIFT_REG;
 logic rnode_241to243_bb4_and269_i168_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_241to243_bb4_and269_i168_0_NO_SHIFT_REG;
 logic rnode_241to243_bb4_and269_i168_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_241to243_bb4_and269_i168_0_reg_243_NO_SHIFT_REG;
 logic rnode_241to243_bb4_and269_i168_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_241to243_bb4_and269_i168_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_241to243_bb4_and269_i168_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_241to243_bb4_and269_i168_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to243_bb4_and269_i168_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to243_bb4_and269_i168_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_241to243_bb4_and269_i168_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_241to243_bb4_and269_i168_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in((local_bb4_and269_i168 & 32'hFF800000)),
	.data_out(rnode_241to243_bb4_and269_i168_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_241to243_bb4_and269_i168_0_reg_243_fifo.DEPTH = 2;
defparam rnode_241to243_bb4_and269_i168_0_reg_243_fifo.DATA_WIDTH = 32;
defparam rnode_241to243_bb4_and269_i168_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to243_bb4_and269_i168_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_241to243_bb4_and269_i168_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_and269_i168_stall_in = 1'b0;
assign rnode_241to243_bb4_and269_i168_0_NO_SHIFT_REG = rnode_241to243_bb4_and269_i168_0_reg_243_NO_SHIFT_REG;
assign rnode_241to243_bb4_and269_i168_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_241to243_bb4_and269_i168_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_241to242_bb4_add245_i154_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4_add245_i154_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4_add245_i154_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4_add245_i154_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_241to242_bb4_add245_i154_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4_add245_i154_1_NO_SHIFT_REG;
 logic rnode_241to242_bb4_add245_i154_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4_add245_i154_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_add245_i154_0_valid_out_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_add245_i154_0_stall_in_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_add245_i154_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_241to242_bb4_add245_i154_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to242_bb4_add245_i154_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to242_bb4_add245_i154_0_stall_in_0_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_241to242_bb4_add245_i154_0_valid_out_0_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_241to242_bb4_add245_i154_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in(local_bb4_add245_i154),
	.data_out(rnode_241to242_bb4_add245_i154_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_241to242_bb4_add245_i154_0_reg_242_fifo.DEPTH = 1;
defparam rnode_241to242_bb4_add245_i154_0_reg_242_fifo.DATA_WIDTH = 32;
defparam rnode_241to242_bb4_add245_i154_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to242_bb4_add245_i154_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_241to242_bb4_add245_i154_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_add245_i154_stall_in = 1'b0;
assign rnode_241to242_bb4_add245_i154_0_stall_in_0_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_add245_i154_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_241to242_bb4_add245_i154_0_NO_SHIFT_REG = rnode_241to242_bb4_add245_i154_0_reg_242_NO_SHIFT_REG;
assign rnode_241to242_bb4_add245_i154_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_241to242_bb4_add245_i154_1_NO_SHIFT_REG = rnode_241to242_bb4_add245_i154_0_reg_242_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_241to242_bb4__45_i146_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4__45_i146_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4__45_i146_1_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4__45_i146_2_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_241to242_bb4__45_i146_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_valid_out_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_stall_in_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4__45_i146_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_241to242_bb4__45_i146_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to242_bb4__45_i146_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to242_bb4__45_i146_0_stall_in_0_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_241to242_bb4__45_i146_0_valid_out_0_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_241to242_bb4__45_i146_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in((local_bb4__45_i146 & 32'hFFFFFFF)),
	.data_out(rnode_241to242_bb4__45_i146_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_241to242_bb4__45_i146_0_reg_242_fifo.DEPTH = 1;
defparam rnode_241to242_bb4__45_i146_0_reg_242_fifo.DATA_WIDTH = 32;
defparam rnode_241to242_bb4__45_i146_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to242_bb4__45_i146_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_241to242_bb4__45_i146_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__45_i146_stall_in = 1'b0;
assign rnode_241to242_bb4__45_i146_0_stall_in_0_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4__45_i146_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_241to242_bb4__45_i146_0_NO_SHIFT_REG = rnode_241to242_bb4__45_i146_0_reg_242_NO_SHIFT_REG;
assign rnode_241to242_bb4__45_i146_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_241to242_bb4__45_i146_1_NO_SHIFT_REG = rnode_241to242_bb4__45_i146_0_reg_242_NO_SHIFT_REG;
assign rnode_241to242_bb4__45_i146_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_241to242_bb4__45_i146_2_NO_SHIFT_REG = rnode_241to242_bb4__45_i146_0_reg_242_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_241to242_bb4_not_cmp37_i142_0_valid_out_NO_SHIFT_REG;
 logic rnode_241to242_bb4_not_cmp37_i142_0_stall_in_NO_SHIFT_REG;
 logic rnode_241to242_bb4_not_cmp37_i142_0_NO_SHIFT_REG;
 logic rnode_241to242_bb4_not_cmp37_i142_0_reg_242_inputs_ready_NO_SHIFT_REG;
 logic rnode_241to242_bb4_not_cmp37_i142_0_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_not_cmp37_i142_0_valid_out_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_not_cmp37_i142_0_stall_in_reg_242_NO_SHIFT_REG;
 logic rnode_241to242_bb4_not_cmp37_i142_0_stall_out_reg_242_NO_SHIFT_REG;

acl_data_fifo rnode_241to242_bb4_not_cmp37_i142_0_reg_242_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_241to242_bb4_not_cmp37_i142_0_reg_242_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_241to242_bb4_not_cmp37_i142_0_stall_in_reg_242_NO_SHIFT_REG),
	.valid_out(rnode_241to242_bb4_not_cmp37_i142_0_valid_out_reg_242_NO_SHIFT_REG),
	.stall_out(rnode_241to242_bb4_not_cmp37_i142_0_stall_out_reg_242_NO_SHIFT_REG),
	.data_in(local_bb4_not_cmp37_i142),
	.data_out(rnode_241to242_bb4_not_cmp37_i142_0_reg_242_NO_SHIFT_REG)
);

defparam rnode_241to242_bb4_not_cmp37_i142_0_reg_242_fifo.DEPTH = 1;
defparam rnode_241to242_bb4_not_cmp37_i142_0_reg_242_fifo.DATA_WIDTH = 1;
defparam rnode_241to242_bb4_not_cmp37_i142_0_reg_242_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_241to242_bb4_not_cmp37_i142_0_reg_242_fifo.IMPL = "shift_reg";

assign rnode_241to242_bb4_not_cmp37_i142_0_reg_242_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_not_cmp37_i142_stall_in_1 = 1'b0;
assign rnode_241to242_bb4_not_cmp37_i142_0_NO_SHIFT_REG = rnode_241to242_bb4_not_cmp37_i142_0_reg_242_NO_SHIFT_REG;
assign rnode_241to242_bb4_not_cmp37_i142_0_stall_in_reg_242_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_not_cmp37_i142_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_notrhs_i159_stall_local;
wire local_bb4_notrhs_i159;

assign local_bb4_notrhs_i159 = ((rnode_241to242_bb4_and250_i157_0_NO_SHIFT_REG & 32'hFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_shl273_i169_stall_local;
wire [31:0] local_bb4_shl273_i169;

assign local_bb4_shl273_i169 = ((rnode_241to243_bb4_and269_i168_0_NO_SHIFT_REG & 32'hFF800000) & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb4_and247_i155_stall_local;
wire [31:0] local_bb4_and247_i155;

assign local_bb4_and247_i155 = (rnode_241to242_bb4_add245_i154_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp258_i162_stall_local;
wire local_bb4_cmp258_i162;

assign local_bb4_cmp258_i162 = ($signed(rnode_241to242_bb4_add245_i154_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb4_and225_i147_stall_local;
wire [31:0] local_bb4_and225_i147;

assign local_bb4_and225_i147 = ((rnode_241to242_bb4__45_i146_0_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_and270_i165_stall_local;
wire [31:0] local_bb4_and270_i165;

assign local_bb4_and270_i165 = ((rnode_241to242_bb4__45_i146_1_NO_SHIFT_REG & 32'hFFFFFFF) & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb4_shr271_i166_valid_out;
wire local_bb4_shr271_i166_stall_in;
wire local_bb4_shr271_i166_inputs_ready;
wire local_bb4_shr271_i166_stall_local;
wire [31:0] local_bb4_shr271_i166;

assign local_bb4_shr271_i166_inputs_ready = rnode_241to242_bb4__45_i146_0_valid_out_2_NO_SHIFT_REG;
assign local_bb4_shr271_i166 = ((rnode_241to242_bb4__45_i146_2_NO_SHIFT_REG & 32'hFFFFFFF) >> 32'h3);
assign local_bb4_shr271_i166_valid_out = 1'b1;
assign rnode_241to242_bb4__45_i146_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb4_notlhs_i158_stall_local;
wire local_bb4_notlhs_i158;

assign local_bb4_notlhs_i158 = ((local_bb4_and247_i155 & 32'h100) != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_i148_stall_local;
wire local_bb4_cmp226_i148;

assign local_bb4_cmp226_i148 = ((local_bb4_and225_i147 & 32'h7FFFFFF) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i180_stall_local;
wire local_bb4_cmp296_i180;

assign local_bb4_cmp296_i180 = ((local_bb4_and270_i165 & 32'h7) > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp296_i180_valid_out;
wire local_bb4_cmp296_i180_stall_in;
wire local_bb4_cmp299_i181_valid_out;
wire local_bb4_cmp299_i181_stall_in;
wire local_bb4_cmp299_i181_inputs_ready;
wire local_bb4_cmp299_i181_stall_local;
wire local_bb4_cmp299_i181;

assign local_bb4_cmp299_i181_inputs_ready = rnode_241to242_bb4__45_i146_0_valid_out_1_NO_SHIFT_REG;
assign local_bb4_cmp299_i181 = ((local_bb4_and270_i165 & 32'h7) == 32'h4);
assign local_bb4_cmp296_i180_valid_out = 1'b1;
assign local_bb4_cmp299_i181_valid_out = 1'b1;
assign rnode_241to242_bb4__45_i146_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4_shr271_i166_0_valid_out_NO_SHIFT_REG;
 logic rnode_242to243_bb4_shr271_i166_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_242to243_bb4_shr271_i166_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_shr271_i166_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_242to243_bb4_shr271_i166_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_shr271_i166_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_shr271_i166_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_shr271_i166_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4_shr271_i166_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4_shr271_i166_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4_shr271_i166_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4_shr271_i166_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4_shr271_i166_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in((local_bb4_shr271_i166 & 32'h1FFFFFF)),
	.data_out(rnode_242to243_bb4_shr271_i166_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4_shr271_i166_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4_shr271_i166_0_reg_243_fifo.DATA_WIDTH = 32;
defparam rnode_242to243_bb4_shr271_i166_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4_shr271_i166_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4_shr271_i166_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_shr271_i166_stall_in = 1'b0;
assign rnode_242to243_bb4_shr271_i166_0_NO_SHIFT_REG = rnode_242to243_bb4_shr271_i166_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_shr271_i166_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_shr271_i166_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_not__46_i160_stall_local;
wire local_bb4_not__46_i160;

assign local_bb4_not__46_i160 = (local_bb4_notrhs_i159 | local_bb4_notlhs_i158);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp226_not_i149_stall_local;
wire local_bb4_cmp226_not_i149;

assign local_bb4_cmp226_not_i149 = (local_bb4_cmp226_i148 ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4_cmp296_i180_0_valid_out_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp296_i180_0_stall_in_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp296_i180_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp296_i180_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp296_i180_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp296_i180_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp296_i180_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp296_i180_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4_cmp296_i180_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4_cmp296_i180_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4_cmp296_i180_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4_cmp296_i180_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4_cmp296_i180_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(local_bb4_cmp296_i180),
	.data_out(rnode_242to243_bb4_cmp296_i180_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4_cmp296_i180_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4_cmp296_i180_0_reg_243_fifo.DATA_WIDTH = 1;
defparam rnode_242to243_bb4_cmp296_i180_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4_cmp296_i180_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4_cmp296_i180_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp296_i180_stall_in = 1'b0;
assign rnode_242to243_bb4_cmp296_i180_0_NO_SHIFT_REG = rnode_242to243_bb4_cmp296_i180_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_cmp296_i180_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_cmp296_i180_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4_cmp299_i181_0_valid_out_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp299_i181_0_stall_in_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp299_i181_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp299_i181_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp299_i181_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp299_i181_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp299_i181_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_cmp299_i181_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4_cmp299_i181_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4_cmp299_i181_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4_cmp299_i181_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4_cmp299_i181_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4_cmp299_i181_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(local_bb4_cmp299_i181),
	.data_out(rnode_242to243_bb4_cmp299_i181_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4_cmp299_i181_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4_cmp299_i181_0_reg_243_fifo.DATA_WIDTH = 1;
defparam rnode_242to243_bb4_cmp299_i181_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4_cmp299_i181_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4_cmp299_i181_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_cmp299_i181_stall_in = 1'b0;
assign rnode_242to243_bb4_cmp299_i181_0_NO_SHIFT_REG = rnode_242to243_bb4_cmp299_i181_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_cmp299_i181_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_cmp299_i181_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb4_and272_i167_stall_local;
wire [31:0] local_bb4_and272_i167;

assign local_bb4_and272_i167 = ((rnode_242to243_bb4_shr271_i166_0_NO_SHIFT_REG & 32'h1FFFFFF) & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4__47_i161_stall_local;
wire local_bb4__47_i161;

assign local_bb4__47_i161 = (local_bb4_cmp226_i148 | local_bb4_not__46_i160);

// This section implements an unregistered operation.
// 
wire local_bb4_brmerge12_i150_stall_local;
wire local_bb4_brmerge12_i150;

assign local_bb4_brmerge12_i150 = (local_bb4_cmp226_not_i149 | rnode_241to242_bb4_not_cmp37_i142_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot262__i163_stall_local;
wire local_bb4_lnot262__i163;

assign local_bb4_lnot262__i163 = (local_bb4_cmp258_i162 & local_bb4_cmp226_not_i149);

// This section implements an unregistered operation.
// 
wire local_bb4_cmp29649_i184_stall_local;
wire [31:0] local_bb4_cmp29649_i184;

assign local_bb4_cmp29649_i184[31:1] = 31'h0;
assign local_bb4_cmp29649_i184[0] = rnode_242to243_bb4_cmp296_i180_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_conv300_i182_stall_local;
wire [31:0] local_bb4_conv300_i182;

assign local_bb4_conv300_i182[31:1] = 31'h0;
assign local_bb4_conv300_i182[0] = rnode_242to243_bb4_cmp299_i181_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or274_i170_stall_local;
wire [31:0] local_bb4_or274_i170;

assign local_bb4_or274_i170 = ((local_bb4_and272_i167 & 32'h7FFFFF) | (local_bb4_shl273_i169 & 32'h7F800000));

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i151_stall_local;
wire [31:0] local_bb4_resultSign_0_i151;

assign local_bb4_resultSign_0_i151 = (local_bb4_brmerge12_i150 ? (rnode_241to242_bb4_and35_i34_0_NO_SHIFT_REG & 32'h80000000) : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_resultSign_0_i151_valid_out;
wire local_bb4_resultSign_0_i151_stall_in;
wire local_bb4__47_i161_valid_out;
wire local_bb4__47_i161_stall_in;
wire local_bb4_or2662_i164_valid_out;
wire local_bb4_or2662_i164_stall_in;
wire local_bb4_or2662_i164_inputs_ready;
wire local_bb4_or2662_i164_stall_local;
wire local_bb4_or2662_i164;

assign local_bb4_or2662_i164_inputs_ready = (rnode_241to242_bb4_and35_i34_0_valid_out_NO_SHIFT_REG & rnode_241to242_bb4_not_cmp37_i142_0_valid_out_NO_SHIFT_REG & rnode_241to242_bb4_add245_i154_0_valid_out_0_NO_SHIFT_REG & rnode_241to242_bb4_and250_i157_0_valid_out_NO_SHIFT_REG & rnode_241to242_bb4__45_i146_0_valid_out_0_NO_SHIFT_REG & rnode_241to242_bb4_add245_i154_0_valid_out_1_NO_SHIFT_REG & rnode_241to242_bb4_var__u83_0_valid_out_NO_SHIFT_REG);
assign local_bb4_or2662_i164 = (rnode_241to242_bb4_var__u83_0_NO_SHIFT_REG | local_bb4_lnot262__i163);
assign local_bb4_resultSign_0_i151_valid_out = 1'b1;
assign local_bb4__47_i161_valid_out = 1'b1;
assign local_bb4_or2662_i164_valid_out = 1'b1;
assign rnode_241to242_bb4_and35_i34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_not_cmp37_i142_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_add245_i154_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_and250_i157_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4__45_i146_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_add245_i154_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_241to242_bb4_var__u83_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4_resultSign_0_i151_0_valid_out_NO_SHIFT_REG;
 logic rnode_242to243_bb4_resultSign_0_i151_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_242to243_bb4_resultSign_0_i151_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_resultSign_0_i151_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_242to243_bb4_resultSign_0_i151_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_resultSign_0_i151_0_valid_out_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_resultSign_0_i151_0_stall_in_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_resultSign_0_i151_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4_resultSign_0_i151_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4_resultSign_0_i151_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4_resultSign_0_i151_0_stall_in_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4_resultSign_0_i151_0_valid_out_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4_resultSign_0_i151_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in((local_bb4_resultSign_0_i151 & 32'h80000000)),
	.data_out(rnode_242to243_bb4_resultSign_0_i151_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4_resultSign_0_i151_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4_resultSign_0_i151_0_reg_243_fifo.DATA_WIDTH = 32;
defparam rnode_242to243_bb4_resultSign_0_i151_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4_resultSign_0_i151_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4_resultSign_0_i151_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_resultSign_0_i151_stall_in = 1'b0;
assign rnode_242to243_bb4_resultSign_0_i151_0_NO_SHIFT_REG = rnode_242to243_bb4_resultSign_0_i151_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_resultSign_0_i151_0_stall_in_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_resultSign_0_i151_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4__47_i161_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_valid_out_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_stall_in_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4__47_i161_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4__47_i161_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4__47_i161_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4__47_i161_0_stall_in_0_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4__47_i161_0_valid_out_0_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4__47_i161_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(local_bb4__47_i161),
	.data_out(rnode_242to243_bb4__47_i161_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4__47_i161_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4__47_i161_0_reg_243_fifo.DATA_WIDTH = 1;
defparam rnode_242to243_bb4__47_i161_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4__47_i161_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4__47_i161_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__47_i161_stall_in = 1'b0;
assign rnode_242to243_bb4__47_i161_0_stall_in_0_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__47_i161_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4__47_i161_0_NO_SHIFT_REG = rnode_242to243_bb4__47_i161_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4__47_i161_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4__47_i161_1_NO_SHIFT_REG = rnode_242to243_bb4__47_i161_0_reg_243_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_242to243_bb4_or2662_i164_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_1_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_2_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_reg_243_inputs_ready_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_valid_out_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_stall_in_0_reg_243_NO_SHIFT_REG;
 logic rnode_242to243_bb4_or2662_i164_0_stall_out_reg_243_NO_SHIFT_REG;

acl_data_fifo rnode_242to243_bb4_or2662_i164_0_reg_243_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_242to243_bb4_or2662_i164_0_reg_243_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_242to243_bb4_or2662_i164_0_stall_in_0_reg_243_NO_SHIFT_REG),
	.valid_out(rnode_242to243_bb4_or2662_i164_0_valid_out_0_reg_243_NO_SHIFT_REG),
	.stall_out(rnode_242to243_bb4_or2662_i164_0_stall_out_reg_243_NO_SHIFT_REG),
	.data_in(local_bb4_or2662_i164),
	.data_out(rnode_242to243_bb4_or2662_i164_0_reg_243_NO_SHIFT_REG)
);

defparam rnode_242to243_bb4_or2662_i164_0_reg_243_fifo.DEPTH = 1;
defparam rnode_242to243_bb4_or2662_i164_0_reg_243_fifo.DATA_WIDTH = 1;
defparam rnode_242to243_bb4_or2662_i164_0_reg_243_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_242to243_bb4_or2662_i164_0_reg_243_fifo.IMPL = "shift_reg";

assign rnode_242to243_bb4_or2662_i164_0_reg_243_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4_or2662_i164_stall_in = 1'b0;
assign rnode_242to243_bb4_or2662_i164_0_stall_in_0_reg_243_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_or2662_i164_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4_or2662_i164_0_NO_SHIFT_REG = rnode_242to243_bb4_or2662_i164_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_or2662_i164_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4_or2662_i164_1_NO_SHIFT_REG = rnode_242to243_bb4_or2662_i164_0_reg_243_NO_SHIFT_REG;
assign rnode_242to243_bb4_or2662_i164_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_242to243_bb4_or2662_i164_2_NO_SHIFT_REG = rnode_242to243_bb4_or2662_i164_0_reg_243_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or275_i171_stall_local;
wire [31:0] local_bb4_or275_i171;

assign local_bb4_or275_i171 = ((local_bb4_or274_i170 & 32'h7FFFFFFF) | (rnode_242to243_bb4_resultSign_0_i151_0_NO_SHIFT_REG & 32'h80000000));

// This section implements an unregistered operation.
// 
wire local_bb4_var__u93_stall_local;
wire [31:0] local_bb4_var__u93;

assign local_bb4_var__u93[31:1] = 31'h0;
assign local_bb4_var__u93[0] = rnode_242to243_bb4__47_i161_1_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_or2804_i172_stall_local;
wire local_bb4_or2804_i172;

assign local_bb4_or2804_i172 = (rnode_242to243_bb4__47_i161_0_NO_SHIFT_REG | rnode_242to243_bb4_or2662_i164_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_or2875_i174_stall_local;
wire local_bb4_or2875_i174;

assign local_bb4_or2875_i174 = (rnode_242to243_bb4_or2662_i164_1_NO_SHIFT_REG | rnode_242to243_bb4__26_i49_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u94_stall_local;
wire [31:0] local_bb4_var__u94;

assign local_bb4_var__u94[31:1] = 31'h0;
assign local_bb4_var__u94[0] = rnode_242to243_bb4_or2662_i164_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext314_i188_stall_local;
wire [31:0] local_bb4_lnot_ext314_i188;

assign local_bb4_lnot_ext314_i188 = ((local_bb4_var__u93 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_cond282_i173_stall_local;
wire [31:0] local_bb4_cond282_i173;

assign local_bb4_cond282_i173 = (local_bb4_or2804_i172 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb4_cond289_i175_stall_local;
wire [31:0] local_bb4_cond289_i175;

assign local_bb4_cond289_i175 = (local_bb4_or2875_i174 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb4_lnot_ext310_i187_stall_local;
wire [31:0] local_bb4_lnot_ext310_i187;

assign local_bb4_lnot_ext310_i187 = ((local_bb4_var__u94 & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb4_and293_i177_stall_local;
wire [31:0] local_bb4_and293_i177;

assign local_bb4_and293_i177 = ((local_bb4_cond282_i173 | 32'h80000000) & local_bb4_or275_i171);

// This section implements an unregistered operation.
// 
wire local_bb4_or294_i178_stall_local;
wire [31:0] local_bb4_or294_i178;

assign local_bb4_or294_i178 = ((local_bb4_cond289_i175 & 32'h7F800000) | (local_bb4_cond292_i176 & 32'h400000));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_0_i189_stall_local;
wire [31:0] local_bb4_reduction_0_i189;

assign local_bb4_reduction_0_i189 = ((local_bb4_lnot_ext310_i187 & 32'h1) & (local_bb4_lnot_ext_i186 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_and302_i183_stall_local;
wire [31:0] local_bb4_and302_i183;

assign local_bb4_and302_i183 = ((local_bb4_conv300_i182 & 32'h1) & local_bb4_and293_i177);

// This section implements an unregistered operation.
// 
wire local_bb4_or295_i179_stall_local;
wire [31:0] local_bb4_or295_i179;

assign local_bb4_or295_i179 = ((local_bb4_or294_i178 & 32'h7FC00000) | local_bb4_and293_i177);

// This section implements an unregistered operation.
// 
wire local_bb4_lor_ext_i185_stall_local;
wire [31:0] local_bb4_lor_ext_i185;

assign local_bb4_lor_ext_i185 = ((local_bb4_cmp29649_i184 & 32'h1) | (local_bb4_and302_i183 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_1_i190_stall_local;
wire [31:0] local_bb4_reduction_1_i190;

assign local_bb4_reduction_1_i190 = ((local_bb4_lnot_ext314_i188 & 32'h1) & (local_bb4_lor_ext_i185 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_reduction_2_i191_stall_local;
wire [31:0] local_bb4_reduction_2_i191;

assign local_bb4_reduction_2_i191 = ((local_bb4_reduction_0_i189 & 32'h1) & (local_bb4_reduction_1_i190 & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb4_add320_i192_stall_local;
wire [31:0] local_bb4_add320_i192;

assign local_bb4_add320_i192 = ((local_bb4_reduction_2_i191 & 32'h1) + local_bb4_or295_i179);

// This section implements an unregistered operation.
// 
wire local_bb4_var__u95_stall_local;
wire [31:0] local_bb4_var__u95;

assign local_bb4_var__u95 = local_bb4_add320_i192;

// This section implements an unregistered operation.
// 
wire local_bb4__46_valid_out;
wire local_bb4__46_stall_in;
wire local_bb4__46_inputs_ready;
wire local_bb4__46_stall_local;
wire [31:0] local_bb4__46;

assign local_bb4__46_inputs_ready = (rnode_242to243_bb4_cmp34_0_valid_out_NO_SHIFT_REG & rnode_242to243_bb4_t_322_pop8_c1_ene3_0_valid_out_NO_SHIFT_REG & rnode_241to243_bb4_and269_i168_0_valid_out_NO_SHIFT_REG & rnode_242to243_bb4_resultSign_0_i151_0_valid_out_NO_SHIFT_REG & rnode_242to243_bb4_or2662_i164_0_valid_out_1_NO_SHIFT_REG & rnode_242to243_bb4__26_i49_0_valid_out_0_NO_SHIFT_REG & rnode_242to243_bb4__26_i49_0_valid_out_1_NO_SHIFT_REG & rnode_242to243_bb4__47_i161_0_valid_out_0_NO_SHIFT_REG & rnode_242to243_bb4_or2662_i164_0_valid_out_0_NO_SHIFT_REG & rnode_242to243_bb4__26_i49_0_valid_out_2_NO_SHIFT_REG & rnode_242to243_bb4_or2662_i164_0_valid_out_2_NO_SHIFT_REG & rnode_242to243_bb4_shr271_i166_0_valid_out_NO_SHIFT_REG & rnode_242to243_bb4__47_i161_0_valid_out_1_NO_SHIFT_REG & rnode_242to243_bb4_cmp296_i180_0_valid_out_NO_SHIFT_REG & rnode_242to243_bb4_cmp299_i181_0_valid_out_NO_SHIFT_REG);
assign local_bb4__46 = (rnode_242to243_bb4_cmp34_0_NO_SHIFT_REG ? local_bb4_var__u95 : rnode_242to243_bb4_t_322_pop8_c1_ene3_0_NO_SHIFT_REG);
assign local_bb4__46_valid_out = 1'b1;
assign rnode_242to243_bb4_cmp34_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_t_322_pop8_c1_ene3_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_241to243_bb4_and269_i168_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_resultSign_0_i151_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_or2662_i164_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__26_i49_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__26_i49_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__47_i161_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_or2662_i164_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__26_i49_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_or2662_i164_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_shr271_i166_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4__47_i161_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_cmp296_i180_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_242to243_bb4_cmp299_i181_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_243to244_bb4__46_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_243to244_bb4__46_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_243to244_bb4__46_0_NO_SHIFT_REG;
 logic rnode_243to244_bb4__46_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_243to244_bb4__46_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_243to244_bb4__46_1_NO_SHIFT_REG;
 logic rnode_243to244_bb4__46_0_reg_244_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_243to244_bb4__46_0_reg_244_NO_SHIFT_REG;
 logic rnode_243to244_bb4__46_0_valid_out_0_reg_244_NO_SHIFT_REG;
 logic rnode_243to244_bb4__46_0_stall_in_0_reg_244_NO_SHIFT_REG;
 logic rnode_243to244_bb4__46_0_stall_out_reg_244_NO_SHIFT_REG;

acl_data_fifo rnode_243to244_bb4__46_0_reg_244_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_243to244_bb4__46_0_reg_244_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_243to244_bb4__46_0_stall_in_0_reg_244_NO_SHIFT_REG),
	.valid_out(rnode_243to244_bb4__46_0_valid_out_0_reg_244_NO_SHIFT_REG),
	.stall_out(rnode_243to244_bb4__46_0_stall_out_reg_244_NO_SHIFT_REG),
	.data_in(local_bb4__46),
	.data_out(rnode_243to244_bb4__46_0_reg_244_NO_SHIFT_REG)
);

defparam rnode_243to244_bb4__46_0_reg_244_fifo.DEPTH = 1;
defparam rnode_243to244_bb4__46_0_reg_244_fifo.DATA_WIDTH = 32;
defparam rnode_243to244_bb4__46_0_reg_244_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_243to244_bb4__46_0_reg_244_fifo.IMPL = "shift_reg";

assign rnode_243to244_bb4__46_0_reg_244_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb4__46_stall_in = 1'b0;
assign rnode_243to244_bb4__46_0_stall_in_0_reg_244_NO_SHIFT_REG = 1'b0;
assign rnode_243to244_bb4__46_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_243to244_bb4__46_0_NO_SHIFT_REG = rnode_243to244_bb4__46_0_reg_244_NO_SHIFT_REG;
assign rnode_243to244_bb4__46_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_243to244_bb4__46_1_NO_SHIFT_REG = rnode_243to244_bb4__46_0_reg_244_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb4_t_322_push8__46_inputs_ready;
 reg local_bb4_t_322_push8__46_valid_out_NO_SHIFT_REG;
wire local_bb4_t_322_push8__46_stall_in;
wire local_bb4_t_322_push8__46_output_regs_ready;
wire [31:0] local_bb4_t_322_push8__46_result;
wire local_bb4_t_322_push8__46_fu_valid_out;
wire local_bb4_t_322_push8__46_fu_stall_out;
 reg [31:0] local_bb4_t_322_push8__46_NO_SHIFT_REG;
wire local_bb4_t_322_push8__46_causedstall;

acl_push local_bb4_t_322_push8__46_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(rnode_243to244_bb4_c1_ene6_0_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(rnode_243to244_bb4__46_0_NO_SHIFT_REG),
	.stall_out(local_bb4_t_322_push8__46_fu_stall_out),
	.valid_in(SFC_3_VALID_243_244_0_NO_SHIFT_REG),
	.valid_out(local_bb4_t_322_push8__46_fu_valid_out),
	.stall_in(1'b0),
	.data_out(local_bb4_t_322_push8__46_result),
	.feedback_out(feedback_data_out_8),
	.feedback_valid_out(feedback_valid_out_8),
	.feedback_stall_in(feedback_stall_in_8)
);

defparam local_bb4_t_322_push8__46_feedback.STALLFREE = 1;
defparam local_bb4_t_322_push8__46_feedback.DATA_WIDTH = 32;
defparam local_bb4_t_322_push8__46_feedback.FIFO_DEPTH = 9;
defparam local_bb4_t_322_push8__46_feedback.MIN_FIFO_LATENCY = 0;
defparam local_bb4_t_322_push8__46_feedback.STYLE = "REGULAR";

assign local_bb4_t_322_push8__46_inputs_ready = 1'b1;
assign local_bb4_t_322_push8__46_output_regs_ready = 1'b1;
assign SFC_3_VALID_243_244_0_stall_in_1 = 1'b0;
assign rnode_243to244_bb4__46_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_243to244_bb4_c1_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_t_322_push8__46_causedstall = (SFC_3_VALID_243_244_0_NO_SHIFT_REG && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_t_322_push8__46_NO_SHIFT_REG <= 'x;
		local_bb4_t_322_push8__46_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_t_322_push8__46_output_regs_ready)
		begin
			local_bb4_t_322_push8__46_NO_SHIFT_REG <= local_bb4_t_322_push8__46_result;
			local_bb4_t_322_push8__46_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb4_t_322_push8__46_stall_in))
			begin
				local_bb4_t_322_push8__46_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_244to245_bb4__46_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_244to245_bb4__46_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4__46_0_NO_SHIFT_REG;
 logic rnode_244to245_bb4__46_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_244to245_bb4__46_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4__46_1_NO_SHIFT_REG;
 logic rnode_244to245_bb4__46_0_reg_245_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_244to245_bb4__46_0_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4__46_0_valid_out_0_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4__46_0_stall_in_0_reg_245_NO_SHIFT_REG;
 logic rnode_244to245_bb4__46_0_stall_out_reg_245_NO_SHIFT_REG;

acl_data_fifo rnode_244to245_bb4__46_0_reg_245_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_244to245_bb4__46_0_reg_245_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_244to245_bb4__46_0_stall_in_0_reg_245_NO_SHIFT_REG),
	.valid_out(rnode_244to245_bb4__46_0_valid_out_0_reg_245_NO_SHIFT_REG),
	.stall_out(rnode_244to245_bb4__46_0_stall_out_reg_245_NO_SHIFT_REG),
	.data_in(rnode_243to244_bb4__46_1_NO_SHIFT_REG),
	.data_out(rnode_244to245_bb4__46_0_reg_245_NO_SHIFT_REG)
);

defparam rnode_244to245_bb4__46_0_reg_245_fifo.DEPTH = 1;
defparam rnode_244to245_bb4__46_0_reg_245_fifo.DATA_WIDTH = 32;
defparam rnode_244to245_bb4__46_0_reg_245_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_244to245_bb4__46_0_reg_245_fifo.IMPL = "shift_reg";

assign rnode_244to245_bb4__46_0_reg_245_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_243to244_bb4__46_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_244to245_bb4__46_0_stall_in_0_reg_245_NO_SHIFT_REG = 1'b0;
assign rnode_244to245_bb4__46_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_244to245_bb4__46_0_NO_SHIFT_REG = rnode_244to245_bb4__46_0_reg_245_NO_SHIFT_REG;
assign rnode_244to245_bb4__46_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_244to245_bb4__46_1_NO_SHIFT_REG = rnode_244to245_bb4__46_0_reg_245_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb4___46_valid_out;
wire local_bb4___46_stall_in;
wire local_bb4___46_inputs_ready;
wire local_bb4___46_stall_local;
 reg [31:0] ffwd_11_0_reg_NO_SHIFT_REG;

assign local_bb4___46_inputs_ready = (SFC_3_VALID_244_245_0_valid_out_2_NO_SHIFT_REG & rnode_244to245_bb4__46_0_valid_out_0_NO_SHIFT_REG);
assign ffwd_11_0 = ffwd_11_0_reg_NO_SHIFT_REG;
assign local_bb4___46_valid_out = 1'b1;
assign SFC_3_VALID_244_245_0_stall_in_2 = 1'b0;
assign rnode_244to245_bb4__46_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock)
begin
	if ((1'b1 & SFC_3_VALID_244_245_0_NO_SHIFT_REG))
	begin
		ffwd_11_0_reg_NO_SHIFT_REG <= rnode_244to245_bb4__46_0_NO_SHIFT_REG;
	end
end


// This section implements an unregistered operation.
// 
wire local_bb4_c1_exi2_valid_out;
wire local_bb4_c1_exi2_stall_in;
wire local_bb4_c1_exi2_inputs_ready;
wire local_bb4_c1_exi2_stall_local;
wire [95:0] local_bb4_c1_exi2;

assign local_bb4_c1_exi2_inputs_ready = (rnode_244to245_bb4__46_0_valid_out_1_NO_SHIFT_REG & rnode_244to245_bb4___0_valid_out_1_NO_SHIFT_REG);
assign local_bb4_c1_exi2[63:0] = local_bb4_c1_exi1[63:0];
assign local_bb4_c1_exi2[95:64] = rnode_244to245_bb4__46_1_NO_SHIFT_REG;
assign local_bb4_c1_exi2_valid_out = 1'b1;
assign rnode_244to245_bb4__46_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_244to245_bb4___0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb4_c1_exit_c1_exi2_inputs_ready;
 reg local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG;
wire local_bb4_c1_exit_c1_exi2_stall_in;
 reg [95:0] local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG;
wire [95:0] local_bb4_c1_exit_c1_exi2_in;
wire local_bb4_c1_exit_c1_exi2_valid;
wire local_bb4_c1_exit_c1_exi2_causedstall;

acl_stall_free_sink local_bb4_c1_exit_c1_exi2_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb4_c1_exi2),
	.data_out(local_bb4_c1_exit_c1_exi2_in),
	.input_accepted(local_bb4_c1_enter_c1_eni6_input_accepted),
	.valid_out(local_bb4_c1_exit_c1_exi2_valid),
	.stall_in(~(local_bb4_c1_exit_c1_exi2_output_regs_ready)),
	.stall_entry(local_bb4_c1_exit_c1_exi2_entry_stall),
	.valid_in(local_bb4_c1_exit_c1_exi2_valid_in),
	.IIphases(local_bb4_c1_exit_c1_exi2_phases),
	.inc_pipelined_thread(local_bb4_c1_enter_c1_eni6_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb4_c1_enter_c1_eni6_dec_pipelined_thread)
);

defparam local_bb4_c1_exit_c1_exi2_instance.DATA_WIDTH = 96;
defparam local_bb4_c1_exit_c1_exi2_instance.PIPELINE_DEPTH = 74;
defparam local_bb4_c1_exit_c1_exi2_instance.SHARINGII = 1;
defparam local_bb4_c1_exit_c1_exi2_instance.SCHEDULEII = 9;
defparam local_bb4_c1_exit_c1_exi2_instance.ALWAYS_THROTTLE = 0;

assign local_bb4_c1_exit_c1_exi2_inputs_ready = 1'b1;
assign local_bb4_c1_exit_c1_exi2_output_regs_ready = (&(~(local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG) | ~(local_bb4_c1_exit_c1_exi2_stall_in)));
assign local_bb4_c1_exit_c1_exi2_valid_in = SFC_3_VALID_244_245_0_NO_SHIFT_REG;
assign local_bb4_c1_exi2_stall_in = 1'b0;
assign local_bb4_t_322_push8__46_stall_in = 1'b0;
assign local_bb4____stall_in = 1'b0;
assign local_bb4___46_stall_in = 1'b0;
assign SFC_3_VALID_244_245_0_stall_in_0 = 1'b0;
assign rnode_244to245_bb4_sum_321_push9___0_stall_in_NO_SHIFT_REG = 1'b0;
assign local_bb4_c1_exit_c1_exi2_causedstall = (1'b1 && (1'b0 && !(~(local_bb4_c1_exit_c1_exi2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG <= 'x;
		local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb4_c1_exit_c1_exi2_output_regs_ready)
		begin
			local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_in;
			local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_valid;
		end
		else
		begin
			if (~(local_bb4_c1_exit_c1_exi2_stall_in))
			begin
				local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [191:0] lvb_bb4_c0_exit28_c0_exi6_0_reg_NO_SHIFT_REG;
 reg lvb_bb4_c0_exe6_0_reg_NO_SHIFT_REG;
 reg [95:0] lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb4_c1_exit_c1_exi2_valid_out_NO_SHIFT_REG & local_bb4_c0_exe6_valid_out & local_bb4_c0_exe331_valid_out & rnode_249to250_bb4_c0_exit28_c0_exi6_0_valid_out_2_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb4_c1_exit_c1_exi2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe6_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb4_c0_exe331_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_249to250_bb4_c0_exit28_c0_exi6_0_stall_in_2_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb4_c0_exit28_c0_exi6_0 = lvb_bb4_c0_exit28_c0_exi6_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exit28_c0_exi6_1 = lvb_bb4_c0_exit28_c0_exi6_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe6_0 = lvb_bb4_c0_exe6_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c0_exe6_1 = lvb_bb4_c0_exe6_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exit_c1_exi2_0 = lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG;
assign lvb_bb4_c1_exit_c1_exi2_1 = lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_bb4_c0_exit28_c0_exi6_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c0_exe6_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb4_c0_exit28_c0_exi6_0_reg_NO_SHIFT_REG <= rnode_249to250_bb4_c0_exit28_c0_exi6_2_NO_SHIFT_REG;
			lvb_bb4_c0_exe6_0_reg_NO_SHIFT_REG <= local_bb4_c0_exe6;
			lvb_bb4_c1_exit_c1_exi2_0_reg_NO_SHIFT_REG <= local_bb4_c1_exit_c1_exi2_NO_SHIFT_REG;
			branch_compare_result_NO_SHIFT_REG <= local_bb4_c0_exe331;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_5
	(
		input 		clock,
		input 		resetn,
		input 		input_wii_cmp1526,
		input [31:0] 		input_wii_sub24,
		input [31:0] 		input_wii_sub27,
		input [31:0] 		input_wii_mul48,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u96,
		input 		valid_in,
		output 		stall_out,
		input [191:0] 		input_c0_exit28_c0_exi6,
		input 		input_c0_exe6,
		input [95:0] 		input_c1_exit_c1_exi2,
		output 		valid_out_0,
		input 		stall_in_0,
		output 		valid_out_1,
		input 		stall_in_1,
		input [31:0] 		workgroup_size,
		input 		start,
		output 		feedback_valid_out_5,
		input 		feedback_stall_in_5,
		output [31:0] 		feedback_data_out_5,
		output 		feedback_valid_out_6,
		input 		feedback_stall_in_6,
		output [31:0] 		feedback_data_out_6
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [191:0] input_c0_exit28_c0_exi6_staging_reg_NO_SHIFT_REG;
 reg input_c0_exe6_staging_reg_NO_SHIFT_REG;
 reg [95:0] input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG;
 reg [191:0] local_lvm_c0_exit28_c0_exi6_NO_SHIFT_REG;
 reg local_lvm_c0_exe6_NO_SHIFT_REG;
 reg [95:0] local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_c0_exit28_c0_exi6_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe6_staging_reg_NO_SHIFT_REG <= 'x;
		input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_c0_exit28_c0_exi6_staging_reg_NO_SHIFT_REG <= input_c0_exit28_c0_exi6;
				input_c0_exe6_staging_reg_NO_SHIFT_REG <= input_c0_exe6;
				input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG <= input_c1_exit_c1_exi2;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_c0_exit28_c0_exi6_NO_SHIFT_REG <= input_c0_exit28_c0_exi6_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe6_NO_SHIFT_REG <= input_c0_exe6_staging_reg_NO_SHIFT_REG;
					local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG <= input_c1_exit_c1_exi2_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_c0_exit28_c0_exi6_NO_SHIFT_REG <= input_c0_exit28_c0_exi6;
					local_lvm_c0_exe6_NO_SHIFT_REG <= input_c0_exe6;
					local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG <= input_c1_exit_c1_exi2;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb5_c1_exe2_valid_out;
wire local_bb5_c1_exe2_stall_in;
wire local_bb5_c1_exe2_inputs_ready;
wire local_bb5_c1_exe2_stall_local;
wire [31:0] local_bb5_c1_exe2;

assign local_bb5_c1_exe2_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb5_c1_exe2 = local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG[95:64];
assign local_bb5_c1_exe2_valid_out = local_bb5_c1_exe2_inputs_ready;
assign local_bb5_c1_exe2_stall_local = local_bb5_c1_exe2_stall_in;
assign merge_node_stall_in_0 = (|local_bb5_c1_exe2_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb5_c1_exe1_valid_out;
wire local_bb5_c1_exe1_stall_in;
wire local_bb5_c1_exe1_inputs_ready;
wire local_bb5_c1_exe1_stall_local;
wire [31:0] local_bb5_c1_exe1;

assign local_bb5_c1_exe1_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb5_c1_exe1 = local_lvm_c1_exit_c1_exi2_NO_SHIFT_REG[63:32];
assign local_bb5_c1_exe1_valid_out = local_bb5_c1_exe1_inputs_ready;
assign local_bb5_c1_exe1_stall_local = local_bb5_c1_exe1_stall_in;
assign merge_node_stall_in_1 = (|local_bb5_c1_exe1_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb5_c0_exe5_valid_out;
wire local_bb5_c0_exe5_stall_in;
wire local_bb5_c0_exe5_inputs_ready;
wire local_bb5_c0_exe5_stall_local;
wire local_bb5_c0_exe5;

assign local_bb5_c0_exe5_inputs_ready = merge_node_valid_out_2_NO_SHIFT_REG;
assign local_bb5_c0_exe5 = local_lvm_c0_exit28_c0_exi6_NO_SHIFT_REG[176];
assign local_bb5_c0_exe5_valid_out = local_bb5_c0_exe5_inputs_ready;
assign local_bb5_c0_exe5_stall_local = local_bb5_c0_exe5_stall_in;
assign merge_node_stall_in_2 = (|local_bb5_c0_exe5_stall_local);

// This section implements a registered operation.
// 
wire local_bb5_t_228_push5_c1_exe2_inputs_ready;
 reg local_bb5_t_228_push5_c1_exe2_valid_out_NO_SHIFT_REG;
wire local_bb5_t_228_push5_c1_exe2_stall_in;
wire local_bb5_t_228_push5_c1_exe2_output_regs_ready;
wire [31:0] local_bb5_t_228_push5_c1_exe2_result;
wire local_bb5_t_228_push5_c1_exe2_fu_valid_out;
wire local_bb5_t_228_push5_c1_exe2_fu_stall_out;
 reg [31:0] local_bb5_t_228_push5_c1_exe2_NO_SHIFT_REG;
wire local_bb5_t_228_push5_c1_exe2_causedstall;

acl_push local_bb5_t_228_push5_c1_exe2_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_c0_exe6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb5_c1_exe2),
	.stall_out(local_bb5_t_228_push5_c1_exe2_fu_stall_out),
	.valid_in(local_bb5_t_228_push5_c1_exe2_inputs_ready),
	.valid_out(local_bb5_t_228_push5_c1_exe2_fu_valid_out),
	.stall_in(~(local_bb5_t_228_push5_c1_exe2_output_regs_ready)),
	.data_out(local_bb5_t_228_push5_c1_exe2_result),
	.feedback_out(feedback_data_out_5),
	.feedback_valid_out(feedback_valid_out_5),
	.feedback_stall_in(feedback_stall_in_5)
);

defparam local_bb5_t_228_push5_c1_exe2_feedback.STALLFREE = 0;
defparam local_bb5_t_228_push5_c1_exe2_feedback.DATA_WIDTH = 32;
defparam local_bb5_t_228_push5_c1_exe2_feedback.FIFO_DEPTH = 3;
defparam local_bb5_t_228_push5_c1_exe2_feedback.MIN_FIFO_LATENCY = 3;
defparam local_bb5_t_228_push5_c1_exe2_feedback.STYLE = "REGULAR";

assign local_bb5_t_228_push5_c1_exe2_inputs_ready = (local_bb5_c1_exe2_valid_out & merge_node_valid_out_4_NO_SHIFT_REG);
assign local_bb5_t_228_push5_c1_exe2_output_regs_ready = (&(~(local_bb5_t_228_push5_c1_exe2_valid_out_NO_SHIFT_REG) | ~(local_bb5_t_228_push5_c1_exe2_stall_in)));
assign local_bb5_c1_exe2_stall_in = (local_bb5_t_228_push5_c1_exe2_fu_stall_out | ~(local_bb5_t_228_push5_c1_exe2_inputs_ready));
assign merge_node_stall_in_4 = (local_bb5_t_228_push5_c1_exe2_fu_stall_out | ~(local_bb5_t_228_push5_c1_exe2_inputs_ready));
assign local_bb5_t_228_push5_c1_exe2_causedstall = (local_bb5_t_228_push5_c1_exe2_inputs_ready && (local_bb5_t_228_push5_c1_exe2_fu_stall_out && !(~(local_bb5_t_228_push5_c1_exe2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_t_228_push5_c1_exe2_NO_SHIFT_REG <= 'x;
		local_bb5_t_228_push5_c1_exe2_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_t_228_push5_c1_exe2_output_regs_ready)
		begin
			local_bb5_t_228_push5_c1_exe2_NO_SHIFT_REG <= local_bb5_t_228_push5_c1_exe2_result;
			local_bb5_t_228_push5_c1_exe2_valid_out_NO_SHIFT_REG <= local_bb5_t_228_push5_c1_exe2_fu_valid_out;
		end
		else
		begin
			if (~(local_bb5_t_228_push5_c1_exe2_stall_in))
			begin
				local_bb5_t_228_push5_c1_exe2_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb5_sum_227_push6_c1_exe1_inputs_ready;
 reg local_bb5_sum_227_push6_c1_exe1_valid_out_NO_SHIFT_REG;
wire local_bb5_sum_227_push6_c1_exe1_stall_in;
wire local_bb5_sum_227_push6_c1_exe1_output_regs_ready;
wire [31:0] local_bb5_sum_227_push6_c1_exe1_result;
wire local_bb5_sum_227_push6_c1_exe1_fu_valid_out;
wire local_bb5_sum_227_push6_c1_exe1_fu_stall_out;
 reg [31:0] local_bb5_sum_227_push6_c1_exe1_NO_SHIFT_REG;
wire local_bb5_sum_227_push6_c1_exe1_causedstall;

acl_push local_bb5_sum_227_push6_c1_exe1_feedback (
	.clock(clock),
	.resetn(resetn),
	.dir(local_lvm_c0_exe6_NO_SHIFT_REG),
	.predicate(1'b0),
	.data_in(local_bb5_c1_exe1),
	.stall_out(local_bb5_sum_227_push6_c1_exe1_fu_stall_out),
	.valid_in(local_bb5_sum_227_push6_c1_exe1_inputs_ready),
	.valid_out(local_bb5_sum_227_push6_c1_exe1_fu_valid_out),
	.stall_in(~(local_bb5_sum_227_push6_c1_exe1_output_regs_ready)),
	.data_out(local_bb5_sum_227_push6_c1_exe1_result),
	.feedback_out(feedback_data_out_6),
	.feedback_valid_out(feedback_valid_out_6),
	.feedback_stall_in(feedback_stall_in_6)
);

defparam local_bb5_sum_227_push6_c1_exe1_feedback.STALLFREE = 0;
defparam local_bb5_sum_227_push6_c1_exe1_feedback.DATA_WIDTH = 32;
defparam local_bb5_sum_227_push6_c1_exe1_feedback.FIFO_DEPTH = 3;
defparam local_bb5_sum_227_push6_c1_exe1_feedback.MIN_FIFO_LATENCY = 3;
defparam local_bb5_sum_227_push6_c1_exe1_feedback.STYLE = "REGULAR";

assign local_bb5_sum_227_push6_c1_exe1_inputs_ready = (local_bb5_c1_exe1_valid_out & merge_node_valid_out_3_NO_SHIFT_REG);
assign local_bb5_sum_227_push6_c1_exe1_output_regs_ready = (&(~(local_bb5_sum_227_push6_c1_exe1_valid_out_NO_SHIFT_REG) | ~(local_bb5_sum_227_push6_c1_exe1_stall_in)));
assign local_bb5_c1_exe1_stall_in = (local_bb5_sum_227_push6_c1_exe1_fu_stall_out | ~(local_bb5_sum_227_push6_c1_exe1_inputs_ready));
assign merge_node_stall_in_3 = (local_bb5_sum_227_push6_c1_exe1_fu_stall_out | ~(local_bb5_sum_227_push6_c1_exe1_inputs_ready));
assign local_bb5_sum_227_push6_c1_exe1_causedstall = (local_bb5_sum_227_push6_c1_exe1_inputs_ready && (local_bb5_sum_227_push6_c1_exe1_fu_stall_out && !(~(local_bb5_sum_227_push6_c1_exe1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb5_sum_227_push6_c1_exe1_NO_SHIFT_REG <= 'x;
		local_bb5_sum_227_push6_c1_exe1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb5_sum_227_push6_c1_exe1_output_regs_ready)
		begin
			local_bb5_sum_227_push6_c1_exe1_NO_SHIFT_REG <= local_bb5_sum_227_push6_c1_exe1_result;
			local_bb5_sum_227_push6_c1_exe1_valid_out_NO_SHIFT_REG <= local_bb5_sum_227_push6_c1_exe1_fu_valid_out;
		end
		else
		begin
			if (~(local_bb5_sum_227_push6_c1_exe1_stall_in))
			begin
				local_bb5_sum_227_push6_c1_exe1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_1to2_bb5_c0_exe5_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe5_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe5_0_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe5_0_reg_2_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe5_0_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe5_0_valid_out_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe5_0_stall_in_reg_2_NO_SHIFT_REG;
 logic rnode_1to2_bb5_c0_exe5_0_stall_out_reg_2_NO_SHIFT_REG;

acl_data_fifo rnode_1to2_bb5_c0_exe5_0_reg_2_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to2_bb5_c0_exe5_0_reg_2_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to2_bb5_c0_exe5_0_stall_in_reg_2_NO_SHIFT_REG),
	.valid_out(rnode_1to2_bb5_c0_exe5_0_valid_out_reg_2_NO_SHIFT_REG),
	.stall_out(rnode_1to2_bb5_c0_exe5_0_stall_out_reg_2_NO_SHIFT_REG),
	.data_in(local_bb5_c0_exe5),
	.data_out(rnode_1to2_bb5_c0_exe5_0_reg_2_NO_SHIFT_REG)
);

defparam rnode_1to2_bb5_c0_exe5_0_reg_2_fifo.DEPTH = 1;
defparam rnode_1to2_bb5_c0_exe5_0_reg_2_fifo.DATA_WIDTH = 1;
defparam rnode_1to2_bb5_c0_exe5_0_reg_2_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_1to2_bb5_c0_exe5_0_reg_2_fifo.IMPL = "ll_reg";

assign rnode_1to2_bb5_c0_exe5_0_reg_2_inputs_ready_NO_SHIFT_REG = local_bb5_c0_exe5_valid_out;
assign local_bb5_c0_exe5_stall_in = rnode_1to2_bb5_c0_exe5_0_stall_out_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb5_c0_exe5_0_NO_SHIFT_REG = rnode_1to2_bb5_c0_exe5_0_reg_2_NO_SHIFT_REG;
assign rnode_1to2_bb5_c0_exe5_0_stall_in_reg_2_NO_SHIFT_REG = rnode_1to2_bb5_c0_exe5_0_stall_in_NO_SHIFT_REG;
assign rnode_1to2_bb5_c0_exe5_0_valid_out_NO_SHIFT_REG = rnode_1to2_bb5_c0_exe5_0_valid_out_reg_2_NO_SHIFT_REG;

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;

assign branch_var__inputs_ready = (local_bb5_t_228_push5_c1_exe2_valid_out_NO_SHIFT_REG & local_bb5_sum_227_push6_c1_exe1_valid_out_NO_SHIFT_REG & rnode_1to2_bb5_c0_exe5_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb5_t_228_push5_c1_exe2_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb5_sum_227_push6_c1_exe1_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to2_bb5_c0_exe5_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			branch_compare_result_NO_SHIFT_REG <= rnode_1to2_bb5_c0_exe5_0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_6
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_out,
		input 		input_wii_cmp1526,
		input [31:0] 		input_wii_sub24,
		input [31:0] 		input_wii_sub27,
		input [31:0] 		input_wii_mul48,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u97,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out_0,
		input 		stall_in_0,
		output [63:0] 		lvb_bb6_indvars_iv_next40_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [63:0] 		lvb_bb6_indvars_iv_next40_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		ffwd_9_0,
		input 		ffwd_5_0,
		input [31:0] 		ffwd_11_0,
		input [31:0] 		ffwd_10_0,
		input [63:0] 		ffwd_6_0,
		input [63:0] 		ffwd_3_0,
		input 		ffwd_8_0,
		output [63:0] 		ffwd_12_0,
		input [511:0] 		avm_local_bb6_st_c0_exe239_readdata,
		input 		avm_local_bb6_st_c0_exe239_readdatavalid,
		input 		avm_local_bb6_st_c0_exe239_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe239_address,
		output 		avm_local_bb6_st_c0_exe239_read,
		output 		avm_local_bb6_st_c0_exe239_write,
		input 		avm_local_bb6_st_c0_exe239_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe239_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe239_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe239_burstcount,
		output 		local_bb6_st_c0_exe239_active,
		input 		clock2x
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb6_c0_enter33__inputs_ready;
 reg local_bb6_c0_enter33__valid_out_0_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_0;
 reg local_bb6_c0_enter33__valid_out_1_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_1;
 reg local_bb6_c0_enter33__valid_out_2_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_2;
 reg local_bb6_c0_enter33__valid_out_3_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_3;
 reg local_bb6_c0_enter33__valid_out_4_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_4;
 reg local_bb6_c0_enter33__valid_out_5_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_5;
 reg local_bb6_c0_enter33__valid_out_6_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_6;
 reg local_bb6_c0_enter33__valid_out_7_NO_SHIFT_REG;
wire local_bb6_c0_enter33__stall_in_7;
wire local_bb6_c0_enter33__output_regs_ready;
 reg [7:0] local_bb6_c0_enter33__NO_SHIFT_REG;
wire local_bb6_c0_enter33__input_accepted;
 reg local_bb6_c0_enter33__valid_bit_NO_SHIFT_REG;
wire local_bb6_c0_exit37_c0_exi336_entry_stall;
wire local_bb6_c0_exit37_c0_exi336_output_regs_ready;
wire [15:0] local_bb6_c0_exit37_c0_exi336_valid_bits;
wire local_bb6_c0_exit37_c0_exi336_valid_in;
wire local_bb6_c0_exit37_c0_exi336_phases;
wire local_bb6_c0_enter33__inc_pipelined_thread;
wire local_bb6_c0_enter33__dec_pipelined_thread;
wire local_bb6_c0_enter33__causedstall;

assign local_bb6_c0_enter33__inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb6_c0_enter33__output_regs_ready = 1'b1;
assign local_bb6_c0_enter33__input_accepted = (local_bb6_c0_enter33__inputs_ready && !(local_bb6_c0_exit37_c0_exi336_entry_stall));
assign local_bb6_c0_enter33__inc_pipelined_thread = 1'b1;
assign local_bb6_c0_enter33__dec_pipelined_thread = ~(1'b0);
assign merge_node_stall_in_0 = ((~(local_bb6_c0_enter33__inputs_ready) | local_bb6_c0_exit37_c0_exi336_entry_stall) | ~(1'b1));
assign local_bb6_c0_enter33__causedstall = (1'b1 && ((~(local_bb6_c0_enter33__inputs_ready) | local_bb6_c0_exit37_c0_exi336_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_enter33__valid_bit_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb6_c0_enter33__valid_bit_NO_SHIFT_REG <= local_bb6_c0_enter33__input_accepted;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_enter33__NO_SHIFT_REG <= 'x;
		local_bb6_c0_enter33__valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter33__valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter33__valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter33__valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter33__valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter33__valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter33__valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_enter33__valid_out_7_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_c0_enter33__output_regs_ready)
		begin
			local_bb6_c0_enter33__NO_SHIFT_REG <= 'x;
			local_bb6_c0_enter33__valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter33__valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter33__valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter33__valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter33__valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter33__valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter33__valid_out_6_NO_SHIFT_REG <= 1'b1;
			local_bb6_c0_enter33__valid_out_7_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb6_c0_enter33__stall_in_0))
			begin
				local_bb6_c0_enter33__valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter33__stall_in_1))
			begin
				local_bb6_c0_enter33__valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter33__stall_in_2))
			begin
				local_bb6_c0_enter33__valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter33__stall_in_3))
			begin
				local_bb6_c0_enter33__valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter33__stall_in_4))
			begin
				local_bb6_c0_enter33__valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter33__stall_in_5))
			begin
				local_bb6_c0_enter33__valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter33__stall_in_6))
			begin
				local_bb6_c0_enter33__valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_enter33__stall_in_7))
			begin
				local_bb6_c0_enter33__valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 18
//  * capacity = 18
 logic rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_reg_19_NO_SHIFT_REG;
 logic rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_reg_19_NO_SHIFT_REG;
 logic rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_out_reg_19_NO_SHIFT_REG;

acl_data_fifo rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_reg_19_NO_SHIFT_REG),
	.valid_out(rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_reg_19_NO_SHIFT_REG),
	.stall_out(rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_out_reg_19_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_fifo.DEPTH = 19;
defparam rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_fifo.DATA_WIDTH = 0;
defparam rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_fifo.IMPL = "ram";

assign rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_19_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign merge_node_stall_in_1 = rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_out_reg_19_NO_SHIFT_REG;
assign rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_reg_19_NO_SHIFT_REG = rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_NO_SHIFT_REG;
assign rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_NO_SHIFT_REG = rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_reg_19_NO_SHIFT_REG;

// Register node:
//  * latency = 179
//  * capacity = 179
 logic rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_fifo.DEPTH = 180;
defparam rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_fifo.DATA_WIDTH = 0;
defparam rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_fifo.IMPL = "ram";

assign rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_180_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign merge_node_stall_in_2 = rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_out_reg_180_NO_SHIFT_REG;
assign rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_reg_180_NO_SHIFT_REG = rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_NO_SHIFT_REG;
assign rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_NO_SHIFT_REG = rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_9_stall_local;
wire local_bb6__acl_ffwd_dest_i1_9;

assign local_bb6__acl_ffwd_dest_i1_9 = ffwd_9_0;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_5_stall_local;
wire local_bb6__acl_ffwd_dest_i1_5;

assign local_bb6__acl_ffwd_dest_i1_5 = ffwd_5_0;

// This section implements an unregistered operation.
// 
wire local_bb6__4610_acl_ffwd_dest_f_11_stall_local;
wire [31:0] local_bb6__4610_acl_ffwd_dest_f_11;

assign local_bb6__4610_acl_ffwd_dest_f_11 = ffwd_11_0;

// This section implements an unregistered operation.
// 
wire local_bb6__9_acl_ffwd_dest_f_10_stall_local;
wire [31:0] local_bb6__9_acl_ffwd_dest_f_10;

assign local_bb6__9_acl_ffwd_dest_f_10 = ffwd_10_0;

// This section implements an unregistered operation.
// 
wire SFC_4_VALID_2_2_0_valid_out;
wire SFC_4_VALID_2_2_0_stall_in;
wire SFC_4_VALID_2_2_0_inputs_ready;
wire SFC_4_VALID_2_2_0_stall_local;
wire SFC_4_VALID_2_2_0;

assign SFC_4_VALID_2_2_0_inputs_ready = local_bb6_c0_enter33__valid_out_4_NO_SHIFT_REG;
assign SFC_4_VALID_2_2_0 = local_bb6_c0_enter33__valid_bit_NO_SHIFT_REG;
assign SFC_4_VALID_2_2_0_valid_out = 1'b1;
assign local_bb6_c0_enter33__stall_in_4 = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_c0_enter33__stall_in_5 = 1'b0;
assign rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_c0_enter33__stall_in_6 = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_fifo.DATA_WIDTH = 0;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_c0_enter33__stall_in_7 = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_NO_SHIFT_REG;
 logic rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_NO_SHIFT_REG;
 logic rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_inputs_ready_NO_SHIFT_REG;
 logic rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_reg_20_NO_SHIFT_REG;
 logic rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_reg_20_NO_SHIFT_REG;
 logic rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_out_reg_20_NO_SHIFT_REG;

acl_data_fifo rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_reg_20_NO_SHIFT_REG),
	.valid_out(rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_reg_20_NO_SHIFT_REG),
	.stall_out(rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_out_reg_20_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_fifo.DEPTH = 1;
defparam rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_fifo.DATA_WIDTH = 0;
defparam rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_fifo.IMPL = "ll_reg";

assign rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_reg_20_inputs_ready_NO_SHIFT_REG = rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_NO_SHIFT_REG;
assign rnode_1to19_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_NO_SHIFT_REG = rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_out_reg_20_NO_SHIFT_REG;
assign rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_reg_20_NO_SHIFT_REG = rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_NO_SHIFT_REG;
assign rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_NO_SHIFT_REG = rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_reg_20_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_fifo.DATA_WIDTH = 0;
defparam rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_fifo.IMPL = "ll_reg";

assign rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_reg_181_inputs_ready_NO_SHIFT_REG = rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_NO_SHIFT_REG;
assign rnode_1to180_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_NO_SHIFT_REG = rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_out_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_reg_181_NO_SHIFT_REG = rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_NO_SHIFT_REG;
assign rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_NO_SHIFT_REG = rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_reg_181_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end57_loopexit_select97_stall_local;
wire local_bb6_do_directly_for_end57_loopexit_select97;

assign local_bb6_do_directly_for_end57_loopexit_select97 = (local_bb6__acl_ffwd_dest_i1_9 ^ 1'b1);

// This section implements a registered operation.
// 
wire SFC_4_VALID_2_3_0_inputs_ready;
 reg SFC_4_VALID_2_3_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_2_3_0_stall_in;
wire SFC_4_VALID_2_3_0_output_regs_ready;
 reg SFC_4_VALID_2_3_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_2_3_0_causedstall;

assign SFC_4_VALID_2_3_0_inputs_ready = 1'b1;
assign SFC_4_VALID_2_3_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_2_2_0_stall_in = 1'b0;
assign SFC_4_VALID_2_3_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_2_3_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_2_3_0_output_regs_ready)
		begin
			SFC_4_VALID_2_3_0_NO_SHIFT_REG <= SFC_4_VALID_2_2_0;
		end
	end
end


// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_fifo.DATA_WIDTH = 0;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb6_idxprom7_acl_ffwd_dest_i64_6_stall_local;
wire [63:0] local_bb6_idxprom7_acl_ffwd_dest_i64_6;

assign local_bb6_idxprom7_acl_ffwd_dest_i64_6 = ffwd_6_0;

// This section implements an unregistered operation.
// 
wire local_bb6_indvars_iv396_acl_ffwd_dest_i64_3_stall_local;
wire [63:0] local_bb6_indvars_iv396_acl_ffwd_dest_i64_3;

assign local_bb6_indvars_iv396_acl_ffwd_dest_i64_3 = ffwd_3_0;

// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end57_loopexit_select_stall_local;
wire local_bb6_do_directly_for_end57_loopexit_select;

assign local_bb6_do_directly_for_end57_loopexit_select = (local_bb6__acl_ffwd_dest_i1_5 & local_bb6_do_directly_for_end57_loopexit_select97);

// This section implements a registered operation.
// 
wire SFC_4_VALID_3_4_0_inputs_ready;
 reg SFC_4_VALID_3_4_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_3_4_0_stall_in;
wire SFC_4_VALID_3_4_0_output_regs_ready;
 reg SFC_4_VALID_3_4_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_3_4_0_causedstall;

assign SFC_4_VALID_3_4_0_inputs_ready = 1'b1;
assign SFC_4_VALID_3_4_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_2_3_0_stall_in = 1'b0;
assign SFC_4_VALID_3_4_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_3_4_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_3_4_0_output_regs_ready)
		begin
			SFC_4_VALID_3_4_0_NO_SHIFT_REG <= SFC_4_VALID_2_3_0_NO_SHIFT_REG;
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_fifo.DATA_WIDTH = 0;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb6_arrayidx62_valid_out;
wire local_bb6_arrayidx62_stall_in;
wire local_bb6_arrayidx62_inputs_ready;
wire local_bb6_arrayidx62_stall_local;
wire [63:0] local_bb6_arrayidx62;

assign local_bb6_arrayidx62_inputs_ready = rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_valid_out_NO_SHIFT_REG;
assign local_bb6_arrayidx62 = ((input_out & 64'hFFFFFFFFFFFFFC00) + (local_bb6_idxprom7_acl_ffwd_dest_i64_6 << 6'h2));
assign local_bb6_arrayidx62_valid_out = local_bb6_arrayidx62_inputs_ready;
assign local_bb6_arrayidx62_stall_local = local_bb6_arrayidx62_stall_in;
assign rnode_19to20_bb6_idxprom7_acl_ffwd_dest_i64_6_0_stall_in_NO_SHIFT_REG = (|local_bb6_arrayidx62_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_indvars_iv_next40_valid_out;
wire local_bb6_indvars_iv_next40_stall_in;
wire local_bb6_indvars_iv_next40_inputs_ready;
wire local_bb6_indvars_iv_next40_stall_local;
wire [63:0] local_bb6_indvars_iv_next40;

assign local_bb6_indvars_iv_next40_inputs_ready = rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_valid_out_NO_SHIFT_REG;
assign local_bb6_indvars_iv_next40 = (local_bb6_indvars_iv396_acl_ffwd_dest_i64_3 + 64'h1);
assign local_bb6_indvars_iv_next40_valid_out = local_bb6_indvars_iv_next40_inputs_ready;
assign local_bb6_indvars_iv_next40_stall_local = local_bb6_indvars_iv_next40_stall_in;
assign rnode_180to181_bb6_indvars_iv396_acl_ffwd_dest_i64_3_0_stall_in_NO_SHIFT_REG = (|local_bb6_indvars_iv_next40_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_select78_stall_local;
wire [31:0] local_bb6_select78;

assign local_bb6_select78 = (local_bb6_do_directly_for_end57_loopexit_select ? local_bb6__4610_acl_ffwd_dest_f_11 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end57_loopexit_select_valid_out_2;
wire local_bb6_do_directly_for_end57_loopexit_select_stall_in_2;
wire local_bb6_select78_valid_out;
wire local_bb6_select78_stall_in;
wire local_bb6_select81_valid_out;
wire local_bb6_select81_stall_in;
wire local_bb6_select81_inputs_ready;
wire local_bb6_select81_stall_local;
wire [31:0] local_bb6_select81;

assign local_bb6_select81_inputs_ready = (local_bb6_c0_enter33__valid_out_0_NO_SHIFT_REG & local_bb6_c0_enter33__valid_out_1_NO_SHIFT_REG & local_bb6_c0_enter33__valid_out_2_NO_SHIFT_REG & local_bb6_c0_enter33__valid_out_3_NO_SHIFT_REG);
assign local_bb6_select81 = (local_bb6_do_directly_for_end57_loopexit_select ? local_bb6__9_acl_ffwd_dest_f_10 : 32'h0);
assign local_bb6_do_directly_for_end57_loopexit_select_valid_out_2 = 1'b1;
assign local_bb6_select78_valid_out = 1'b1;
assign local_bb6_select81_valid_out = 1'b1;
assign local_bb6_c0_enter33__stall_in_0 = 1'b0;
assign local_bb6_c0_enter33__stall_in_1 = 1'b0;
assign local_bb6_c0_enter33__stall_in_2 = 1'b0;
assign local_bb6_c0_enter33__stall_in_3 = 1'b0;

// This section implements a registered operation.
// 
wire SFC_4_VALID_4_5_0_inputs_ready;
 reg SFC_4_VALID_4_5_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_4_5_0_stall_in;
wire SFC_4_VALID_4_5_0_output_regs_ready;
 reg SFC_4_VALID_4_5_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_4_5_0_causedstall;

assign SFC_4_VALID_4_5_0_inputs_ready = 1'b1;
assign SFC_4_VALID_4_5_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_3_4_0_stall_in = 1'b0;
assign SFC_4_VALID_4_5_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_4_5_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_4_5_0_output_regs_ready)
		begin
			SFC_4_VALID_4_5_0_NO_SHIFT_REG <= SFC_4_VALID_3_4_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_cmp88_acl_ffwd_dest_i1_8_stall_local;
wire local_bb6_cmp88_acl_ffwd_dest_i1_8;

assign local_bb6_cmp88_acl_ffwd_dest_i1_8 = ffwd_8_0;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_5_u98_stall_local;
wire local_bb6__acl_ffwd_dest_i1_5_u98;

assign local_bb6__acl_ffwd_dest_i1_5_u98 = ffwd_5_0;

// This section implements an unregistered operation.
// 
wire local_bb6__acl_ffwd_dest_i1_9_u99_stall_local;
wire local_bb6__acl_ffwd_dest_i1_9_u99;

assign local_bb6__acl_ffwd_dest_i1_9_u99 = ffwd_9_0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_20to21_bb6_arrayidx62_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx62_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx62_0_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx62_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx62_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx62_1_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx62_0_reg_21_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_20to21_bb6_arrayidx62_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx62_0_valid_out_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx62_0_stall_in_0_reg_21_NO_SHIFT_REG;
 logic rnode_20to21_bb6_arrayidx62_0_stall_out_reg_21_NO_SHIFT_REG;
 reg rnode_20to21_bb6_arrayidx62_0_consumed_0_NO_SHIFT_REG;
 reg rnode_20to21_bb6_arrayidx62_0_consumed_1_NO_SHIFT_REG;

acl_data_fifo rnode_20to21_bb6_arrayidx62_0_reg_21_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_20to21_bb6_arrayidx62_0_reg_21_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_20to21_bb6_arrayidx62_0_stall_in_0_reg_21_NO_SHIFT_REG),
	.valid_out(rnode_20to21_bb6_arrayidx62_0_valid_out_0_reg_21_NO_SHIFT_REG),
	.stall_out(rnode_20to21_bb6_arrayidx62_0_stall_out_reg_21_NO_SHIFT_REG),
	.data_in((local_bb6_arrayidx62 & 64'hFFFFFFFFFFFFFFFC)),
	.data_out(rnode_20to21_bb6_arrayidx62_0_reg_21_NO_SHIFT_REG)
);

defparam rnode_20to21_bb6_arrayidx62_0_reg_21_fifo.DEPTH = 2;
defparam rnode_20to21_bb6_arrayidx62_0_reg_21_fifo.DATA_WIDTH = 64;
defparam rnode_20to21_bb6_arrayidx62_0_reg_21_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_20to21_bb6_arrayidx62_0_reg_21_fifo.IMPL = "ll_reg";

assign rnode_20to21_bb6_arrayidx62_0_reg_21_inputs_ready_NO_SHIFT_REG = local_bb6_arrayidx62_valid_out;
assign local_bb6_arrayidx62_stall_in = rnode_20to21_bb6_arrayidx62_0_stall_out_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb6_arrayidx62_0_stall_in_0_reg_21_NO_SHIFT_REG = ((rnode_20to21_bb6_arrayidx62_0_stall_in_0_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx62_0_consumed_0_NO_SHIFT_REG)) | (rnode_20to21_bb6_arrayidx62_0_stall_in_1_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx62_0_consumed_1_NO_SHIFT_REG)));
assign rnode_20to21_bb6_arrayidx62_0_valid_out_0_NO_SHIFT_REG = (rnode_20to21_bb6_arrayidx62_0_valid_out_0_reg_21_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx62_0_consumed_0_NO_SHIFT_REG));
assign rnode_20to21_bb6_arrayidx62_0_valid_out_1_NO_SHIFT_REG = (rnode_20to21_bb6_arrayidx62_0_valid_out_0_reg_21_NO_SHIFT_REG & ~(rnode_20to21_bb6_arrayidx62_0_consumed_1_NO_SHIFT_REG));
assign rnode_20to21_bb6_arrayidx62_0_NO_SHIFT_REG = rnode_20to21_bb6_arrayidx62_0_reg_21_NO_SHIFT_REG;
assign rnode_20to21_bb6_arrayidx62_1_NO_SHIFT_REG = rnode_20to21_bb6_arrayidx62_0_reg_21_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rnode_20to21_bb6_arrayidx62_0_consumed_0_NO_SHIFT_REG <= 1'b0;
		rnode_20to21_bb6_arrayidx62_0_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rnode_20to21_bb6_arrayidx62_0_consumed_0_NO_SHIFT_REG <= (rnode_20to21_bb6_arrayidx62_0_valid_out_0_reg_21_NO_SHIFT_REG & (rnode_20to21_bb6_arrayidx62_0_consumed_0_NO_SHIFT_REG | ~(rnode_20to21_bb6_arrayidx62_0_stall_in_0_NO_SHIFT_REG)) & rnode_20to21_bb6_arrayidx62_0_stall_in_0_reg_21_NO_SHIFT_REG);
		rnode_20to21_bb6_arrayidx62_0_consumed_1_NO_SHIFT_REG <= (rnode_20to21_bb6_arrayidx62_0_valid_out_0_reg_21_NO_SHIFT_REG & (rnode_20to21_bb6_arrayidx62_0_consumed_1_NO_SHIFT_REG | ~(rnode_20to21_bb6_arrayidx62_0_stall_in_1_NO_SHIFT_REG)) & rnode_20to21_bb6_arrayidx62_0_stall_in_0_reg_21_NO_SHIFT_REG);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_valid_out_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_stall_in_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_inputs_ready_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_valid_out_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_3_NO_SHIFT_REG;
 logic rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_stall_out_reg_3_NO_SHIFT_REG;

acl_data_fifo rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_3_NO_SHIFT_REG),
	.valid_out(rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_valid_out_reg_3_NO_SHIFT_REG),
	.stall_out(rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_stall_out_reg_3_NO_SHIFT_REG),
	.data_in(local_bb6_do_directly_for_end57_loopexit_select),
	.data_out(rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_NO_SHIFT_REG)
);

defparam rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_fifo.DEPTH = 1;
defparam rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_fifo.DATA_WIDTH = 1;
defparam rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_fifo.IMPL = "shift_reg";

assign rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb6_do_directly_for_end57_loopexit_select_stall_in_2 = 1'b0;
assign rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG = rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_reg_3_NO_SHIFT_REG;
assign rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_3_NO_SHIFT_REG = 1'b0;
assign rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb6_div58_inputs_ready;
 reg local_bb6_div58_valid_out_NO_SHIFT_REG;
wire local_bb6_div58_stall_in;
wire local_bb6_div58_output_regs_ready;
wire [31:0] local_bb6_div58;
 reg local_bb6_div58_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_1_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_2_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_3_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_4_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_5_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_6_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_7_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_8_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_9_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_10_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_11_NO_SHIFT_REG;
 reg local_bb6_div58_valid_pipe_12_NO_SHIFT_REG;
wire local_bb6_div58_causedstall;

acl_fp_div_s5 fp_module_local_bb6_div58 (
	.clock(clock),
	.dataa(local_bb6_select78),
	.datab(local_bb6_select81),
	.enable(local_bb6_div58_output_regs_ready),
	.result(local_bb6_div58)
);


assign local_bb6_div58_inputs_ready = 1'b1;
assign local_bb6_div58_output_regs_ready = 1'b1;
assign local_bb6_select78_stall_in = 1'b0;
assign local_bb6_select81_stall_in = 1'b0;
assign local_bb6_div58_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_div58_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_2_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_3_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_4_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_5_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_6_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_7_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_8_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_9_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_10_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_11_NO_SHIFT_REG <= 1'b0;
		local_bb6_div58_valid_pipe_12_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_div58_output_regs_ready)
		begin
			local_bb6_div58_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb6_div58_valid_pipe_1_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_0_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_2_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_1_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_3_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_2_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_4_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_3_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_5_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_4_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_6_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_5_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_7_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_6_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_8_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_7_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_9_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_8_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_10_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_9_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_11_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_10_NO_SHIFT_REG;
			local_bb6_div58_valid_pipe_12_NO_SHIFT_REG <= local_bb6_div58_valid_pipe_11_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_div58_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_div58_output_regs_ready)
		begin
			local_bb6_div58_valid_out_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb6_div58_stall_in))
			begin
				local_bb6_div58_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_5_6_0_inputs_ready;
 reg SFC_4_VALID_5_6_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_5_6_0_stall_in;
wire SFC_4_VALID_5_6_0_output_regs_ready;
 reg SFC_4_VALID_5_6_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_5_6_0_causedstall;

assign SFC_4_VALID_5_6_0_inputs_ready = 1'b1;
assign SFC_4_VALID_5_6_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_4_5_0_stall_in = 1'b0;
assign SFC_4_VALID_5_6_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_5_6_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_5_6_0_output_regs_ready)
		begin
			SFC_4_VALID_5_6_0_NO_SHIFT_REG <= SFC_4_VALID_4_5_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_cmp8_not_stall_local;
wire local_bb6_cmp8_not;

assign local_bb6_cmp8_not = (local_bb6_cmp88_acl_ffwd_dest_i1_8 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb6__arrayidx62_valid_out;
wire local_bb6__arrayidx62_stall_in;
wire local_bb6__arrayidx62_inputs_ready;
wire local_bb6__arrayidx62_stall_local;
 reg [63:0] ffwd_12_0_reg_NO_SHIFT_REG;

assign local_bb6__arrayidx62_inputs_ready = rnode_20to21_bb6_arrayidx62_0_valid_out_1_NO_SHIFT_REG;
assign ffwd_12_0 = ffwd_12_0_reg_NO_SHIFT_REG;
assign local_bb6__arrayidx62_valid_out = local_bb6__arrayidx62_inputs_ready;
assign local_bb6__arrayidx62_stall_local = local_bb6__arrayidx62_stall_in;
assign rnode_20to21_bb6_arrayidx62_0_stall_in_1_NO_SHIFT_REG = (|local_bb6__arrayidx62_stall_local);

always @(posedge clock)
begin
	if ((1'b1 & local_bb6__arrayidx62_inputs_ready))
	begin
		ffwd_12_0_reg_NO_SHIFT_REG <= (rnode_20to21_bb6_arrayidx62_1_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC);
	end
end


// Register node:
//  * latency = 12
//  * capacity = 12
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_valid_out_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_stall_in_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_inputs_ready_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_valid_out_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_15_NO_SHIFT_REG;
 logic rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_stall_out_reg_15_NO_SHIFT_REG;

acl_data_fifo rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_15_NO_SHIFT_REG),
	.valid_out(rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_valid_out_reg_15_NO_SHIFT_REG),
	.stall_out(rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_stall_out_reg_15_NO_SHIFT_REG),
	.data_in(rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG),
	.data_out(rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_NO_SHIFT_REG)
);

defparam rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_fifo.DEPTH = 12;
defparam rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_fifo.DATA_WIDTH = 1;
defparam rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_fifo.IMPL = "shift_reg";

assign rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_2to3_bb6_do_directly_for_end57_loopexit_select_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG = rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_reg_15_NO_SHIFT_REG;
assign rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_15_NO_SHIFT_REG = 1'b0;
assign rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_4_VALID_6_7_0_inputs_ready;
 reg SFC_4_VALID_6_7_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_6_7_0_stall_in;
wire SFC_4_VALID_6_7_0_output_regs_ready;
 reg SFC_4_VALID_6_7_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_6_7_0_causedstall;

assign SFC_4_VALID_6_7_0_inputs_ready = 1'b1;
assign SFC_4_VALID_6_7_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_5_6_0_stall_in = 1'b0;
assign SFC_4_VALID_6_7_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_6_7_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_6_7_0_output_regs_ready)
		begin
			SFC_4_VALID_6_7_0_NO_SHIFT_REG <= SFC_4_VALID_5_6_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_not__phi_decision91_select_stall_local;
wire local_bb6_not__phi_decision91_select;

assign local_bb6_not__phi_decision91_select = (local_bb6__acl_ffwd_dest_i1_5_u98 & local_bb6_cmp8_not);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_valid_out_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_stall_in_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_inputs_ready_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_valid_out_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_16_NO_SHIFT_REG;
 logic rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_stall_out_reg_16_NO_SHIFT_REG;

acl_data_fifo rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_16_NO_SHIFT_REG),
	.valid_out(rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_valid_out_reg_16_NO_SHIFT_REG),
	.stall_out(rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_stall_out_reg_16_NO_SHIFT_REG),
	.data_in(rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG),
	.data_out(rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_NO_SHIFT_REG)
);

defparam rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_fifo.DEPTH = 1;
defparam rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_fifo.DATA_WIDTH = 1;
defparam rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_fifo.IMPL = "shift_reg";

assign rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_3to15_bb6_do_directly_for_end57_loopexit_select_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG = rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_reg_16_NO_SHIFT_REG;
assign rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_stall_in_reg_16_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire SFC_4_VALID_7_8_0_inputs_ready;
 reg SFC_4_VALID_7_8_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_7_8_0_stall_in;
wire SFC_4_VALID_7_8_0_output_regs_ready;
 reg SFC_4_VALID_7_8_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_7_8_0_causedstall;

assign SFC_4_VALID_7_8_0_inputs_ready = 1'b1;
assign SFC_4_VALID_7_8_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_6_7_0_stall_in = 1'b0;
assign SFC_4_VALID_7_8_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_7_8_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_7_8_0_output_regs_ready)
		begin
			SFC_4_VALID_7_8_0_NO_SHIFT_REG <= SFC_4_VALID_6_7_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_do_directly_for_end57_select_stall_local;
wire local_bb6_do_directly_for_end57_select;

assign local_bb6_do_directly_for_end57_select = (local_bb6__acl_ffwd_dest_i1_9_u99 & local_bb6_not__phi_decision91_select);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exi134_stall_local;
wire [95:0] local_bb6_c0_exi134;

assign local_bb6_c0_exi134[7:0] = 8'bx;
assign local_bb6_c0_exi134[8] = local_bb6_not__phi_decision91_select;
assign local_bb6_c0_exi134[95:9] = 87'bx;

// This section implements a registered operation.
// 
wire SFC_4_VALID_8_9_0_inputs_ready;
 reg SFC_4_VALID_8_9_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_8_9_0_stall_in;
wire SFC_4_VALID_8_9_0_output_regs_ready;
 reg SFC_4_VALID_8_9_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_8_9_0_causedstall;

assign SFC_4_VALID_8_9_0_inputs_ready = 1'b1;
assign SFC_4_VALID_8_9_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_7_8_0_stall_in = 1'b0;
assign SFC_4_VALID_8_9_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_8_9_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_8_9_0_output_regs_ready)
		begin
			SFC_4_VALID_8_9_0_NO_SHIFT_REG <= SFC_4_VALID_7_8_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_or_stall_local;
wire local_bb6_or;

assign local_bb6_or = (local_bb6_do_directly_for_end57_select | rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exi235_stall_local;
wire [95:0] local_bb6_c0_exi235;

assign local_bb6_c0_exi235[31:0] = local_bb6_c0_exi134[31:0];
assign local_bb6_c0_exi235[63:32] = local_bb6_div58;
assign local_bb6_c0_exi235[95:64] = local_bb6_c0_exi134[95:64];

// This section implements a registered operation.
// 
wire SFC_4_VALID_9_10_0_inputs_ready;
 reg SFC_4_VALID_9_10_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_9_10_0_stall_in;
wire SFC_4_VALID_9_10_0_output_regs_ready;
 reg SFC_4_VALID_9_10_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_9_10_0_causedstall;

assign SFC_4_VALID_9_10_0_inputs_ready = 1'b1;
assign SFC_4_VALID_9_10_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_8_9_0_stall_in = 1'b0;
assign SFC_4_VALID_9_10_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_9_10_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_9_10_0_output_regs_ready)
		begin
			SFC_4_VALID_9_10_0_NO_SHIFT_REG <= SFC_4_VALID_8_9_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_cmp_phi_decision85_xor_or_stall_local;
wire local_bb6_cmp_phi_decision85_xor_or;

assign local_bb6_cmp_phi_decision85_xor_or = (local_bb6_or ^ 1'b1);

// This section implements a registered operation.
// 
wire SFC_4_VALID_10_11_0_inputs_ready;
 reg SFC_4_VALID_10_11_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_10_11_0_stall_in;
wire SFC_4_VALID_10_11_0_output_regs_ready;
 reg SFC_4_VALID_10_11_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_10_11_0_causedstall;

assign SFC_4_VALID_10_11_0_inputs_ready = 1'b1;
assign SFC_4_VALID_10_11_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_9_10_0_stall_in = 1'b0;
assign SFC_4_VALID_10_11_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_10_11_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_10_11_0_output_regs_ready)
		begin
			SFC_4_VALID_10_11_0_NO_SHIFT_REG <= SFC_4_VALID_9_10_0_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_c0_exi336_valid_out;
wire local_bb6_c0_exi336_stall_in;
wire local_bb6_c0_exi336_inputs_ready;
wire local_bb6_c0_exi336_stall_local;
wire [95:0] local_bb6_c0_exi336;

assign local_bb6_c0_exi336_inputs_ready = (local_bb6_div58_valid_out_NO_SHIFT_REG & rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_valid_out_NO_SHIFT_REG & rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_valid_out_NO_SHIFT_REG & rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_valid_out_NO_SHIFT_REG & rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_valid_out_NO_SHIFT_REG);
assign local_bb6_c0_exi336[63:0] = local_bb6_c0_exi235[63:0];
assign local_bb6_c0_exi336[64] = local_bb6_cmp_phi_decision85_xor_or;
assign local_bb6_c0_exi336[95:65] = local_bb6_c0_exi235[95:65];
assign local_bb6_c0_exi336_valid_out = 1'b1;
assign local_bb6_div58_stall_in = 1'b0;
assign rnode_15to16_bb6_cmp88_acl_ffwd_dest_i1_8_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_5_u98_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6__acl_ffwd_dest_i1_9_u99_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_15to16_bb6_do_directly_for_end57_loopexit_select_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire SFC_4_VALID_11_12_0_inputs_ready;
 reg SFC_4_VALID_11_12_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_11_12_0_stall_in;
wire SFC_4_VALID_11_12_0_output_regs_ready;
 reg SFC_4_VALID_11_12_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_11_12_0_causedstall;

assign SFC_4_VALID_11_12_0_inputs_ready = 1'b1;
assign SFC_4_VALID_11_12_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_10_11_0_stall_in = 1'b0;
assign SFC_4_VALID_11_12_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_11_12_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_11_12_0_output_regs_ready)
		begin
			SFC_4_VALID_11_12_0_NO_SHIFT_REG <= SFC_4_VALID_10_11_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_12_13_0_inputs_ready;
 reg SFC_4_VALID_12_13_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_12_13_0_stall_in;
wire SFC_4_VALID_12_13_0_output_regs_ready;
 reg SFC_4_VALID_12_13_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_12_13_0_causedstall;

assign SFC_4_VALID_12_13_0_inputs_ready = 1'b1;
assign SFC_4_VALID_12_13_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_11_12_0_stall_in = 1'b0;
assign SFC_4_VALID_12_13_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_12_13_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_12_13_0_output_regs_ready)
		begin
			SFC_4_VALID_12_13_0_NO_SHIFT_REG <= SFC_4_VALID_11_12_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_13_14_0_inputs_ready;
 reg SFC_4_VALID_13_14_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_13_14_0_stall_in;
wire SFC_4_VALID_13_14_0_output_regs_ready;
 reg SFC_4_VALID_13_14_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_13_14_0_causedstall;

assign SFC_4_VALID_13_14_0_inputs_ready = 1'b1;
assign SFC_4_VALID_13_14_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_12_13_0_stall_in = 1'b0;
assign SFC_4_VALID_13_14_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_13_14_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_13_14_0_output_regs_ready)
		begin
			SFC_4_VALID_13_14_0_NO_SHIFT_REG <= SFC_4_VALID_12_13_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_14_15_0_inputs_ready;
 reg SFC_4_VALID_14_15_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_14_15_0_stall_in;
wire SFC_4_VALID_14_15_0_output_regs_ready;
 reg SFC_4_VALID_14_15_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_14_15_0_causedstall;

assign SFC_4_VALID_14_15_0_inputs_ready = 1'b1;
assign SFC_4_VALID_14_15_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_13_14_0_stall_in = 1'b0;
assign SFC_4_VALID_14_15_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_14_15_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_14_15_0_output_regs_ready)
		begin
			SFC_4_VALID_14_15_0_NO_SHIFT_REG <= SFC_4_VALID_13_14_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire SFC_4_VALID_15_16_0_inputs_ready;
 reg SFC_4_VALID_15_16_0_valid_out_NO_SHIFT_REG;
wire SFC_4_VALID_15_16_0_stall_in;
wire SFC_4_VALID_15_16_0_output_regs_ready;
 reg SFC_4_VALID_15_16_0_NO_SHIFT_REG /* synthesis  preserve  */;
wire SFC_4_VALID_15_16_0_causedstall;

assign SFC_4_VALID_15_16_0_inputs_ready = 1'b1;
assign SFC_4_VALID_15_16_0_output_regs_ready = 1'b1;
assign SFC_4_VALID_14_15_0_stall_in = 1'b0;
assign SFC_4_VALID_15_16_0_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		SFC_4_VALID_15_16_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (SFC_4_VALID_15_16_0_output_regs_ready)
		begin
			SFC_4_VALID_15_16_0_NO_SHIFT_REG <= SFC_4_VALID_14_15_0_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb6_c0_exit37_c0_exi336_inputs_ready;
 reg local_bb6_c0_exit37_c0_exi336_valid_out_0_NO_SHIFT_REG;
wire local_bb6_c0_exit37_c0_exi336_stall_in_0;
 reg local_bb6_c0_exit37_c0_exi336_valid_out_1_NO_SHIFT_REG;
wire local_bb6_c0_exit37_c0_exi336_stall_in_1;
 reg local_bb6_c0_exit37_c0_exi336_valid_out_2_NO_SHIFT_REG;
wire local_bb6_c0_exit37_c0_exi336_stall_in_2;
 reg [95:0] local_bb6_c0_exit37_c0_exi336_NO_SHIFT_REG;
wire [95:0] local_bb6_c0_exit37_c0_exi336_in;
wire local_bb6_c0_exit37_c0_exi336_valid;
wire local_bb6_c0_exit37_c0_exi336_causedstall;

acl_stall_free_sink local_bb6_c0_exit37_c0_exi336_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb6_c0_exi336),
	.data_out(local_bb6_c0_exit37_c0_exi336_in),
	.input_accepted(local_bb6_c0_enter33__input_accepted),
	.valid_out(local_bb6_c0_exit37_c0_exi336_valid),
	.stall_in(~(local_bb6_c0_exit37_c0_exi336_output_regs_ready)),
	.stall_entry(local_bb6_c0_exit37_c0_exi336_entry_stall),
	.valid_in(local_bb6_c0_exit37_c0_exi336_valid_in),
	.IIphases(local_bb6_c0_exit37_c0_exi336_phases),
	.inc_pipelined_thread(local_bb6_c0_enter33__inc_pipelined_thread),
	.dec_pipelined_thread(local_bb6_c0_enter33__dec_pipelined_thread)
);

defparam local_bb6_c0_exit37_c0_exi336_instance.DATA_WIDTH = 96;
defparam local_bb6_c0_exit37_c0_exi336_instance.PIPELINE_DEPTH = 20;
defparam local_bb6_c0_exit37_c0_exi336_instance.SHARINGII = 1;
defparam local_bb6_c0_exit37_c0_exi336_instance.SCHEDULEII = 1;
defparam local_bb6_c0_exit37_c0_exi336_instance.ALWAYS_THROTTLE = 0;

assign local_bb6_c0_exit37_c0_exi336_inputs_ready = 1'b1;
assign local_bb6_c0_exit37_c0_exi336_output_regs_ready = ((~(local_bb6_c0_exit37_c0_exi336_valid_out_0_NO_SHIFT_REG) | ~(local_bb6_c0_exit37_c0_exi336_stall_in_0)) & (~(local_bb6_c0_exit37_c0_exi336_valid_out_1_NO_SHIFT_REG) | ~(local_bb6_c0_exit37_c0_exi336_stall_in_1)) & (~(local_bb6_c0_exit37_c0_exi336_valid_out_2_NO_SHIFT_REG) | ~(local_bb6_c0_exit37_c0_exi336_stall_in_2)));
assign local_bb6_c0_exit37_c0_exi336_valid_in = SFC_4_VALID_15_16_0_NO_SHIFT_REG;
assign local_bb6_c0_exi336_stall_in = 1'b0;
assign SFC_4_VALID_15_16_0_stall_in = 1'b0;
assign local_bb6_c0_exit37_c0_exi336_causedstall = (1'b1 && (1'b0 && !(~(local_bb6_c0_exit37_c0_exi336_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_c0_exit37_c0_exi336_NO_SHIFT_REG <= 'x;
		local_bb6_c0_exit37_c0_exi336_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_exit37_c0_exi336_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb6_c0_exit37_c0_exi336_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_c0_exit37_c0_exi336_output_regs_ready)
		begin
			local_bb6_c0_exit37_c0_exi336_NO_SHIFT_REG <= local_bb6_c0_exit37_c0_exi336_in;
			local_bb6_c0_exit37_c0_exi336_valid_out_0_NO_SHIFT_REG <= local_bb6_c0_exit37_c0_exi336_valid;
			local_bb6_c0_exit37_c0_exi336_valid_out_1_NO_SHIFT_REG <= local_bb6_c0_exit37_c0_exi336_valid;
			local_bb6_c0_exit37_c0_exi336_valid_out_2_NO_SHIFT_REG <= local_bb6_c0_exit37_c0_exi336_valid;
		end
		else
		begin
			if (~(local_bb6_c0_exit37_c0_exi336_stall_in_0))
			begin
				local_bb6_c0_exit37_c0_exi336_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_exit37_c0_exi336_stall_in_1))
			begin
				local_bb6_c0_exit37_c0_exi336_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb6_c0_exit37_c0_exi336_stall_in_2))
			begin
				local_bb6_c0_exit37_c0_exi336_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb6_c0_exe138_valid_out;
wire local_bb6_c0_exe138_stall_in;
wire local_bb6_c0_exe138_inputs_ready;
wire local_bb6_c0_exe138_stall_local;
wire local_bb6_c0_exe138;

assign local_bb6_c0_exe138_inputs_ready = local_bb6_c0_exit37_c0_exi336_valid_out_0_NO_SHIFT_REG;
assign local_bb6_c0_exe138 = local_bb6_c0_exit37_c0_exi336_NO_SHIFT_REG[8];
assign local_bb6_c0_exe138_valid_out = local_bb6_c0_exe138_inputs_ready;
assign local_bb6_c0_exe138_stall_local = local_bb6_c0_exe138_stall_in;
assign local_bb6_c0_exit37_c0_exi336_stall_in_0 = (|local_bb6_c0_exe138_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exe239_valid_out;
wire local_bb6_c0_exe239_stall_in;
wire local_bb6_c0_exe239_inputs_ready;
wire local_bb6_c0_exe239_stall_local;
wire [31:0] local_bb6_c0_exe239;

assign local_bb6_c0_exe239_inputs_ready = local_bb6_c0_exit37_c0_exi336_valid_out_1_NO_SHIFT_REG;
assign local_bb6_c0_exe239 = local_bb6_c0_exit37_c0_exi336_NO_SHIFT_REG[63:32];
assign local_bb6_c0_exe239_valid_out = local_bb6_c0_exe239_inputs_ready;
assign local_bb6_c0_exe239_stall_local = local_bb6_c0_exe239_stall_in;
assign local_bb6_c0_exit37_c0_exi336_stall_in_1 = (|local_bb6_c0_exe239_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb6_c0_exe340_valid_out;
wire local_bb6_c0_exe340_stall_in;
wire local_bb6_c0_exe340_inputs_ready;
wire local_bb6_c0_exe340_stall_local;
wire local_bb6_c0_exe340;
wire rci_rcnode_21to180_rc0_bb6__arrayidx62_0_reg_21;

assign local_bb6_c0_exe340_inputs_ready = local_bb6_c0_exit37_c0_exi336_valid_out_2_NO_SHIFT_REG;
assign local_bb6_c0_exe340 = local_bb6_c0_exit37_c0_exi336_NO_SHIFT_REG[64];
assign local_bb6_c0_exe340_valid_out = local_bb6_c0_exe340_inputs_ready;
assign local_bb6_c0_exe340_stall_local = local_bb6_c0_exe340_stall_in;
assign local_bb6_c0_exit37_c0_exi336_stall_in_2 = (|local_bb6_c0_exe340_stall_local);
assign rci_rcnode_21to180_rc0_bb6__arrayidx62_0_reg_21 = local_bb6_c0_exe138;

// Register node:
//  * latency = 159
//  * capacity = 159
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_valid_out_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_stall_in_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_stall_out_0_reg_180_IP_NO_SHIFT_REG;
 logic rcnode_21to180_rc0_bb6__arrayidx62_0_stall_out_0_reg_180_NO_SHIFT_REG;

acl_data_fifo rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_21to180_rc0_bb6__arrayidx62_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rcnode_21to180_rc0_bb6__arrayidx62_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rcnode_21to180_rc0_bb6__arrayidx62_0_stall_out_0_reg_180_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_21to180_rc0_bb6__arrayidx62_0_reg_21),
	.data_out(rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_NO_SHIFT_REG)
);

defparam rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_fifo.DEPTH = 160;
defparam rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_fifo.ALLOW_FULL_WRITE = 0;
defparam rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_fifo.IMPL = "ram";

assign rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_inputs_ready_NO_SHIFT_REG = (local_bb6__arrayidx62_valid_out & local_bb6_c0_exe138_valid_out);
assign rcnode_21to180_rc0_bb6__arrayidx62_0_stall_out_0_reg_180_NO_SHIFT_REG = (~(rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_inputs_ready_NO_SHIFT_REG) | rcnode_21to180_rc0_bb6__arrayidx62_0_stall_out_0_reg_180_IP_NO_SHIFT_REG);
assign local_bb6__arrayidx62_stall_in = rcnode_21to180_rc0_bb6__arrayidx62_0_stall_out_0_reg_180_NO_SHIFT_REG;
assign local_bb6_c0_exe138_stall_in = rcnode_21to180_rc0_bb6__arrayidx62_0_stall_out_0_reg_180_NO_SHIFT_REG;
assign rcnode_21to180_rc0_bb6__arrayidx62_0_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx62_0_reg_180_NO_SHIFT_REG;
assign rcnode_21to180_rc0_bb6__arrayidx62_0_stall_in_reg_180_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx62_0_stall_in_NO_SHIFT_REG;
assign rcnode_21to180_rc0_bb6__arrayidx62_0_valid_out_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx62_0_valid_out_reg_180_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb6_st_c0_exe239_inputs_ready;
 reg local_bb6_st_c0_exe239_valid_out_NO_SHIFT_REG;
wire local_bb6_st_c0_exe239_stall_in;
wire local_bb6_st_c0_exe239_output_regs_ready;
wire local_bb6_st_c0_exe239_fu_stall_out;
wire local_bb6_st_c0_exe239_fu_valid_out;
wire local_bb6_st_c0_exe239_causedstall;
wire rci_rcnode_180to181_rc0_bb6__arrayidx62_0_reg_180;

lsu_top lsu_local_bb6_st_c0_exe239 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb6_st_c0_exe239_fu_stall_out),
	.i_valid(local_bb6_st_c0_exe239_inputs_ready),
	.i_address((rnode_20to21_bb6_arrayidx62_0_NO_SHIFT_REG & 64'hFFFFFFFFFFFFFFFC)),
	.i_writedata(local_bb6_c0_exe239),
	.i_cmpdata(),
	.i_predicate(local_bb6_c0_exe340),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb6_st_c0_exe239_output_regs_ready)),
	.o_valid(local_bb6_st_c0_exe239_fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb6_st_c0_exe239_active),
	.avm_address(avm_local_bb6_st_c0_exe239_address),
	.avm_read(avm_local_bb6_st_c0_exe239_read),
	.avm_readdata(avm_local_bb6_st_c0_exe239_readdata),
	.avm_write(avm_local_bb6_st_c0_exe239_write),
	.avm_writeack(avm_local_bb6_st_c0_exe239_writeack),
	.avm_burstcount(avm_local_bb6_st_c0_exe239_burstcount),
	.avm_writedata(avm_local_bb6_st_c0_exe239_writedata),
	.avm_byteenable(avm_local_bb6_st_c0_exe239_byteenable),
	.avm_waitrequest(avm_local_bb6_st_c0_exe239_waitrequest),
	.avm_readdatavalid(avm_local_bb6_st_c0_exe239_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb6_st_c0_exe239.AWIDTH = 33;
defparam lsu_local_bb6_st_c0_exe239.WIDTH_BYTES = 4;
defparam lsu_local_bb6_st_c0_exe239.MWIDTH_BYTES = 64;
defparam lsu_local_bb6_st_c0_exe239.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb6_st_c0_exe239.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb6_st_c0_exe239.READ = 0;
defparam lsu_local_bb6_st_c0_exe239.ATOMIC = 0;
defparam lsu_local_bb6_st_c0_exe239.WIDTH = 32;
defparam lsu_local_bb6_st_c0_exe239.MWIDTH = 512;
defparam lsu_local_bb6_st_c0_exe239.ATOMIC_WIDTH = 3;
defparam lsu_local_bb6_st_c0_exe239.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb6_st_c0_exe239.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb6_st_c0_exe239.MEMORY_SIDE_MEM_LATENCY = 10;
defparam lsu_local_bb6_st_c0_exe239.USE_WRITE_ACK = 1;
defparam lsu_local_bb6_st_c0_exe239.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb6_st_c0_exe239.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb6_st_c0_exe239.NUMBER_BANKS = 1;
defparam lsu_local_bb6_st_c0_exe239.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb6_st_c0_exe239.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb6_st_c0_exe239.USEINPUTFIFO = 0;
defparam lsu_local_bb6_st_c0_exe239.USECACHING = 0;
defparam lsu_local_bb6_st_c0_exe239.USEOUTPUTFIFO = 1;
defparam lsu_local_bb6_st_c0_exe239.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb6_st_c0_exe239.HIGH_FMAX = 1;
defparam lsu_local_bb6_st_c0_exe239.ADDRSPACE = 1;
defparam lsu_local_bb6_st_c0_exe239.STYLE = "BURST-COALESCED";
defparam lsu_local_bb6_st_c0_exe239.USE_BYTE_EN = 0;

assign local_bb6_st_c0_exe239_inputs_ready = (local_bb6_c0_exe239_valid_out & local_bb6_c0_exe340_valid_out & rnode_20to21_bb6_arrayidx62_0_valid_out_0_NO_SHIFT_REG);
assign local_bb6_st_c0_exe239_output_regs_ready = (&(~(local_bb6_st_c0_exe239_valid_out_NO_SHIFT_REG) | ~(local_bb6_st_c0_exe239_stall_in)));
assign local_bb6_c0_exe239_stall_in = (local_bb6_st_c0_exe239_fu_stall_out | ~(local_bb6_st_c0_exe239_inputs_ready));
assign local_bb6_c0_exe340_stall_in = (local_bb6_st_c0_exe239_fu_stall_out | ~(local_bb6_st_c0_exe239_inputs_ready));
assign rnode_20to21_bb6_arrayidx62_0_stall_in_0_NO_SHIFT_REG = (local_bb6_st_c0_exe239_fu_stall_out | ~(local_bb6_st_c0_exe239_inputs_ready));
assign local_bb6_st_c0_exe239_causedstall = (local_bb6_st_c0_exe239_inputs_ready && (local_bb6_st_c0_exe239_fu_stall_out && !(~(local_bb6_st_c0_exe239_output_regs_ready))));
assign rci_rcnode_180to181_rc0_bb6__arrayidx62_0_reg_180 = rcnode_21to180_rc0_bb6__arrayidx62_0_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb6_st_c0_exe239_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb6_st_c0_exe239_output_regs_ready)
		begin
			local_bb6_st_c0_exe239_valid_out_NO_SHIFT_REG <= local_bb6_st_c0_exe239_fu_valid_out;
		end
		else
		begin
			if (~(local_bb6_st_c0_exe239_stall_in))
			begin
				local_bb6_st_c0_exe239_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_valid_out_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_stall_in_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_stall_out_reg_181_IP_NO_SHIFT_REG;
 logic rcnode_180to181_rc0_bb6__arrayidx62_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rcnode_180to181_rc0_bb6__arrayidx62_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rcnode_180to181_rc0_bb6__arrayidx62_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rcnode_180to181_rc0_bb6__arrayidx62_0_stall_out_reg_181_IP_NO_SHIFT_REG),
	.data_in(rci_rcnode_180to181_rc0_bb6__arrayidx62_0_reg_180),
	.data_out(rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_NO_SHIFT_REG)
);

defparam rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_fifo.DEPTH = 1;
defparam rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_fifo.IMPL = "ll_reg";

assign rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_inputs_ready_NO_SHIFT_REG = rcnode_21to180_rc0_bb6__arrayidx62_0_valid_out_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx62_0_stall_out_reg_181_NO_SHIFT_REG = (~(rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_inputs_ready_NO_SHIFT_REG) | rcnode_180to181_rc0_bb6__arrayidx62_0_stall_out_reg_181_IP_NO_SHIFT_REG);
assign rcnode_21to180_rc0_bb6__arrayidx62_0_stall_in_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx62_0_stall_out_reg_181_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx62_0_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx62_0_reg_181_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx62_0_stall_in_reg_181_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx62_0_stall_in_NO_SHIFT_REG;
assign rcnode_180to181_rc0_bb6__arrayidx62_0_valid_out_NO_SHIFT_REG = rcnode_180to181_rc0_bb6__arrayidx62_0_valid_out_reg_181_NO_SHIFT_REG;

// This section implements a staging register.
// 
wire rstag_181to181_bb6_st_c0_exe239_valid_out;
wire rstag_181to181_bb6_st_c0_exe239_stall_in;
wire rstag_181to181_bb6_st_c0_exe239_inputs_ready;
wire rstag_181to181_bb6_st_c0_exe239_stall_local;
 reg rstag_181to181_bb6_st_c0_exe239_staging_valid_NO_SHIFT_REG;
wire rstag_181to181_bb6_st_c0_exe239_combined_valid;

assign rstag_181to181_bb6_st_c0_exe239_inputs_ready = local_bb6_st_c0_exe239_valid_out_NO_SHIFT_REG;
assign rstag_181to181_bb6_st_c0_exe239_combined_valid = (rstag_181to181_bb6_st_c0_exe239_staging_valid_NO_SHIFT_REG | rstag_181to181_bb6_st_c0_exe239_inputs_ready);
assign rstag_181to181_bb6_st_c0_exe239_valid_out = rstag_181to181_bb6_st_c0_exe239_combined_valid;
assign rstag_181to181_bb6_st_c0_exe239_stall_local = rstag_181to181_bb6_st_c0_exe239_stall_in;
assign local_bb6_st_c0_exe239_stall_in = (|rstag_181to181_bb6_st_c0_exe239_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_181to181_bb6_st_c0_exe239_staging_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (rstag_181to181_bb6_st_c0_exe239_stall_local)
		begin
			if (~(rstag_181to181_bb6_st_c0_exe239_staging_valid_NO_SHIFT_REG))
			begin
				rstag_181to181_bb6_st_c0_exe239_staging_valid_NO_SHIFT_REG <= rstag_181to181_bb6_st_c0_exe239_inputs_ready;
			end
		end
		else
		begin
			rstag_181to181_bb6_st_c0_exe239_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_bb6_indvars_iv_next40_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb6_indvars_iv_next40_valid_out & rcnode_180to181_rc0_bb6__arrayidx62_0_valid_out_NO_SHIFT_REG & rstag_181to181_bb6_st_c0_exe239_valid_out);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb6_indvars_iv_next40_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rcnode_180to181_rc0_bb6__arrayidx62_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rstag_181to181_bb6_st_c0_exe239_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb6_indvars_iv_next40_0 = lvb_bb6_indvars_iv_next40_0_reg_NO_SHIFT_REG;
assign lvb_bb6_indvars_iv_next40_1 = lvb_bb6_indvars_iv_next40_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_bb6_indvars_iv_next40_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb6_indvars_iv_next40_0_reg_NO_SHIFT_REG <= local_bb6_indvars_iv_next40;
			branch_compare_result_NO_SHIFT_REG <= rcnode_180to181_rc0_bb6__arrayidx62_0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_7
	(
		input 		clock,
		input 		resetn,
		input 		input_wii_cmp1526,
		input [31:0] 		input_wii_sub24,
		input [31:0] 		input_wii_sub27,
		input [31:0] 		input_wii_mul48,
		input [63:0] 		input_wii_var_,
		input [63:0] 		input_wii_var__u100,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out_0,
		input 		stall_in_0,
		output [31:0] 		lvb_bb7_inc67_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [31:0] 		lvb_bb7_inc67_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input 		ffwd_1_0,
		input [31:0] 		ffwd_0_0,
		input 		ffwd_5_0,
		output [31:0] 		ffwd_13_0
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb7_cmp3_acl_ffwd_dest_i1_1_stall_local;
wire local_bb7_cmp3_acl_ffwd_dest_i1_1;

assign local_bb7_cmp3_acl_ffwd_dest_i1_1 = ffwd_1_0;

// This section implements an unregistered operation.
// 
wire local_bb7_pos_y_01_acl_ffwd_dest_i32_0_stall_local;
wire [31:0] local_bb7_pos_y_01_acl_ffwd_dest_i32_0;

assign local_bb7_pos_y_01_acl_ffwd_dest_i32_0 = ffwd_0_0;

// This section implements an unregistered operation.
// 
wire local_bb7__acl_ffwd_dest_i1_5_stall_local;
wire local_bb7__acl_ffwd_dest_i1_5;

assign local_bb7__acl_ffwd_dest_i1_5 = ffwd_5_0;

// This section implements an unregistered operation.
// 
wire local_bb7_var__stall_local;
wire [31:0] local_bb7_var_;

assign local_bb7_var_[31:1] = 31'h0;
assign local_bb7_var_[0] = local_bb7_cmp3_acl_ffwd_dest_i1_1;

// This section implements an unregistered operation.
// 
wire local_bb7_inc67_stall_local;
wire [31:0] local_bb7_inc67;

assign local_bb7_inc67 = (local_bb7_pos_y_01_acl_ffwd_dest_i32_0 + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb7_came_from_for_cond_select_stall_local;
wire [31:0] local_bb7_came_from_for_cond_select;

assign local_bb7_came_from_for_cond_select = ((local_bb7_var_ & 32'h1) ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb7_select49_stall_local;
wire [31:0] local_bb7_select49;

assign local_bb7_select49 = (local_bb7__acl_ffwd_dest_i1_5 ? 32'h2 : (local_bb7_came_from_for_cond_select & 32'h1));

// This section implements an unregistered operation.
// 
wire local_bb7_for_cond_branch_back_stall_local;
wire local_bb7_for_cond_branch_back;

assign local_bb7_for_cond_branch_back = ((local_bb7_select49 & 32'h3) == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb7_for_cond_branch_back_valid_out;
wire local_bb7_for_cond_branch_back_stall_in;
wire local_bb7__select49_valid_out;
wire local_bb7__select49_stall_in;
wire local_bb7_inc67_valid_out;
wire local_bb7_inc67_stall_in;
wire local_bb7__select49_inputs_ready;
wire local_bb7__select49_stall_local;
 reg [31:0] ffwd_13_0_reg_NO_SHIFT_REG;

assign local_bb7__select49_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG);
assign ffwd_13_0 = ffwd_13_0_reg_NO_SHIFT_REG;
assign local_bb7__select49_stall_local = (local_bb7_for_cond_branch_back_stall_in | local_bb7__select49_stall_in | local_bb7_inc67_stall_in);
assign local_bb7_for_cond_branch_back_valid_out = local_bb7__select49_inputs_ready;
assign local_bb7__select49_valid_out = local_bb7__select49_inputs_ready;
assign local_bb7_inc67_valid_out = local_bb7__select49_inputs_ready;
assign merge_node_stall_in_0 = (local_bb7__select49_stall_local | ~(local_bb7__select49_inputs_ready));
assign merge_node_stall_in_2 = (local_bb7__select49_stall_local | ~(local_bb7__select49_inputs_ready));
assign merge_node_stall_in_1 = (local_bb7__select49_stall_local | ~(local_bb7__select49_inputs_ready));

always @(posedge clock)
begin
	if ((1'b1 & local_bb7__select49_inputs_ready))
	begin
		ffwd_13_0_reg_NO_SHIFT_REG <= (local_bb7_select49 & 32'h3);
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [31:0] lvb_bb7_inc67_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb7__select49_valid_out & local_bb7_for_cond_branch_back_valid_out & local_bb7_inc67_valid_out);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb7__select49_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb7_for_cond_branch_back_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb7_inc67_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb7_inc67_0 = lvb_bb7_inc67_0_reg_NO_SHIFT_REG;
assign lvb_bb7_inc67_1 = lvb_bb7_inc67_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_bb7_inc67_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb7_inc67_0_reg_NO_SHIFT_REG <= local_bb7_inc67;
			branch_compare_result_NO_SHIFT_REG <= local_bb7_for_cond_branch_back;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_basic_block_8
	(
		input 		clock,
		input 		resetn,
		input 		valid_in,
		output 		stall_out,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start,
		input [31:0] 		ffwd_13_0,
		input [63:0] 		ffwd_12_0,
		input [511:0] 		avm_local_bb8_st__readdata,
		input 		avm_local_bb8_st__readdatavalid,
		input 		avm_local_bb8_st__waitrequest,
		output [32:0] 		avm_local_bb8_st__address,
		output 		avm_local_bb8_st__read,
		output 		avm_local_bb8_st__write,
		input 		avm_local_bb8_st__writeack,
		output [511:0] 		avm_local_bb8_st__writedata,
		output [63:0] 		avm_local_bb8_st__byteenable,
		output [4:0] 		avm_local_bb8_st__burstcount,
		output 		local_bb8_st__active,
		input 		clock2x
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb8_select4912_acl_ffwd_dest_i32_13_stall_local;
wire [31:0] local_bb8_select4912_acl_ffwd_dest_i32_13;

assign local_bb8_select4912_acl_ffwd_dest_i32_13 = ffwd_13_0;

// This section implements an unregistered operation.
// 
wire local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_valid_out;
wire local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_stall_in;
wire local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_inputs_ready;
wire local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_stall_local;
wire [63:0] local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12;

assign local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12 = ffwd_12_0;
assign local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_valid_out = local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_inputs_ready;
assign local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_stall_local = local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_stall_in;
assign merge_node_stall_in_1 = (|local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb8_for_cond_branch_to_dummy_valid_out;
wire local_bb8_for_cond_branch_to_dummy_stall_in;
wire local_bb8_for_cond_branch_to_dummy_inputs_ready;
wire local_bb8_for_cond_branch_to_dummy_stall_local;
wire local_bb8_for_cond_branch_to_dummy;

assign local_bb8_for_cond_branch_to_dummy_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb8_for_cond_branch_to_dummy = (local_bb8_select4912_acl_ffwd_dest_i32_13 == 32'h1);
assign local_bb8_for_cond_branch_to_dummy_valid_out = local_bb8_for_cond_branch_to_dummy_inputs_ready;
assign local_bb8_for_cond_branch_to_dummy_stall_local = local_bb8_for_cond_branch_to_dummy_stall_in;
assign merge_node_stall_in_0 = (|local_bb8_for_cond_branch_to_dummy_stall_local);

// This section implements a registered operation.
// 
wire local_bb8_st__inputs_ready;
 reg local_bb8_st__valid_out_NO_SHIFT_REG;
wire local_bb8_st__stall_in;
wire local_bb8_st__output_regs_ready;
wire local_bb8_st__fu_stall_out;
wire local_bb8_st__fu_valid_out;
wire local_bb8_st__causedstall;

lsu_top lsu_local_bb8_st_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb8_st__fu_stall_out),
	.i_valid(local_bb8_st__inputs_ready),
	.i_address(local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12),
	.i_writedata(32'h0),
	.i_cmpdata(),
	.i_predicate(local_bb8_for_cond_branch_to_dummy),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb8_st__output_regs_ready)),
	.o_valid(local_bb8_st__fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb8_st__active),
	.avm_address(avm_local_bb8_st__address),
	.avm_read(avm_local_bb8_st__read),
	.avm_readdata(avm_local_bb8_st__readdata),
	.avm_write(avm_local_bb8_st__write),
	.avm_writeack(avm_local_bb8_st__writeack),
	.avm_burstcount(avm_local_bb8_st__burstcount),
	.avm_writedata(avm_local_bb8_st__writedata),
	.avm_byteenable(avm_local_bb8_st__byteenable),
	.avm_waitrequest(avm_local_bb8_st__waitrequest),
	.avm_readdatavalid(avm_local_bb8_st__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb8_st_.AWIDTH = 33;
defparam lsu_local_bb8_st_.WIDTH_BYTES = 4;
defparam lsu_local_bb8_st_.MWIDTH_BYTES = 64;
defparam lsu_local_bb8_st_.WRITEDATAWIDTH_BYTES = 64;
defparam lsu_local_bb8_st_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb8_st_.READ = 0;
defparam lsu_local_bb8_st_.ATOMIC = 0;
defparam lsu_local_bb8_st_.WIDTH = 32;
defparam lsu_local_bb8_st_.MWIDTH = 512;
defparam lsu_local_bb8_st_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb8_st_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb8_st_.KERNEL_SIDE_MEM_LATENCY = 4;
defparam lsu_local_bb8_st_.MEMORY_SIDE_MEM_LATENCY = 10;
defparam lsu_local_bb8_st_.USE_WRITE_ACK = 0;
defparam lsu_local_bb8_st_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb8_st_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb8_st_.NUMBER_BANKS = 1;
defparam lsu_local_bb8_st_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb8_st_.INTENDED_DEVICE_FAMILY = "Stratix V";
defparam lsu_local_bb8_st_.USEINPUTFIFO = 0;
defparam lsu_local_bb8_st_.USECACHING = 0;
defparam lsu_local_bb8_st_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb8_st_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb8_st_.HIGH_FMAX = 1;
defparam lsu_local_bb8_st_.ADDRSPACE = 1;
defparam lsu_local_bb8_st_.STYLE = "BURST-COALESCED";
defparam lsu_local_bb8_st_.USE_BYTE_EN = 0;

assign local_bb8_st__inputs_ready = (local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_valid_out & local_bb8_for_cond_branch_to_dummy_valid_out);
assign local_bb8_st__output_regs_ready = (&(~(local_bb8_st__valid_out_NO_SHIFT_REG) | ~(local_bb8_st__stall_in)));
assign local_bb8_arrayidx6211_acl_ffwd_dest_p1f_12_stall_in = (local_bb8_st__fu_stall_out | ~(local_bb8_st__inputs_ready));
assign local_bb8_for_cond_branch_to_dummy_stall_in = (local_bb8_st__fu_stall_out | ~(local_bb8_st__inputs_ready));
assign local_bb8_st__causedstall = (local_bb8_st__inputs_ready && (local_bb8_st__fu_stall_out && !(~(local_bb8_st__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb8_st__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb8_st__output_regs_ready)
		begin
			local_bb8_st__valid_out_NO_SHIFT_REG <= local_bb8_st__fu_valid_out;
		end
		else
		begin
			if (~(local_bb8_st__stall_in))
			begin
				local_bb8_st__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_5to5_bb8_st__valid_out;
wire rstag_5to5_bb8_st__stall_in;
wire rstag_5to5_bb8_st__inputs_ready;
wire rstag_5to5_bb8_st__stall_local;
 reg rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb8_st__combined_valid;

assign rstag_5to5_bb8_st__inputs_ready = local_bb8_st__valid_out_NO_SHIFT_REG;
assign rstag_5to5_bb8_st__combined_valid = (rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG | rstag_5to5_bb8_st__inputs_ready);
assign rstag_5to5_bb8_st__valid_out = rstag_5to5_bb8_st__combined_valid;
assign rstag_5to5_bb8_st__stall_local = rstag_5to5_bb8_st__stall_in;
assign local_bb8_st__stall_in = (|rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (rstag_5to5_bb8_st__stall_local)
		begin
			if (~(rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG <= rstag_5to5_bb8_st__inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb8_st__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
wire branch_var__output_regs_ready;

assign branch_var__inputs_ready = rstag_5to5_bb8_st__valid_out;
assign branch_var__output_regs_ready = ~(stall_in);
assign rstag_5to5_bb8_st__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out = branch_var__inputs_ready;

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_function
	(
		input 		clock,
		input 		resetn,
		output 		stall_out,
		input 		valid_in,
		output 		valid_out,
		input 		stall_in,
		input [511:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [32:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [511:0] 		avm_local_bb2_ld__writedata,
		output [63:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		input [511:0] 		avm_local_bb4_ld__readdata,
		input 		avm_local_bb4_ld__readdatavalid,
		input 		avm_local_bb4_ld__waitrequest,
		output [32:0] 		avm_local_bb4_ld__address,
		output 		avm_local_bb4_ld__read,
		output 		avm_local_bb4_ld__write,
		input 		avm_local_bb4_ld__writeack,
		output [511:0] 		avm_local_bb4_ld__writedata,
		output [63:0] 		avm_local_bb4_ld__byteenable,
		output [4:0] 		avm_local_bb4_ld__burstcount,
		input [511:0] 		avm_local_bb6_st_c0_exe239_readdata,
		input 		avm_local_bb6_st_c0_exe239_readdatavalid,
		input 		avm_local_bb6_st_c0_exe239_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe239_address,
		output 		avm_local_bb6_st_c0_exe239_read,
		output 		avm_local_bb6_st_c0_exe239_write,
		input 		avm_local_bb6_st_c0_exe239_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe239_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe239_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe239_burstcount,
		input [511:0] 		avm_local_bb8_st__readdata,
		input 		avm_local_bb8_st__readdatavalid,
		input 		avm_local_bb8_st__waitrequest,
		output [32:0] 		avm_local_bb8_st__address,
		output 		avm_local_bb8_st__read,
		output 		avm_local_bb8_st__write,
		input 		avm_local_bb8_st__writeack,
		output [511:0] 		avm_local_bb8_st__writedata,
		output [63:0] 		avm_local_bb8_st__byteenable,
		output [4:0] 		avm_local_bb8_st__burstcount,
		input 		start,
		input [31:0] 		input_r,
		input [31:0] 		input_global_size_0,
		input [31:0] 		input_global_size_1,
		input [31:0] 		input_e_d,
		input 		clock2x,
		input [63:0] 		input_in,
		input [63:0] 		input_out,
		output reg 		has_a_write_pending,
		output reg 		has_a_lsu_active
	);


wire [31:0] workgroup_size;
wire [31:0] cur_cycle;
wire bb_0_stall_out;
wire bb_0_valid_out;
wire bb_0_lvb_bb0_cmp1526;
wire [31:0] bb_0_lvb_bb0_sub24;
wire [31:0] bb_0_lvb_bb0_sub27;
wire [31:0] bb_0_lvb_bb0_mul48;
wire [63:0] bb_0_lvb_bb0_var_;
wire [63:0] bb_0_lvb_bb0_var__u0;
wire bb_1_stall_out_0;
wire bb_1_stall_out_1;
wire bb_1_valid_out;
wire [31:0] ffwd_0_0;
wire ffwd_1_0;
wire [31:0] ffwd_2_0;
wire bb_2_stall_out_0;
wire bb_2_stall_out_1;
wire bb_2_valid_out;
wire [63:0] ffwd_3_0;
wire [31:0] ffwd_4_0;
wire [63:0] ffwd_6_0;
wire ffwd_5_0;
wire bb_2_local_bb2_ld__active;
wire [31:0] ffwd_7_0;
wire ffwd_8_0;
wire ffwd_9_0;
wire bb_3_stall_out_0;
wire bb_3_stall_out_1;
wire bb_3_valid_out;
wire [31:0] bb_3_lvb_bb3_c0_exe1;
wire [31:0] bb_3_lvb_bb3_c0_exe2;
wire bb_3_lvb_bb3_c0_exe3;
wire bb_3_lvb_bb3_c0_exe4;
wire [31:0] bb_3_lvb_bb3_t_228_pop5_;
wire [31:0] bb_3_lvb_bb3_sum_227_pop6_;
wire bb_3_feedback_stall_out_5;
wire bb_3_feedback_stall_out_6;
wire bb_3_feedback_stall_out_4;
wire bb_3_feedback_stall_out_2;
wire bb_3_feedback_stall_out_3;
wire bb_3_acl_pipelined_valid;
wire bb_3_acl_pipelined_exiting_valid;
wire bb_3_acl_pipelined_exiting_stall;
wire bb_3_feedback_valid_out_3;
wire bb_3_feedback_data_out_3;
wire bb_3_feedback_valid_out_4;
wire [63:0] bb_3_feedback_data_out_4;
wire bb_4_stall_out_0;
wire bb_4_stall_out_1;
wire bb_4_valid_out_0;
wire [191:0] bb_4_lvb_bb4_c0_exit28_c0_exi6_0;
wire bb_4_lvb_bb4_c0_exe6_0;
wire [95:0] bb_4_lvb_bb4_c1_exit_c1_exi2_0;
wire bb_4_valid_out_1;
wire [191:0] bb_4_lvb_bb4_c0_exit28_c0_exi6_1;
wire bb_4_lvb_bb4_c0_exe6_1;
wire [95:0] bb_4_lvb_bb4_c1_exit_c1_exi2_1;
wire bb_4_feedback_stall_out_7;
wire bb_4_feedback_stall_out_11;
wire bb_4_feedback_stall_out_0;
wire bb_4_feedback_stall_out_1;
wire bb_4_acl_pipelined_valid;
wire bb_4_acl_pipelined_exiting_valid;
wire bb_4_acl_pipelined_exiting_stall;
wire bb_4_feedback_stall_out_10;
wire bb_4_feedback_stall_out_12;
wire bb_4_feedback_stall_out_13;
wire bb_4_feedback_valid_out_7;
wire [63:0] bb_4_feedback_data_out_7;
wire bb_4_feedback_valid_out_1;
wire bb_4_feedback_data_out_1;
wire bb_4_feedback_valid_out_10;
wire [31:0] bb_4_feedback_data_out_10;
wire bb_4_feedback_valid_out_12;
wire bb_4_feedback_data_out_12;
wire bb_4_feedback_valid_out_13;
wire bb_4_feedback_data_out_13;
wire bb_4_feedback_valid_out_11;
wire [31:0] bb_4_feedback_data_out_11;
wire bb_4_local_bb4_ld__active;
wire bb_4_feedback_stall_out_9;
wire bb_4_feedback_stall_out_8;
wire bb_4_feedback_valid_out_9;
wire [31:0] bb_4_feedback_data_out_9;
wire [31:0] ffwd_10_0;
wire bb_4_feedback_valid_out_8;
wire [31:0] bb_4_feedback_data_out_8;
wire [31:0] ffwd_11_0;
wire bb_5_stall_out;
wire bb_5_valid_out_0;
wire bb_5_valid_out_1;
wire bb_5_feedback_valid_out_5;
wire [31:0] bb_5_feedback_data_out_5;
wire bb_5_feedback_valid_out_6;
wire [31:0] bb_5_feedback_data_out_6;
wire bb_6_stall_out;
wire bb_6_valid_out_0;
wire [63:0] bb_6_lvb_bb6_indvars_iv_next40_0;
wire bb_6_valid_out_1;
wire [63:0] bb_6_lvb_bb6_indvars_iv_next40_1;
wire [63:0] ffwd_12_0;
wire bb_6_local_bb6_st_c0_exe239_active;
wire bb_7_stall_out;
wire bb_7_valid_out_0;
wire [31:0] bb_7_lvb_bb7_inc67_0;
wire bb_7_valid_out_1;
wire [31:0] bb_7_lvb_bb7_inc67_1;
wire [31:0] ffwd_13_0;
wire bb_8_stall_out;
wire bb_8_valid_out;
wire bb_8_local_bb8_st__active;
wire feedback_stall_3;
wire feedback_valid_3;
wire feedback_data_3;
wire feedback_stall_4;
wire feedback_valid_4;
wire [63:0] feedback_data_4;
wire feedback_stall_1;
wire feedback_valid_1;
wire feedback_data_1;
wire feedback_stall_11;
wire feedback_valid_11;
wire [31:0] feedback_data_11;
wire feedback_stall_10;
wire feedback_valid_10;
wire [31:0] feedback_data_10;
wire feedback_stall_7;
wire feedback_valid_7;
wire [63:0] feedback_data_7;
wire feedback_stall_12;
wire feedback_valid_12;
wire feedback_data_12;
wire feedback_stall_13;
wire feedback_valid_13;
wire feedback_data_13;
wire feedback_stall_9;
wire feedback_valid_9;
wire [31:0] feedback_data_9;
wire feedback_stall_8;
wire feedback_valid_8;
wire [31:0] feedback_data_8;
wire feedback_stall_6;
wire feedback_valid_6;
wire [31:0] feedback_data_6;
wire feedback_stall_5;
wire feedback_valid_5;
wire [31:0] feedback_data_5;
wire loop_limiter_1_stall_out;
wire loop_limiter_1_valid_out;
wire loop_limiter_2_stall_out;
wire loop_limiter_2_valid_out;
wire loop_limiter_3_stall_out;
wire loop_limiter_3_valid_out;
wire [1:0] writes_pending;
wire [3:0] lsus_active;

AOCbilateralFilterkernel_basic_block_0 AOCbilateralFilterkernel_basic_block_0 (
	.clock(clock),
	.resetn(resetn),
	.start(start),
	.input_r(input_r),
	.input_global_size_0(input_global_size_0),
	.input_global_size_1(input_global_size_1),
	.input_e_d(input_e_d),
	.valid_in(valid_in),
	.stall_out(bb_0_stall_out),
	.valid_out(bb_0_valid_out),
	.stall_in(bb_1_stall_out_1),
	.lvb_bb0_cmp1526(bb_0_lvb_bb0_cmp1526),
	.lvb_bb0_sub24(bb_0_lvb_bb0_sub24),
	.lvb_bb0_sub27(bb_0_lvb_bb0_sub27),
	.lvb_bb0_mul48(bb_0_lvb_bb0_mul48),
	.lvb_bb0_var_(bb_0_lvb_bb0_var_),
	.lvb_bb0_var__u0(bb_0_lvb_bb0_var__u0),
	.workgroup_size(workgroup_size)
);


AOCbilateralFilterkernel_basic_block_1 AOCbilateralFilterkernel_basic_block_1 (
	.clock(clock),
	.resetn(resetn),
	.input_global_size_1(input_global_size_1),
	.input_global_size_0(input_global_size_0),
	.input_wii_cmp1526(bb_0_lvb_bb0_cmp1526),
	.input_wii_sub24(bb_0_lvb_bb0_sub24),
	.input_wii_sub27(bb_0_lvb_bb0_sub27),
	.input_wii_mul48(bb_0_lvb_bb0_mul48),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u3(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_7_valid_out_0),
	.stall_out_0(bb_1_stall_out_0),
	.input_pos_y_0_0(bb_7_lvb_bb7_inc67_0),
	.valid_in_1(bb_0_valid_out),
	.stall_out_1(bb_1_stall_out_1),
	.input_pos_y_0_1(32'h0),
	.valid_out(bb_1_valid_out),
	.stall_in(loop_limiter_1_stall_out),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_0_0(ffwd_0_0),
	.ffwd_1_0(ffwd_1_0),
	.ffwd_2_0(ffwd_2_0)
);


AOCbilateralFilterkernel_basic_block_2 AOCbilateralFilterkernel_basic_block_2 (
	.clock(clock),
	.resetn(resetn),
	.input_global_size_0(input_global_size_0),
	.input_in(input_in),
	.input_wii_cmp1526(bb_0_lvb_bb0_cmp1526),
	.input_wii_sub24(bb_0_lvb_bb0_sub24),
	.input_wii_sub27(bb_0_lvb_bb0_sub27),
	.input_wii_mul48(bb_0_lvb_bb0_mul48),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u4(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_6_valid_out_0),
	.stall_out_0(bb_2_stall_out_0),
	.input_indvars_iv39_0(bb_6_lvb_bb6_indvars_iv_next40_0),
	.valid_in_1(loop_limiter_1_valid_out),
	.stall_out_1(bb_2_stall_out_1),
	.input_indvars_iv39_1(64'h0),
	.valid_out(bb_2_valid_out),
	.stall_in(loop_limiter_2_stall_out),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_2_0(ffwd_2_0),
	.ffwd_3_0(ffwd_3_0),
	.ffwd_1_0(ffwd_1_0),
	.ffwd_4_0(ffwd_4_0),
	.ffwd_6_0(ffwd_6_0),
	.ffwd_5_0(ffwd_5_0),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__burstcount),
	.local_bb2_ld__active(bb_2_local_bb2_ld__active),
	.clock2x(clock2x),
	.ffwd_7_0(ffwd_7_0),
	.ffwd_8_0(ffwd_8_0),
	.ffwd_9_0(ffwd_9_0)
);


AOCbilateralFilterkernel_basic_block_3 AOCbilateralFilterkernel_basic_block_3 (
	.clock(clock),
	.resetn(resetn),
	.input_r(input_r),
	.input_wii_cmp1526(bb_0_lvb_bb0_cmp1526),
	.input_wii_sub24(bb_0_lvb_bb0_sub24),
	.input_wii_sub27(bb_0_lvb_bb0_sub27),
	.input_wii_mul48(bb_0_lvb_bb0_mul48),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u11(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_3_acl_pipelined_valid),
	.stall_out_0(bb_3_stall_out_0),
	.input_forked_0(1'b0),
	.valid_in_1(loop_limiter_2_valid_out),
	.stall_out_1(bb_3_stall_out_1),
	.input_forked_1(1'b1),
	.valid_out(bb_3_valid_out),
	.stall_in(loop_limiter_3_stall_out),
	.lvb_bb3_c0_exe1(bb_3_lvb_bb3_c0_exe1),
	.lvb_bb3_c0_exe2(bb_3_lvb_bb3_c0_exe2),
	.lvb_bb3_c0_exe3(bb_3_lvb_bb3_c0_exe3),
	.lvb_bb3_c0_exe4(bb_3_lvb_bb3_c0_exe4),
	.lvb_bb3_t_228_pop5_(bb_3_lvb_bb3_t_228_pop5_),
	.lvb_bb3_sum_227_pop6_(bb_3_lvb_bb3_sum_227_pop6_),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_in_5(feedback_valid_5),
	.feedback_stall_out_5(feedback_stall_5),
	.feedback_data_in_5(feedback_data_5),
	.feedback_valid_in_6(feedback_valid_6),
	.feedback_stall_out_6(feedback_stall_6),
	.feedback_data_in_6(feedback_data_6),
	.feedback_valid_in_4(feedback_valid_4),
	.feedback_stall_out_4(feedback_stall_4),
	.feedback_data_in_4(feedback_data_4),
	.ffwd_9_0(ffwd_9_0),
	.feedback_stall_out_2(bb_3_feedback_stall_out_2),
	.feedback_valid_in_3(feedback_valid_3),
	.feedback_stall_out_3(feedback_stall_3),
	.feedback_data_in_3(feedback_data_3),
	.acl_pipelined_valid(bb_3_acl_pipelined_valid),
	.acl_pipelined_stall(bb_3_stall_out_0),
	.acl_pipelined_exiting_valid(bb_3_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_3_acl_pipelined_exiting_stall),
	.ffwd_4_0(ffwd_4_0),
	.feedback_valid_out_3(feedback_valid_3),
	.feedback_stall_in_3(feedback_stall_3),
	.feedback_data_out_3(feedback_data_3),
	.feedback_valid_out_4(feedback_valid_4),
	.feedback_stall_in_4(feedback_stall_4),
	.feedback_data_out_4(feedback_data_4)
);


AOCbilateralFilterkernel_basic_block_4 AOCbilateralFilterkernel_basic_block_4 (
	.clock(clock),
	.resetn(resetn),
	.input_global_size_0(input_global_size_0),
	.input_in(input_in),
	.input_r(input_r),
	.input_wii_cmp1526(bb_0_lvb_bb0_cmp1526),
	.input_wii_sub24(bb_0_lvb_bb0_sub24),
	.input_wii_sub27(bb_0_lvb_bb0_sub27),
	.input_wii_mul48(bb_0_lvb_bb0_mul48),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u15(bb_0_lvb_bb0_var__u0),
	.valid_in_0(bb_4_acl_pipelined_valid),
	.stall_out_0(bb_4_stall_out_0),
	.input_t_322_0('x),
	.input_sum_321_0('x),
	.input_forked17_0(1'b0),
	.input_sub24_add2318_0('x),
	.input_gaussian_ROM4119_0('x),
	.input_var__u16_0('x),
	.input_notexitcond1520_0('x),
	.valid_in_1(loop_limiter_3_valid_out),
	.stall_out_1(bb_4_stall_out_1),
	.input_t_322_1(bb_3_lvb_bb3_t_228_pop5_),
	.input_sum_321_1(bb_3_lvb_bb3_sum_227_pop6_),
	.input_forked17_1(1'b1),
	.input_sub24_add2318_1(bb_3_lvb_bb3_c0_exe1),
	.input_gaussian_ROM4119_1(bb_3_lvb_bb3_c0_exe2),
	.input_var__u16_1(bb_3_lvb_bb3_c0_exe3),
	.input_notexitcond1520_1(bb_3_lvb_bb3_c0_exe4),
	.valid_out_0(bb_4_valid_out_0),
	.stall_in_0(bb_5_stall_out),
	.lvb_bb4_c0_exit28_c0_exi6_0(bb_4_lvb_bb4_c0_exit28_c0_exi6_0),
	.lvb_bb4_c0_exe6_0(bb_4_lvb_bb4_c0_exe6_0),
	.lvb_bb4_c1_exit_c1_exi2_0(bb_4_lvb_bb4_c1_exit_c1_exi2_0),
	.valid_out_1(bb_4_valid_out_1),
	.stall_in_1(1'b0),
	.lvb_bb4_c0_exit28_c0_exi6_1(bb_4_lvb_bb4_c0_exit28_c0_exi6_1),
	.lvb_bb4_c0_exe6_1(bb_4_lvb_bb4_c0_exe6_1),
	.lvb_bb4_c1_exit_c1_exi2_1(bb_4_lvb_bb4_c1_exit_c1_exi2_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_9_0(ffwd_9_0),
	.ffwd_0_0(ffwd_0_0),
	.feedback_valid_in_7(feedback_valid_7),
	.feedback_stall_out_7(feedback_stall_7),
	.feedback_data_in_7(feedback_data_7),
	.feedback_valid_in_11(feedback_valid_11),
	.feedback_stall_out_11(feedback_stall_11),
	.feedback_data_in_11(feedback_data_11),
	.feedback_stall_out_0(bb_4_feedback_stall_out_0),
	.feedback_valid_in_1(feedback_valid_1),
	.feedback_stall_out_1(feedback_stall_1),
	.feedback_data_in_1(feedback_data_1),
	.acl_pipelined_valid(bb_4_acl_pipelined_valid),
	.acl_pipelined_stall(bb_4_stall_out_0),
	.acl_pipelined_exiting_valid(bb_4_acl_pipelined_exiting_valid),
	.acl_pipelined_exiting_stall(bb_4_acl_pipelined_exiting_stall),
	.feedback_valid_in_10(feedback_valid_10),
	.feedback_stall_out_10(feedback_stall_10),
	.feedback_data_in_10(feedback_data_10),
	.feedback_valid_in_12(feedback_valid_12),
	.feedback_stall_out_12(feedback_stall_12),
	.feedback_data_in_12(feedback_data_12),
	.feedback_valid_in_13(feedback_valid_13),
	.feedback_stall_out_13(feedback_stall_13),
	.feedback_data_in_13(feedback_data_13),
	.feedback_valid_out_7(feedback_valid_7),
	.feedback_stall_in_7(feedback_stall_7),
	.feedback_data_out_7(feedback_data_7),
	.feedback_valid_out_1(feedback_valid_1),
	.feedback_stall_in_1(feedback_stall_1),
	.feedback_data_out_1(feedback_data_1),
	.feedback_valid_out_10(feedback_valid_10),
	.feedback_stall_in_10(feedback_stall_10),
	.feedback_data_out_10(feedback_data_10),
	.feedback_valid_out_12(feedback_valid_12),
	.feedback_stall_in_12(feedback_stall_12),
	.feedback_data_out_12(feedback_data_12),
	.feedback_valid_out_13(feedback_valid_13),
	.feedback_stall_in_13(feedback_stall_13),
	.feedback_data_out_13(feedback_data_13),
	.feedback_valid_out_11(feedback_valid_11),
	.feedback_stall_in_11(feedback_stall_11),
	.feedback_data_out_11(feedback_data_11),
	.avm_local_bb4_ld__readdata(avm_local_bb4_ld__readdata),
	.avm_local_bb4_ld__readdatavalid(avm_local_bb4_ld__readdatavalid),
	.avm_local_bb4_ld__waitrequest(avm_local_bb4_ld__waitrequest),
	.avm_local_bb4_ld__address(avm_local_bb4_ld__address),
	.avm_local_bb4_ld__read(avm_local_bb4_ld__read),
	.avm_local_bb4_ld__write(avm_local_bb4_ld__write),
	.avm_local_bb4_ld__writeack(avm_local_bb4_ld__writeack),
	.avm_local_bb4_ld__writedata(avm_local_bb4_ld__writedata),
	.avm_local_bb4_ld__byteenable(avm_local_bb4_ld__byteenable),
	.avm_local_bb4_ld__burstcount(avm_local_bb4_ld__burstcount),
	.local_bb4_ld__active(bb_4_local_bb4_ld__active),
	.clock2x(clock2x),
	.ffwd_7_0(ffwd_7_0),
	.feedback_valid_in_9(feedback_valid_9),
	.feedback_stall_out_9(feedback_stall_9),
	.feedback_data_in_9(feedback_data_9),
	.feedback_valid_in_8(feedback_valid_8),
	.feedback_stall_out_8(feedback_stall_8),
	.feedback_data_in_8(feedback_data_8),
	.feedback_valid_out_9(feedback_valid_9),
	.feedback_stall_in_9(feedback_stall_9),
	.feedback_data_out_9(feedback_data_9),
	.ffwd_10_0(ffwd_10_0),
	.feedback_valid_out_8(feedback_valid_8),
	.feedback_stall_in_8(feedback_stall_8),
	.feedback_data_out_8(feedback_data_8),
	.ffwd_11_0(ffwd_11_0)
);


AOCbilateralFilterkernel_basic_block_5 AOCbilateralFilterkernel_basic_block_5 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_cmp1526(bb_0_lvb_bb0_cmp1526),
	.input_wii_sub24(bb_0_lvb_bb0_sub24),
	.input_wii_sub27(bb_0_lvb_bb0_sub27),
	.input_wii_mul48(bb_0_lvb_bb0_mul48),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u96(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_4_valid_out_0),
	.stall_out(bb_5_stall_out),
	.input_c0_exit28_c0_exi6(bb_4_lvb_bb4_c0_exit28_c0_exi6_0),
	.input_c0_exe6(bb_4_lvb_bb4_c0_exe6_0),
	.input_c1_exit_c1_exi2(bb_4_lvb_bb4_c1_exit_c1_exi2_0),
	.valid_out_0(bb_5_valid_out_0),
	.stall_in_0(bb_6_stall_out),
	.valid_out_1(bb_5_valid_out_1),
	.stall_in_1(1'b0),
	.workgroup_size(workgroup_size),
	.start(start),
	.feedback_valid_out_5(feedback_valid_5),
	.feedback_stall_in_5(feedback_stall_5),
	.feedback_data_out_5(feedback_data_5),
	.feedback_valid_out_6(feedback_valid_6),
	.feedback_stall_in_6(feedback_stall_6),
	.feedback_data_out_6(feedback_data_6)
);


AOCbilateralFilterkernel_basic_block_6 AOCbilateralFilterkernel_basic_block_6 (
	.clock(clock),
	.resetn(resetn),
	.input_out(input_out),
	.input_wii_cmp1526(bb_0_lvb_bb0_cmp1526),
	.input_wii_sub24(bb_0_lvb_bb0_sub24),
	.input_wii_sub27(bb_0_lvb_bb0_sub27),
	.input_wii_mul48(bb_0_lvb_bb0_mul48),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u97(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_5_valid_out_0),
	.stall_out(bb_6_stall_out),
	.valid_out_0(bb_6_valid_out_0),
	.stall_in_0(bb_2_stall_out_0),
	.lvb_bb6_indvars_iv_next40_0(bb_6_lvb_bb6_indvars_iv_next40_0),
	.valid_out_1(bb_6_valid_out_1),
	.stall_in_1(bb_7_stall_out),
	.lvb_bb6_indvars_iv_next40_1(bb_6_lvb_bb6_indvars_iv_next40_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_9_0(ffwd_9_0),
	.ffwd_5_0(ffwd_5_0),
	.ffwd_11_0(ffwd_11_0),
	.ffwd_10_0(ffwd_10_0),
	.ffwd_6_0(ffwd_6_0),
	.ffwd_3_0(ffwd_3_0),
	.ffwd_8_0(ffwd_8_0),
	.ffwd_12_0(ffwd_12_0),
	.avm_local_bb6_st_c0_exe239_readdata(avm_local_bb6_st_c0_exe239_readdata),
	.avm_local_bb6_st_c0_exe239_readdatavalid(avm_local_bb6_st_c0_exe239_readdatavalid),
	.avm_local_bb6_st_c0_exe239_waitrequest(avm_local_bb6_st_c0_exe239_waitrequest),
	.avm_local_bb6_st_c0_exe239_address(avm_local_bb6_st_c0_exe239_address),
	.avm_local_bb6_st_c0_exe239_read(avm_local_bb6_st_c0_exe239_read),
	.avm_local_bb6_st_c0_exe239_write(avm_local_bb6_st_c0_exe239_write),
	.avm_local_bb6_st_c0_exe239_writeack(avm_local_bb6_st_c0_exe239_writeack),
	.avm_local_bb6_st_c0_exe239_writedata(avm_local_bb6_st_c0_exe239_writedata),
	.avm_local_bb6_st_c0_exe239_byteenable(avm_local_bb6_st_c0_exe239_byteenable),
	.avm_local_bb6_st_c0_exe239_burstcount(avm_local_bb6_st_c0_exe239_burstcount),
	.local_bb6_st_c0_exe239_active(bb_6_local_bb6_st_c0_exe239_active),
	.clock2x(clock2x)
);


AOCbilateralFilterkernel_basic_block_7 AOCbilateralFilterkernel_basic_block_7 (
	.clock(clock),
	.resetn(resetn),
	.input_wii_cmp1526(bb_0_lvb_bb0_cmp1526),
	.input_wii_sub24(bb_0_lvb_bb0_sub24),
	.input_wii_sub27(bb_0_lvb_bb0_sub27),
	.input_wii_mul48(bb_0_lvb_bb0_mul48),
	.input_wii_var_(bb_0_lvb_bb0_var_),
	.input_wii_var__u100(bb_0_lvb_bb0_var__u0),
	.valid_in(bb_6_valid_out_1),
	.stall_out(bb_7_stall_out),
	.valid_out_0(bb_7_valid_out_0),
	.stall_in_0(bb_1_stall_out_0),
	.lvb_bb7_inc67_0(bb_7_lvb_bb7_inc67_0),
	.valid_out_1(bb_7_valid_out_1),
	.stall_in_1(bb_8_stall_out),
	.lvb_bb7_inc67_1(bb_7_lvb_bb7_inc67_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_1_0(ffwd_1_0),
	.ffwd_0_0(ffwd_0_0),
	.ffwd_5_0(ffwd_5_0),
	.ffwd_13_0(ffwd_13_0)
);


AOCbilateralFilterkernel_basic_block_8 AOCbilateralFilterkernel_basic_block_8 (
	.clock(clock),
	.resetn(resetn),
	.valid_in(bb_7_valid_out_1),
	.stall_out(bb_8_stall_out),
	.valid_out(bb_8_valid_out),
	.stall_in(stall_in),
	.workgroup_size(workgroup_size),
	.start(start),
	.ffwd_13_0(ffwd_13_0),
	.ffwd_12_0(ffwd_12_0),
	.avm_local_bb8_st__readdata(avm_local_bb8_st__readdata),
	.avm_local_bb8_st__readdatavalid(avm_local_bb8_st__readdatavalid),
	.avm_local_bb8_st__waitrequest(avm_local_bb8_st__waitrequest),
	.avm_local_bb8_st__address(avm_local_bb8_st__address),
	.avm_local_bb8_st__read(avm_local_bb8_st__read),
	.avm_local_bb8_st__write(avm_local_bb8_st__write),
	.avm_local_bb8_st__writeack(avm_local_bb8_st__writeack),
	.avm_local_bb8_st__writedata(avm_local_bb8_st__writedata),
	.avm_local_bb8_st__byteenable(avm_local_bb8_st__byteenable),
	.avm_local_bb8_st__burstcount(avm_local_bb8_st__burstcount),
	.local_bb8_st__active(bb_8_local_bb8_st__active),
	.clock2x(clock2x)
);


acl_loop_limiter loop_limiter_1 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_1_valid_out),
	.i_stall(bb_2_stall_out_1),
	.i_valid_exit(bb_6_valid_out_1),
	.i_stall_exit(bb_7_stall_out),
	.o_valid(loop_limiter_1_valid_out),
	.o_stall(loop_limiter_1_stall_out)
);

defparam loop_limiter_1.ENTRY_WIDTH = 1;
defparam loop_limiter_1.EXIT_WIDTH = 1;
defparam loop_limiter_1.THRESHOLD = 614;

acl_loop_limiter loop_limiter_2 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_2_valid_out),
	.i_stall(bb_3_stall_out_1),
	.i_valid_exit(bb_3_acl_pipelined_exiting_valid),
	.i_stall_exit(bb_3_acl_pipelined_exiting_stall),
	.o_valid(loop_limiter_2_valid_out),
	.o_stall(loop_limiter_2_stall_out)
);

defparam loop_limiter_2.ENTRY_WIDTH = 1;
defparam loop_limiter_2.EXIT_WIDTH = 1;
defparam loop_limiter_2.THRESHOLD = 2;

acl_loop_limiter loop_limiter_3 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_3_valid_out),
	.i_stall(bb_4_stall_out_1),
	.i_valid_exit(bb_4_acl_pipelined_exiting_valid),
	.i_stall_exit(bb_4_acl_pipelined_exiting_stall),
	.o_valid(loop_limiter_3_valid_out),
	.o_stall(loop_limiter_3_stall_out)
);

defparam loop_limiter_3.ENTRY_WIDTH = 1;
defparam loop_limiter_3.EXIT_WIDTH = 1;
defparam loop_limiter_3.THRESHOLD = 9;

AOCbilateralFilterkernel_sys_cycle_time system_cycle_time_module (
	.clock(clock),
	.resetn(resetn),
	.cur_cycle(cur_cycle)
);


assign workgroup_size = 32'h1;
assign valid_out = bb_8_valid_out;
assign stall_out = bb_0_stall_out;
assign writes_pending[0] = bb_6_local_bb6_st_c0_exe239_active;
assign writes_pending[1] = bb_8_local_bb8_st__active;
assign lsus_active[0] = bb_2_local_bb2_ld__active;
assign lsus_active[1] = bb_4_local_bb4_ld__active;
assign lsus_active[2] = bb_6_local_bb6_st_c0_exe239_active;
assign lsus_active[3] = bb_8_local_bb8_st__active;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		has_a_write_pending <= 1'b0;
		has_a_lsu_active <= 1'b0;
	end
	else
	begin
		has_a_write_pending <= (|writes_pending);
		has_a_lsu_active <= (|lsus_active);
	end
end

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_function_wrapper
	(
		input 		clock,
		input 		resetn,
		input 		clock2x,
		input 		local_router_hang,
		input 		avs_cra_read,
		input 		avs_cra_write,
		input [3:0] 		avs_cra_address,
		input [63:0] 		avs_cra_writedata,
		input [7:0] 		avs_cra_byteenable,
		output reg [63:0] 		avs_cra_readdata,
		output reg 		avs_cra_readdatavalid,
		output 		cra_irq,
		input [511:0] 		avm_local_bb2_ld__inst0_readdata,
		input 		avm_local_bb2_ld__inst0_readdatavalid,
		input 		avm_local_bb2_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb2_ld__inst0_address,
		output 		avm_local_bb2_ld__inst0_read,
		output 		avm_local_bb2_ld__inst0_write,
		input 		avm_local_bb2_ld__inst0_writeack,
		output [511:0] 		avm_local_bb2_ld__inst0_writedata,
		output [63:0] 		avm_local_bb2_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb4_ld__inst0_readdata,
		input 		avm_local_bb4_ld__inst0_readdatavalid,
		input 		avm_local_bb4_ld__inst0_waitrequest,
		output [32:0] 		avm_local_bb4_ld__inst0_address,
		output 		avm_local_bb4_ld__inst0_read,
		output 		avm_local_bb4_ld__inst0_write,
		input 		avm_local_bb4_ld__inst0_writeack,
		output [511:0] 		avm_local_bb4_ld__inst0_writedata,
		output [63:0] 		avm_local_bb4_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb4_ld__inst0_burstcount,
		input [511:0] 		avm_local_bb6_st_c0_exe239_inst0_readdata,
		input 		avm_local_bb6_st_c0_exe239_inst0_readdatavalid,
		input 		avm_local_bb6_st_c0_exe239_inst0_waitrequest,
		output [32:0] 		avm_local_bb6_st_c0_exe239_inst0_address,
		output 		avm_local_bb6_st_c0_exe239_inst0_read,
		output 		avm_local_bb6_st_c0_exe239_inst0_write,
		input 		avm_local_bb6_st_c0_exe239_inst0_writeack,
		output [511:0] 		avm_local_bb6_st_c0_exe239_inst0_writedata,
		output [63:0] 		avm_local_bb6_st_c0_exe239_inst0_byteenable,
		output [4:0] 		avm_local_bb6_st_c0_exe239_inst0_burstcount,
		input [511:0] 		avm_local_bb8_st__inst0_readdata,
		input 		avm_local_bb8_st__inst0_readdatavalid,
		input 		avm_local_bb8_st__inst0_waitrequest,
		output [32:0] 		avm_local_bb8_st__inst0_address,
		output 		avm_local_bb8_st__inst0_read,
		output 		avm_local_bb8_st__inst0_write,
		input 		avm_local_bb8_st__inst0_writeack,
		output [511:0] 		avm_local_bb8_st__inst0_writedata,
		output [63:0] 		avm_local_bb8_st__inst0_byteenable,
		output [4:0] 		avm_local_bb8_st__inst0_burstcount
	);

// Responsible for interfacing a kernel with the outside world. It comprises a
// slave interface to specify the kernel arguments and retain kernel status. 

// This section of the wrapper implements the slave interface.
// twoXclock_consumer uses clock2x, even if nobody inside the kernel does. Keeps interface to acl_iface consistent for all kernels.
 reg start_NO_SHIFT_REG;
 reg started_NO_SHIFT_REG;
wire finish;
 reg [31:0] status_NO_SHIFT_REG;
wire has_a_write_pending;
wire has_a_lsu_active;
 reg [191:0] kernel_arguments_NO_SHIFT_REG;
 reg twoXclock_consumer_NO_SHIFT_REG /* synthesis  preserve  noprune  */;
 reg [31:0] workgroup_size_NO_SHIFT_REG;
 reg [31:0] global_size_NO_SHIFT_REG[2:0];
 reg [31:0] num_groups_NO_SHIFT_REG[2:0];
 reg [31:0] local_size_NO_SHIFT_REG[2:0];
 reg [31:0] work_dim_NO_SHIFT_REG;
 reg [31:0] global_offset_NO_SHIFT_REG[2:0];
 reg [63:0] profile_data_NO_SHIFT_REG;
 reg [31:0] profile_ctrl_NO_SHIFT_REG;
 reg [63:0] profile_start_cycle_NO_SHIFT_REG;
 reg [63:0] profile_stop_cycle_NO_SHIFT_REG;
wire dispatched_all_groups;
wire [31:0] group_id_tmp[2:0];
wire [31:0] global_id_base_out[2:0];
wire start_out;
wire [31:0] local_id[0:0][2:0];
wire [31:0] global_id[0:0][2:0];
wire [31:0] group_id[0:0][2:0];
wire iter_valid_in;
wire iter_stall_out;
wire stall_in;
wire stall_out;
wire valid_in;
wire valid_out;

always @(posedge clock2x or negedge resetn)
begin
	if (~(resetn))
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b1;
	end
end



// Work group dispatcher is responsible for issuing work-groups to id iterator(s)
acl_work_group_dispatcher group_dispatcher (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.num_groups(num_groups_NO_SHIFT_REG),
	.local_size(local_size_NO_SHIFT_REG),
	.stall_in(iter_stall_out),
	.valid_out(iter_valid_in),
	.group_id_out(group_id_tmp),
	.global_id_base_out(global_id_base_out),
	.start_out(start_out),
	.dispatched_all_groups(dispatched_all_groups)
);

defparam group_dispatcher.NUM_COPIES = 1;
defparam group_dispatcher.RUN_FOREVER = 0;


// This section of the wrapper implements an Avalon Slave Interface used to configure a kernel invocation.
// The few words words contain the status and the workgroup size registers.
// The remaining addressable space is reserved for kernel arguments.
 reg [63:0] cra_readdata_st1_NO_SHIFT_REG;
 reg [3:0] cra_addr_st1_NO_SHIFT_REG;
 reg cra_read_st1_NO_SHIFT_REG;
wire [63:0] bitenable;

assign bitenable[7:0] = (avs_cra_byteenable[0] ? 8'hFF : 8'h0);
assign bitenable[15:8] = (avs_cra_byteenable[1] ? 8'hFF : 8'h0);
assign bitenable[23:16] = (avs_cra_byteenable[2] ? 8'hFF : 8'h0);
assign bitenable[31:24] = (avs_cra_byteenable[3] ? 8'hFF : 8'h0);
assign bitenable[39:32] = (avs_cra_byteenable[4] ? 8'hFF : 8'h0);
assign bitenable[47:40] = (avs_cra_byteenable[5] ? 8'hFF : 8'h0);
assign bitenable[55:48] = (avs_cra_byteenable[6] ? 8'hFF : 8'h0);
assign bitenable[63:56] = (avs_cra_byteenable[7] ? 8'hFF : 8'h0);
assign cra_irq = (status_NO_SHIFT_REG[1] | status_NO_SHIFT_REG[3]);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		start_NO_SHIFT_REG <= 1'b0;
		started_NO_SHIFT_REG <= 1'b0;
		kernel_arguments_NO_SHIFT_REG <= 192'h0;
		status_NO_SHIFT_REG <= 32'h30000;
		profile_ctrl_NO_SHIFT_REG <= 32'h4;
		profile_start_cycle_NO_SHIFT_REG <= 64'h0;
		profile_stop_cycle_NO_SHIFT_REG <= 64'hFFFFFFFFFFFFFFFF;
		work_dim_NO_SHIFT_REG <= 32'h0;
		workgroup_size_NO_SHIFT_REG <= 32'h0;
		global_size_NO_SHIFT_REG[0] <= 32'h0;
		global_size_NO_SHIFT_REG[1] <= 32'h0;
		global_size_NO_SHIFT_REG[2] <= 32'h0;
		num_groups_NO_SHIFT_REG[0] <= 32'h0;
		num_groups_NO_SHIFT_REG[1] <= 32'h0;
		num_groups_NO_SHIFT_REG[2] <= 32'h0;
		local_size_NO_SHIFT_REG[0] <= 32'h0;
		local_size_NO_SHIFT_REG[1] <= 32'h0;
		local_size_NO_SHIFT_REG[2] <= 32'h0;
		global_offset_NO_SHIFT_REG[0] <= 32'h0;
		global_offset_NO_SHIFT_REG[1] <= 32'h0;
		global_offset_NO_SHIFT_REG[2] <= 32'h0;
	end
	else
	begin
		if (avs_cra_write)
		begin
			case (avs_cra_address)
				4'h0:
				begin
					status_NO_SHIFT_REG[31:16] <= 16'h3;
					status_NO_SHIFT_REG[15:0] <= ((status_NO_SHIFT_REG[15:0] & ~(bitenable[15:0])) | (avs_cra_writedata[15:0] & bitenable[15:0]));
				end

				4'h1:
				begin
					profile_ctrl_NO_SHIFT_REG <= ((profile_ctrl_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'h3:
				begin
					profile_start_cycle_NO_SHIFT_REG[31:0] <= ((profile_start_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_start_cycle_NO_SHIFT_REG[63:32] <= ((profile_start_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'h4:
				begin
					profile_stop_cycle_NO_SHIFT_REG[31:0] <= ((profile_stop_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_stop_cycle_NO_SHIFT_REG[63:32] <= ((profile_stop_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'h5:
				begin
					work_dim_NO_SHIFT_REG <= ((work_dim_NO_SHIFT_REG & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					workgroup_size_NO_SHIFT_REG <= ((workgroup_size_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'h6:
				begin
					global_size_NO_SHIFT_REG[0] <= ((global_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_size_NO_SHIFT_REG[1] <= ((global_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'h7:
				begin
					global_size_NO_SHIFT_REG[2] <= ((global_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[0] <= ((num_groups_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'h8:
				begin
					num_groups_NO_SHIFT_REG[1] <= ((num_groups_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[2] <= ((num_groups_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'h9:
				begin
					local_size_NO_SHIFT_REG[0] <= ((local_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					local_size_NO_SHIFT_REG[1] <= ((local_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'hA:
				begin
					local_size_NO_SHIFT_REG[2] <= ((local_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[0] <= ((global_offset_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'hB:
				begin
					global_offset_NO_SHIFT_REG[1] <= ((global_offset_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[2] <= ((global_offset_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'hC:
				begin
					kernel_arguments_NO_SHIFT_REG[31:0] <= ((kernel_arguments_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[63:32] <= ((kernel_arguments_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'hD:
				begin
					kernel_arguments_NO_SHIFT_REG[95:64] <= ((kernel_arguments_NO_SHIFT_REG[95:64] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[127:96] <= ((kernel_arguments_NO_SHIFT_REG[127:96] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				4'hE:
				begin
					kernel_arguments_NO_SHIFT_REG[159:128] <= ((kernel_arguments_NO_SHIFT_REG[159:128] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[191:160] <= ((kernel_arguments_NO_SHIFT_REG[191:160] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				default:
				begin
				end

			endcase
		end
		else
		begin
			if (status_NO_SHIFT_REG[0])
			begin
				start_NO_SHIFT_REG <= 1'b1;
			end
			if (start_NO_SHIFT_REG)
			begin
				status_NO_SHIFT_REG[0] <= 1'b0;
				started_NO_SHIFT_REG <= 1'b1;
			end
			if (started_NO_SHIFT_REG)
			begin
				start_NO_SHIFT_REG <= 1'b0;
			end
			if (finish)
			begin
				status_NO_SHIFT_REG[1] <= 1'b1;
				started_NO_SHIFT_REG <= 1'b0;
			end
		end
		status_NO_SHIFT_REG[11] <= 1'b0;
		status_NO_SHIFT_REG[12] <= (|has_a_lsu_active);
		status_NO_SHIFT_REG[13] <= (|has_a_write_pending);
		status_NO_SHIFT_REG[14] <= (|valid_in);
		status_NO_SHIFT_REG[15] <= started_NO_SHIFT_REG;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cra_read_st1_NO_SHIFT_REG <= 1'b0;
		cra_addr_st1_NO_SHIFT_REG <= 4'h0;
		cra_readdata_st1_NO_SHIFT_REG <= 64'h0;
	end
	else
	begin
		cra_read_st1_NO_SHIFT_REG <= avs_cra_read;
		cra_addr_st1_NO_SHIFT_REG <= avs_cra_address;
		case (avs_cra_address)
			4'h0:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= status_NO_SHIFT_REG;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			4'h1:
			begin
				cra_readdata_st1_NO_SHIFT_REG[31:0] <= 'x;
				cra_readdata_st1_NO_SHIFT_REG[63:32] <= 32'h0;
			end

			4'h2:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			4'h3:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			4'h4:
			begin
				cra_readdata_st1_NO_SHIFT_REG[63:0] <= 64'h0;
			end

			default:
			begin
				cra_readdata_st1_NO_SHIFT_REG <= status_NO_SHIFT_REG;
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		avs_cra_readdatavalid <= 1'b0;
		avs_cra_readdata <= 64'h0;
	end
	else
	begin
		avs_cra_readdatavalid <= cra_read_st1_NO_SHIFT_REG;
		case (cra_addr_st1_NO_SHIFT_REG)
			4'h2:
			begin
				avs_cra_readdata[63:0] <= profile_data_NO_SHIFT_REG;
			end

			default:
			begin
				avs_cra_readdata <= cra_readdata_st1_NO_SHIFT_REG;
			end

		endcase
	end
end


// Handshaking signals used to control data through the pipeline

// Determine when the kernel is finished.
acl_kernel_finish_detector kernel_finish_detector (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.wg_size(workgroup_size_NO_SHIFT_REG),
	.wg_dispatch_valid_out(iter_valid_in),
	.wg_dispatch_stall_in(iter_stall_out),
	.dispatched_all_groups(dispatched_all_groups),
	.kernel_copy_valid_out(valid_out),
	.kernel_copy_stall_in(stall_in),
	.pending_writes(has_a_write_pending),
	.finish(finish)
);

defparam kernel_finish_detector.TESSELLATION_SIZE = 0;
defparam kernel_finish_detector.NUM_COPIES = 1;
defparam kernel_finish_detector.WG_SIZE_W = 32;

assign stall_in = 1'b0;

// Creating ID iterator and kernel instance for every requested kernel copy

// ID iterator is responsible for iterating over all local ids for given work-groups
acl_id_iterator id_iter_inst0 (
	.clock(clock),
	.resetn(resetn),
	.start(start_out),
	.valid_in(iter_valid_in),
	.stall_out(iter_stall_out),
	.stall_in(stall_out),
	.valid_out(valid_in),
	.group_id_in(group_id_tmp),
	.global_id_base_in(global_id_base_out),
	.local_size(local_size_NO_SHIFT_REG),
	.global_size(global_size_NO_SHIFT_REG),
	.local_id(local_id[0]),
	.global_id(global_id[0]),
	.group_id(group_id[0])
);



// This section instantiates a kernel function block
AOCbilateralFilterkernel_function AOCbilateralFilterkernel_function_inst0 (
	.clock(clock),
	.resetn(resetn),
	.stall_out(stall_out),
	.valid_in(valid_in),
	.valid_out(valid_out),
	.stall_in(stall_in),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__inst0_readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__inst0_readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__inst0_waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__inst0_address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__inst0_read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__inst0_write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__inst0_writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__inst0_writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__inst0_byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__inst0_burstcount),
	.avm_local_bb4_ld__readdata(avm_local_bb4_ld__inst0_readdata),
	.avm_local_bb4_ld__readdatavalid(avm_local_bb4_ld__inst0_readdatavalid),
	.avm_local_bb4_ld__waitrequest(avm_local_bb4_ld__inst0_waitrequest),
	.avm_local_bb4_ld__address(avm_local_bb4_ld__inst0_address),
	.avm_local_bb4_ld__read(avm_local_bb4_ld__inst0_read),
	.avm_local_bb4_ld__write(avm_local_bb4_ld__inst0_write),
	.avm_local_bb4_ld__writeack(avm_local_bb4_ld__inst0_writeack),
	.avm_local_bb4_ld__writedata(avm_local_bb4_ld__inst0_writedata),
	.avm_local_bb4_ld__byteenable(avm_local_bb4_ld__inst0_byteenable),
	.avm_local_bb4_ld__burstcount(avm_local_bb4_ld__inst0_burstcount),
	.avm_local_bb6_st_c0_exe239_readdata(avm_local_bb6_st_c0_exe239_inst0_readdata),
	.avm_local_bb6_st_c0_exe239_readdatavalid(avm_local_bb6_st_c0_exe239_inst0_readdatavalid),
	.avm_local_bb6_st_c0_exe239_waitrequest(avm_local_bb6_st_c0_exe239_inst0_waitrequest),
	.avm_local_bb6_st_c0_exe239_address(avm_local_bb6_st_c0_exe239_inst0_address),
	.avm_local_bb6_st_c0_exe239_read(avm_local_bb6_st_c0_exe239_inst0_read),
	.avm_local_bb6_st_c0_exe239_write(avm_local_bb6_st_c0_exe239_inst0_write),
	.avm_local_bb6_st_c0_exe239_writeack(avm_local_bb6_st_c0_exe239_inst0_writeack),
	.avm_local_bb6_st_c0_exe239_writedata(avm_local_bb6_st_c0_exe239_inst0_writedata),
	.avm_local_bb6_st_c0_exe239_byteenable(avm_local_bb6_st_c0_exe239_inst0_byteenable),
	.avm_local_bb6_st_c0_exe239_burstcount(avm_local_bb6_st_c0_exe239_inst0_burstcount),
	.avm_local_bb8_st__readdata(avm_local_bb8_st__inst0_readdata),
	.avm_local_bb8_st__readdatavalid(avm_local_bb8_st__inst0_readdatavalid),
	.avm_local_bb8_st__waitrequest(avm_local_bb8_st__inst0_waitrequest),
	.avm_local_bb8_st__address(avm_local_bb8_st__inst0_address),
	.avm_local_bb8_st__read(avm_local_bb8_st__inst0_read),
	.avm_local_bb8_st__write(avm_local_bb8_st__inst0_write),
	.avm_local_bb8_st__writeack(avm_local_bb8_st__inst0_writeack),
	.avm_local_bb8_st__writedata(avm_local_bb8_st__inst0_writedata),
	.avm_local_bb8_st__byteenable(avm_local_bb8_st__inst0_byteenable),
	.avm_local_bb8_st__burstcount(avm_local_bb8_st__inst0_burstcount),
	.start(start_out),
	.input_r(kernel_arguments_NO_SHIFT_REG[191:160]),
	.input_global_size_0(global_size_NO_SHIFT_REG[0]),
	.input_global_size_1(global_size_NO_SHIFT_REG[1]),
	.input_e_d(kernel_arguments_NO_SHIFT_REG[159:128]),
	.clock2x(clock2x),
	.input_in(kernel_arguments_NO_SHIFT_REG[127:64]),
	.input_out(kernel_arguments_NO_SHIFT_REG[63:0]),
	.has_a_write_pending(has_a_write_pending),
	.has_a_lsu_active(has_a_lsu_active)
);



endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

// altera message_off 10036
// altera message_off 10230
// altera message_off 10858
module AOCbilateralFilterkernel_sys_cycle_time
	(
		input 		clock,
		input 		resetn,
		output [31:0] 		cur_cycle
	);


 reg [31:0] cur_count_NO_SHIFT_REG;

assign cur_cycle = cur_count_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cur_count_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		cur_count_NO_SHIFT_REG <= (cur_count_NO_SHIFT_REG + 32'h1);
	end
end

endmodule

